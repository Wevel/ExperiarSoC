// This is the unpowered netlist.
module ExperiarCore (clk0,
    clk1,
    core_wb_ack_i,
    core_wb_cyc_o,
    core_wb_error_i,
    core_wb_stall_i,
    core_wb_stb_o,
    core_wb_we_o,
    jtag_tck,
    jtag_tdi,
    jtag_tdo,
    jtag_tms,
    localMemory_wb_ack_o,
    localMemory_wb_cyc_i,
    localMemory_wb_error_o,
    localMemory_wb_stall_o,
    localMemory_wb_stb_i,
    localMemory_wb_we_i,
    probe_state,
    wb_clk_i,
    wb_rst_i,
    web0,
    addr0,
    addr1,
    coreIndex,
    core_wb_adr_o,
    core_wb_data_i,
    core_wb_data_o,
    core_wb_sel_o,
    csb0,
    csb1,
    din0,
    dout0,
    dout1,
    irq,
    localMemory_wb_adr_i,
    localMemory_wb_data_i,
    localMemory_wb_data_o,
    localMemory_wb_sel_i,
    manufacturerID,
    partID,
    probe_env,
    probe_jtagInstruction,
    probe_programCounter,
    versionID,
    wmask0);
 output clk0;
 output clk1;
 input core_wb_ack_i;
 output core_wb_cyc_o;
 input core_wb_error_i;
 input core_wb_stall_i;
 output core_wb_stb_o;
 output core_wb_we_o;
 input jtag_tck;
 input jtag_tdi;
 output jtag_tdo;
 input jtag_tms;
 output localMemory_wb_ack_o;
 input localMemory_wb_cyc_i;
 output localMemory_wb_error_o;
 output localMemory_wb_stall_o;
 input localMemory_wb_stb_i;
 input localMemory_wb_we_i;
 output probe_state;
 input wb_clk_i;
 input wb_rst_i;
 output web0;
 output [8:0] addr0;
 output [8:0] addr1;
 input [7:0] coreIndex;
 output [27:0] core_wb_adr_o;
 input [31:0] core_wb_data_i;
 output [31:0] core_wb_data_o;
 output [3:0] core_wb_sel_o;
 output [1:0] csb0;
 output [1:0] csb1;
 output [31:0] din0;
 input [63:0] dout0;
 input [63:0] dout1;
 input [15:0] irq;
 input [23:0] localMemory_wb_adr_i;
 input [31:0] localMemory_wb_data_i;
 output [31:0] localMemory_wb_data_o;
 input [3:0] localMemory_wb_sel_i;
 input [10:0] manufacturerID;
 input [15:0] partID;
 output [1:0] probe_env;
 output [4:0] probe_jtagInstruction;
 output [31:0] probe_programCounter;
 input [3:0] versionID;
 output [3:0] wmask0;

 wire net1911;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0_0_wb_clk_i;
 wire clknet_2_1_0_wb_clk_i;
 wire clknet_2_2_0_wb_clk_i;
 wire clknet_2_3_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_131_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_133_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_leaf_136_wb_clk_i;
 wire clknet_leaf_137_wb_clk_i;
 wire clknet_leaf_138_wb_clk_i;
 wire clknet_leaf_139_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_140_wb_clk_i;
 wire clknet_leaf_141_wb_clk_i;
 wire clknet_leaf_142_wb_clk_i;
 wire clknet_leaf_143_wb_clk_i;
 wire clknet_leaf_144_wb_clk_i;
 wire clknet_leaf_145_wb_clk_i;
 wire clknet_leaf_146_wb_clk_i;
 wire clknet_leaf_147_wb_clk_i;
 wire clknet_leaf_148_wb_clk_i;
 wire clknet_leaf_149_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_150_wb_clk_i;
 wire clknet_leaf_151_wb_clk_i;
 wire clknet_leaf_152_wb_clk_i;
 wire clknet_leaf_153_wb_clk_i;
 wire clknet_leaf_154_wb_clk_i;
 wire clknet_leaf_155_wb_clk_i;
 wire clknet_leaf_156_wb_clk_i;
 wire clknet_leaf_157_wb_clk_i;
 wire clknet_leaf_158_wb_clk_i;
 wire clknet_leaf_159_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_160_wb_clk_i;
 wire clknet_leaf_161_wb_clk_i;
 wire clknet_leaf_162_wb_clk_i;
 wire clknet_leaf_163_wb_clk_i;
 wire clknet_leaf_164_wb_clk_i;
 wire clknet_leaf_165_wb_clk_i;
 wire clknet_leaf_166_wb_clk_i;
 wire clknet_leaf_167_wb_clk_i;
 wire clknet_leaf_168_wb_clk_i;
 wire clknet_leaf_169_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_170_wb_clk_i;
 wire clknet_leaf_171_wb_clk_i;
 wire clknet_leaf_172_wb_clk_i;
 wire clknet_leaf_173_wb_clk_i;
 wire clknet_leaf_174_wb_clk_i;
 wire clknet_leaf_175_wb_clk_i;
 wire clknet_leaf_176_wb_clk_i;
 wire clknet_leaf_177_wb_clk_i;
 wire clknet_leaf_178_wb_clk_i;
 wire clknet_leaf_179_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_180_wb_clk_i;
 wire clknet_leaf_181_wb_clk_i;
 wire clknet_leaf_182_wb_clk_i;
 wire clknet_leaf_183_wb_clk_i;
 wire clknet_leaf_184_wb_clk_i;
 wire clknet_leaf_185_wb_clk_i;
 wire clknet_leaf_186_wb_clk_i;
 wire clknet_leaf_187_wb_clk_i;
 wire clknet_leaf_188_wb_clk_i;
 wire clknet_leaf_189_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_190_wb_clk_i;
 wire clknet_leaf_191_wb_clk_i;
 wire clknet_leaf_192_wb_clk_i;
 wire clknet_leaf_193_wb_clk_i;
 wire clknet_leaf_194_wb_clk_i;
 wire clknet_leaf_195_wb_clk_i;
 wire clknet_leaf_196_wb_clk_i;
 wire clknet_leaf_197_wb_clk_i;
 wire clknet_leaf_198_wb_clk_i;
 wire clknet_leaf_199_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_200_wb_clk_i;
 wire clknet_leaf_201_wb_clk_i;
 wire clknet_leaf_202_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire \core.cancelStall ;
 wire \core.csr.currentInstruction[0] ;
 wire \core.csr.currentInstruction[10] ;
 wire \core.csr.currentInstruction[11] ;
 wire \core.csr.currentInstruction[12] ;
 wire \core.csr.currentInstruction[13] ;
 wire \core.csr.currentInstruction[14] ;
 wire \core.csr.currentInstruction[15] ;
 wire \core.csr.currentInstruction[16] ;
 wire \core.csr.currentInstruction[17] ;
 wire \core.csr.currentInstruction[18] ;
 wire \core.csr.currentInstruction[19] ;
 wire \core.csr.currentInstruction[1] ;
 wire \core.csr.currentInstruction[20] ;
 wire \core.csr.currentInstruction[21] ;
 wire \core.csr.currentInstruction[22] ;
 wire \core.csr.currentInstruction[23] ;
 wire \core.csr.currentInstruction[24] ;
 wire \core.csr.currentInstruction[25] ;
 wire \core.csr.currentInstruction[26] ;
 wire \core.csr.currentInstruction[27] ;
 wire \core.csr.currentInstruction[28] ;
 wire \core.csr.currentInstruction[29] ;
 wire \core.csr.currentInstruction[2] ;
 wire \core.csr.currentInstruction[30] ;
 wire \core.csr.currentInstruction[31] ;
 wire \core.csr.currentInstruction[3] ;
 wire \core.csr.currentInstruction[4] ;
 wire \core.csr.currentInstruction[5] ;
 wire \core.csr.currentInstruction[6] ;
 wire \core.csr.currentInstruction[7] ;
 wire \core.csr.currentInstruction[8] ;
 wire \core.csr.currentInstruction[9] ;
 wire \core.csr.cycleTimer.currentValue[0] ;
 wire \core.csr.cycleTimer.currentValue[10] ;
 wire \core.csr.cycleTimer.currentValue[11] ;
 wire \core.csr.cycleTimer.currentValue[12] ;
 wire \core.csr.cycleTimer.currentValue[13] ;
 wire \core.csr.cycleTimer.currentValue[14] ;
 wire \core.csr.cycleTimer.currentValue[15] ;
 wire \core.csr.cycleTimer.currentValue[16] ;
 wire \core.csr.cycleTimer.currentValue[17] ;
 wire \core.csr.cycleTimer.currentValue[18] ;
 wire \core.csr.cycleTimer.currentValue[19] ;
 wire \core.csr.cycleTimer.currentValue[1] ;
 wire \core.csr.cycleTimer.currentValue[20] ;
 wire \core.csr.cycleTimer.currentValue[21] ;
 wire \core.csr.cycleTimer.currentValue[22] ;
 wire \core.csr.cycleTimer.currentValue[23] ;
 wire \core.csr.cycleTimer.currentValue[24] ;
 wire \core.csr.cycleTimer.currentValue[25] ;
 wire \core.csr.cycleTimer.currentValue[26] ;
 wire \core.csr.cycleTimer.currentValue[27] ;
 wire \core.csr.cycleTimer.currentValue[28] ;
 wire \core.csr.cycleTimer.currentValue[29] ;
 wire \core.csr.cycleTimer.currentValue[2] ;
 wire \core.csr.cycleTimer.currentValue[30] ;
 wire \core.csr.cycleTimer.currentValue[31] ;
 wire \core.csr.cycleTimer.currentValue[32] ;
 wire \core.csr.cycleTimer.currentValue[33] ;
 wire \core.csr.cycleTimer.currentValue[34] ;
 wire \core.csr.cycleTimer.currentValue[35] ;
 wire \core.csr.cycleTimer.currentValue[36] ;
 wire \core.csr.cycleTimer.currentValue[37] ;
 wire \core.csr.cycleTimer.currentValue[38] ;
 wire \core.csr.cycleTimer.currentValue[39] ;
 wire \core.csr.cycleTimer.currentValue[3] ;
 wire \core.csr.cycleTimer.currentValue[40] ;
 wire \core.csr.cycleTimer.currentValue[41] ;
 wire \core.csr.cycleTimer.currentValue[42] ;
 wire \core.csr.cycleTimer.currentValue[43] ;
 wire \core.csr.cycleTimer.currentValue[44] ;
 wire \core.csr.cycleTimer.currentValue[45] ;
 wire \core.csr.cycleTimer.currentValue[46] ;
 wire \core.csr.cycleTimer.currentValue[47] ;
 wire \core.csr.cycleTimer.currentValue[48] ;
 wire \core.csr.cycleTimer.currentValue[49] ;
 wire \core.csr.cycleTimer.currentValue[4] ;
 wire \core.csr.cycleTimer.currentValue[50] ;
 wire \core.csr.cycleTimer.currentValue[51] ;
 wire \core.csr.cycleTimer.currentValue[52] ;
 wire \core.csr.cycleTimer.currentValue[53] ;
 wire \core.csr.cycleTimer.currentValue[54] ;
 wire \core.csr.cycleTimer.currentValue[55] ;
 wire \core.csr.cycleTimer.currentValue[56] ;
 wire \core.csr.cycleTimer.currentValue[57] ;
 wire \core.csr.cycleTimer.currentValue[58] ;
 wire \core.csr.cycleTimer.currentValue[59] ;
 wire \core.csr.cycleTimer.currentValue[5] ;
 wire \core.csr.cycleTimer.currentValue[60] ;
 wire \core.csr.cycleTimer.currentValue[61] ;
 wire \core.csr.cycleTimer.currentValue[62] ;
 wire \core.csr.cycleTimer.currentValue[63] ;
 wire \core.csr.cycleTimer.currentValue[6] ;
 wire \core.csr.cycleTimer.currentValue[7] ;
 wire \core.csr.cycleTimer.currentValue[8] ;
 wire \core.csr.cycleTimer.currentValue[9] ;
 wire \core.csr.instretTimer.currentValue[0] ;
 wire \core.csr.instretTimer.currentValue[10] ;
 wire \core.csr.instretTimer.currentValue[11] ;
 wire \core.csr.instretTimer.currentValue[12] ;
 wire \core.csr.instretTimer.currentValue[13] ;
 wire \core.csr.instretTimer.currentValue[14] ;
 wire \core.csr.instretTimer.currentValue[15] ;
 wire \core.csr.instretTimer.currentValue[16] ;
 wire \core.csr.instretTimer.currentValue[17] ;
 wire \core.csr.instretTimer.currentValue[18] ;
 wire \core.csr.instretTimer.currentValue[19] ;
 wire \core.csr.instretTimer.currentValue[1] ;
 wire \core.csr.instretTimer.currentValue[20] ;
 wire \core.csr.instretTimer.currentValue[21] ;
 wire \core.csr.instretTimer.currentValue[22] ;
 wire \core.csr.instretTimer.currentValue[23] ;
 wire \core.csr.instretTimer.currentValue[24] ;
 wire \core.csr.instretTimer.currentValue[25] ;
 wire \core.csr.instretTimer.currentValue[26] ;
 wire \core.csr.instretTimer.currentValue[27] ;
 wire \core.csr.instretTimer.currentValue[28] ;
 wire \core.csr.instretTimer.currentValue[29] ;
 wire \core.csr.instretTimer.currentValue[2] ;
 wire \core.csr.instretTimer.currentValue[30] ;
 wire \core.csr.instretTimer.currentValue[31] ;
 wire \core.csr.instretTimer.currentValue[32] ;
 wire \core.csr.instretTimer.currentValue[33] ;
 wire \core.csr.instretTimer.currentValue[34] ;
 wire \core.csr.instretTimer.currentValue[35] ;
 wire \core.csr.instretTimer.currentValue[36] ;
 wire \core.csr.instretTimer.currentValue[37] ;
 wire \core.csr.instretTimer.currentValue[38] ;
 wire \core.csr.instretTimer.currentValue[39] ;
 wire \core.csr.instretTimer.currentValue[3] ;
 wire \core.csr.instretTimer.currentValue[40] ;
 wire \core.csr.instretTimer.currentValue[41] ;
 wire \core.csr.instretTimer.currentValue[42] ;
 wire \core.csr.instretTimer.currentValue[43] ;
 wire \core.csr.instretTimer.currentValue[44] ;
 wire \core.csr.instretTimer.currentValue[45] ;
 wire \core.csr.instretTimer.currentValue[46] ;
 wire \core.csr.instretTimer.currentValue[47] ;
 wire \core.csr.instretTimer.currentValue[48] ;
 wire \core.csr.instretTimer.currentValue[49] ;
 wire \core.csr.instretTimer.currentValue[4] ;
 wire \core.csr.instretTimer.currentValue[50] ;
 wire \core.csr.instretTimer.currentValue[51] ;
 wire \core.csr.instretTimer.currentValue[52] ;
 wire \core.csr.instretTimer.currentValue[53] ;
 wire \core.csr.instretTimer.currentValue[54] ;
 wire \core.csr.instretTimer.currentValue[55] ;
 wire \core.csr.instretTimer.currentValue[56] ;
 wire \core.csr.instretTimer.currentValue[57] ;
 wire \core.csr.instretTimer.currentValue[58] ;
 wire \core.csr.instretTimer.currentValue[59] ;
 wire \core.csr.instretTimer.currentValue[5] ;
 wire \core.csr.instretTimer.currentValue[60] ;
 wire \core.csr.instretTimer.currentValue[61] ;
 wire \core.csr.instretTimer.currentValue[62] ;
 wire \core.csr.instretTimer.currentValue[63] ;
 wire \core.csr.instretTimer.currentValue[6] ;
 wire \core.csr.instretTimer.currentValue[7] ;
 wire \core.csr.instretTimer.currentValue[8] ;
 wire \core.csr.instretTimer.currentValue[9] ;
 wire \core.csr.mconfigptr.currentValue[0] ;
 wire \core.csr.mconfigptr.currentValue[10] ;
 wire \core.csr.mconfigptr.currentValue[11] ;
 wire \core.csr.mconfigptr.currentValue[12] ;
 wire \core.csr.mconfigptr.currentValue[13] ;
 wire \core.csr.mconfigptr.currentValue[14] ;
 wire \core.csr.mconfigptr.currentValue[15] ;
 wire \core.csr.mconfigptr.currentValue[16] ;
 wire \core.csr.mconfigptr.currentValue[17] ;
 wire \core.csr.mconfigptr.currentValue[18] ;
 wire \core.csr.mconfigptr.currentValue[19] ;
 wire \core.csr.mconfigptr.currentValue[1] ;
 wire \core.csr.mconfigptr.currentValue[20] ;
 wire \core.csr.mconfigptr.currentValue[21] ;
 wire \core.csr.mconfigptr.currentValue[22] ;
 wire \core.csr.mconfigptr.currentValue[23] ;
 wire \core.csr.mconfigptr.currentValue[24] ;
 wire \core.csr.mconfigptr.currentValue[25] ;
 wire \core.csr.mconfigptr.currentValue[26] ;
 wire \core.csr.mconfigptr.currentValue[27] ;
 wire \core.csr.mconfigptr.currentValue[28] ;
 wire \core.csr.mconfigptr.currentValue[29] ;
 wire \core.csr.mconfigptr.currentValue[2] ;
 wire \core.csr.mconfigptr.currentValue[30] ;
 wire \core.csr.mconfigptr.currentValue[31] ;
 wire \core.csr.mconfigptr.currentValue[3] ;
 wire \core.csr.mconfigptr.currentValue[4] ;
 wire \core.csr.mconfigptr.currentValue[5] ;
 wire \core.csr.mconfigptr.currentValue[6] ;
 wire \core.csr.mconfigptr.currentValue[7] ;
 wire \core.csr.mconfigptr.currentValue[8] ;
 wire \core.csr.mconfigptr.currentValue[9] ;
 wire \core.csr.trapReturnVector[0] ;
 wire \core.csr.trapReturnVector[10] ;
 wire \core.csr.trapReturnVector[11] ;
 wire \core.csr.trapReturnVector[12] ;
 wire \core.csr.trapReturnVector[13] ;
 wire \core.csr.trapReturnVector[14] ;
 wire \core.csr.trapReturnVector[15] ;
 wire \core.csr.trapReturnVector[16] ;
 wire \core.csr.trapReturnVector[17] ;
 wire \core.csr.trapReturnVector[18] ;
 wire \core.csr.trapReturnVector[19] ;
 wire \core.csr.trapReturnVector[1] ;
 wire \core.csr.trapReturnVector[20] ;
 wire \core.csr.trapReturnVector[21] ;
 wire \core.csr.trapReturnVector[22] ;
 wire \core.csr.trapReturnVector[23] ;
 wire \core.csr.trapReturnVector[24] ;
 wire \core.csr.trapReturnVector[25] ;
 wire \core.csr.trapReturnVector[26] ;
 wire \core.csr.trapReturnVector[27] ;
 wire \core.csr.trapReturnVector[28] ;
 wire \core.csr.trapReturnVector[29] ;
 wire \core.csr.trapReturnVector[2] ;
 wire \core.csr.trapReturnVector[30] ;
 wire \core.csr.trapReturnVector[31] ;
 wire \core.csr.trapReturnVector[3] ;
 wire \core.csr.trapReturnVector[4] ;
 wire \core.csr.trapReturnVector[5] ;
 wire \core.csr.trapReturnVector[6] ;
 wire \core.csr.trapReturnVector[7] ;
 wire \core.csr.trapReturnVector[8] ;
 wire \core.csr.trapReturnVector[9] ;
 wire \core.csr.traps.machineInterruptEnable ;
 wire \core.csr.traps.machinePreviousInterruptEnable ;
 wire \core.csr.traps.mcause.csrReadData[0] ;
 wire \core.csr.traps.mcause.csrReadData[10] ;
 wire \core.csr.traps.mcause.csrReadData[11] ;
 wire \core.csr.traps.mcause.csrReadData[12] ;
 wire \core.csr.traps.mcause.csrReadData[13] ;
 wire \core.csr.traps.mcause.csrReadData[14] ;
 wire \core.csr.traps.mcause.csrReadData[15] ;
 wire \core.csr.traps.mcause.csrReadData[16] ;
 wire \core.csr.traps.mcause.csrReadData[17] ;
 wire \core.csr.traps.mcause.csrReadData[18] ;
 wire \core.csr.traps.mcause.csrReadData[19] ;
 wire \core.csr.traps.mcause.csrReadData[1] ;
 wire \core.csr.traps.mcause.csrReadData[20] ;
 wire \core.csr.traps.mcause.csrReadData[21] ;
 wire \core.csr.traps.mcause.csrReadData[22] ;
 wire \core.csr.traps.mcause.csrReadData[23] ;
 wire \core.csr.traps.mcause.csrReadData[24] ;
 wire \core.csr.traps.mcause.csrReadData[25] ;
 wire \core.csr.traps.mcause.csrReadData[26] ;
 wire \core.csr.traps.mcause.csrReadData[27] ;
 wire \core.csr.traps.mcause.csrReadData[28] ;
 wire \core.csr.traps.mcause.csrReadData[29] ;
 wire \core.csr.traps.mcause.csrReadData[2] ;
 wire \core.csr.traps.mcause.csrReadData[30] ;
 wire \core.csr.traps.mcause.csrReadData[31] ;
 wire \core.csr.traps.mcause.csrReadData[3] ;
 wire \core.csr.traps.mcause.csrReadData[4] ;
 wire \core.csr.traps.mcause.csrReadData[5] ;
 wire \core.csr.traps.mcause.csrReadData[6] ;
 wire \core.csr.traps.mcause.csrReadData[7] ;
 wire \core.csr.traps.mcause.csrReadData[8] ;
 wire \core.csr.traps.mcause.csrReadData[9] ;
 wire \core.csr.traps.mie.currentValue[0] ;
 wire \core.csr.traps.mie.currentValue[10] ;
 wire \core.csr.traps.mie.currentValue[11] ;
 wire \core.csr.traps.mie.currentValue[12] ;
 wire \core.csr.traps.mie.currentValue[13] ;
 wire \core.csr.traps.mie.currentValue[14] ;
 wire \core.csr.traps.mie.currentValue[15] ;
 wire \core.csr.traps.mie.currentValue[16] ;
 wire \core.csr.traps.mie.currentValue[17] ;
 wire \core.csr.traps.mie.currentValue[18] ;
 wire \core.csr.traps.mie.currentValue[19] ;
 wire \core.csr.traps.mie.currentValue[1] ;
 wire \core.csr.traps.mie.currentValue[20] ;
 wire \core.csr.traps.mie.currentValue[21] ;
 wire \core.csr.traps.mie.currentValue[22] ;
 wire \core.csr.traps.mie.currentValue[23] ;
 wire \core.csr.traps.mie.currentValue[24] ;
 wire \core.csr.traps.mie.currentValue[25] ;
 wire \core.csr.traps.mie.currentValue[26] ;
 wire \core.csr.traps.mie.currentValue[27] ;
 wire \core.csr.traps.mie.currentValue[28] ;
 wire \core.csr.traps.mie.currentValue[29] ;
 wire \core.csr.traps.mie.currentValue[2] ;
 wire \core.csr.traps.mie.currentValue[30] ;
 wire \core.csr.traps.mie.currentValue[31] ;
 wire \core.csr.traps.mie.currentValue[3] ;
 wire \core.csr.traps.mie.currentValue[4] ;
 wire \core.csr.traps.mie.currentValue[5] ;
 wire \core.csr.traps.mie.currentValue[6] ;
 wire \core.csr.traps.mie.currentValue[7] ;
 wire \core.csr.traps.mie.currentValue[8] ;
 wire \core.csr.traps.mie.currentValue[9] ;
 wire \core.csr.traps.mip.csrReadData[0] ;
 wire \core.csr.traps.mip.csrReadData[10] ;
 wire \core.csr.traps.mip.csrReadData[11] ;
 wire \core.csr.traps.mip.csrReadData[12] ;
 wire \core.csr.traps.mip.csrReadData[13] ;
 wire \core.csr.traps.mip.csrReadData[14] ;
 wire \core.csr.traps.mip.csrReadData[15] ;
 wire \core.csr.traps.mip.csrReadData[16] ;
 wire \core.csr.traps.mip.csrReadData[17] ;
 wire \core.csr.traps.mip.csrReadData[18] ;
 wire \core.csr.traps.mip.csrReadData[19] ;
 wire \core.csr.traps.mip.csrReadData[1] ;
 wire \core.csr.traps.mip.csrReadData[20] ;
 wire \core.csr.traps.mip.csrReadData[21] ;
 wire \core.csr.traps.mip.csrReadData[22] ;
 wire \core.csr.traps.mip.csrReadData[23] ;
 wire \core.csr.traps.mip.csrReadData[24] ;
 wire \core.csr.traps.mip.csrReadData[25] ;
 wire \core.csr.traps.mip.csrReadData[26] ;
 wire \core.csr.traps.mip.csrReadData[27] ;
 wire \core.csr.traps.mip.csrReadData[28] ;
 wire \core.csr.traps.mip.csrReadData[29] ;
 wire \core.csr.traps.mip.csrReadData[2] ;
 wire \core.csr.traps.mip.csrReadData[30] ;
 wire \core.csr.traps.mip.csrReadData[31] ;
 wire \core.csr.traps.mip.csrReadData[3] ;
 wire \core.csr.traps.mip.csrReadData[4] ;
 wire \core.csr.traps.mip.csrReadData[5] ;
 wire \core.csr.traps.mip.csrReadData[6] ;
 wire \core.csr.traps.mip.csrReadData[7] ;
 wire \core.csr.traps.mip.csrReadData[8] ;
 wire \core.csr.traps.mip.csrReadData[9] ;
 wire \core.csr.traps.mscratch.currentValue[0] ;
 wire \core.csr.traps.mscratch.currentValue[10] ;
 wire \core.csr.traps.mscratch.currentValue[11] ;
 wire \core.csr.traps.mscratch.currentValue[12] ;
 wire \core.csr.traps.mscratch.currentValue[13] ;
 wire \core.csr.traps.mscratch.currentValue[14] ;
 wire \core.csr.traps.mscratch.currentValue[15] ;
 wire \core.csr.traps.mscratch.currentValue[16] ;
 wire \core.csr.traps.mscratch.currentValue[17] ;
 wire \core.csr.traps.mscratch.currentValue[18] ;
 wire \core.csr.traps.mscratch.currentValue[19] ;
 wire \core.csr.traps.mscratch.currentValue[1] ;
 wire \core.csr.traps.mscratch.currentValue[20] ;
 wire \core.csr.traps.mscratch.currentValue[21] ;
 wire \core.csr.traps.mscratch.currentValue[22] ;
 wire \core.csr.traps.mscratch.currentValue[23] ;
 wire \core.csr.traps.mscratch.currentValue[24] ;
 wire \core.csr.traps.mscratch.currentValue[25] ;
 wire \core.csr.traps.mscratch.currentValue[26] ;
 wire \core.csr.traps.mscratch.currentValue[27] ;
 wire \core.csr.traps.mscratch.currentValue[28] ;
 wire \core.csr.traps.mscratch.currentValue[29] ;
 wire \core.csr.traps.mscratch.currentValue[2] ;
 wire \core.csr.traps.mscratch.currentValue[30] ;
 wire \core.csr.traps.mscratch.currentValue[31] ;
 wire \core.csr.traps.mscratch.currentValue[3] ;
 wire \core.csr.traps.mscratch.currentValue[4] ;
 wire \core.csr.traps.mscratch.currentValue[5] ;
 wire \core.csr.traps.mscratch.currentValue[6] ;
 wire \core.csr.traps.mscratch.currentValue[7] ;
 wire \core.csr.traps.mscratch.currentValue[8] ;
 wire \core.csr.traps.mscratch.currentValue[9] ;
 wire \core.csr.traps.mtval.csrReadData[0] ;
 wire \core.csr.traps.mtval.csrReadData[10] ;
 wire \core.csr.traps.mtval.csrReadData[11] ;
 wire \core.csr.traps.mtval.csrReadData[12] ;
 wire \core.csr.traps.mtval.csrReadData[13] ;
 wire \core.csr.traps.mtval.csrReadData[14] ;
 wire \core.csr.traps.mtval.csrReadData[15] ;
 wire \core.csr.traps.mtval.csrReadData[16] ;
 wire \core.csr.traps.mtval.csrReadData[17] ;
 wire \core.csr.traps.mtval.csrReadData[18] ;
 wire \core.csr.traps.mtval.csrReadData[19] ;
 wire \core.csr.traps.mtval.csrReadData[1] ;
 wire \core.csr.traps.mtval.csrReadData[20] ;
 wire \core.csr.traps.mtval.csrReadData[21] ;
 wire \core.csr.traps.mtval.csrReadData[22] ;
 wire \core.csr.traps.mtval.csrReadData[23] ;
 wire \core.csr.traps.mtval.csrReadData[24] ;
 wire \core.csr.traps.mtval.csrReadData[25] ;
 wire \core.csr.traps.mtval.csrReadData[26] ;
 wire \core.csr.traps.mtval.csrReadData[27] ;
 wire \core.csr.traps.mtval.csrReadData[28] ;
 wire \core.csr.traps.mtval.csrReadData[29] ;
 wire \core.csr.traps.mtval.csrReadData[2] ;
 wire \core.csr.traps.mtval.csrReadData[30] ;
 wire \core.csr.traps.mtval.csrReadData[31] ;
 wire \core.csr.traps.mtval.csrReadData[3] ;
 wire \core.csr.traps.mtval.csrReadData[4] ;
 wire \core.csr.traps.mtval.csrReadData[5] ;
 wire \core.csr.traps.mtval.csrReadData[6] ;
 wire \core.csr.traps.mtval.csrReadData[7] ;
 wire \core.csr.traps.mtval.csrReadData[8] ;
 wire \core.csr.traps.mtval.csrReadData[9] ;
 wire \core.csr.traps.mtvec.csrReadData[0] ;
 wire \core.csr.traps.mtvec.csrReadData[10] ;
 wire \core.csr.traps.mtvec.csrReadData[11] ;
 wire \core.csr.traps.mtvec.csrReadData[12] ;
 wire \core.csr.traps.mtvec.csrReadData[13] ;
 wire \core.csr.traps.mtvec.csrReadData[14] ;
 wire \core.csr.traps.mtvec.csrReadData[15] ;
 wire \core.csr.traps.mtvec.csrReadData[16] ;
 wire \core.csr.traps.mtvec.csrReadData[17] ;
 wire \core.csr.traps.mtvec.csrReadData[18] ;
 wire \core.csr.traps.mtvec.csrReadData[19] ;
 wire \core.csr.traps.mtvec.csrReadData[1] ;
 wire \core.csr.traps.mtvec.csrReadData[20] ;
 wire \core.csr.traps.mtvec.csrReadData[21] ;
 wire \core.csr.traps.mtvec.csrReadData[22] ;
 wire \core.csr.traps.mtvec.csrReadData[23] ;
 wire \core.csr.traps.mtvec.csrReadData[24] ;
 wire \core.csr.traps.mtvec.csrReadData[25] ;
 wire \core.csr.traps.mtvec.csrReadData[26] ;
 wire \core.csr.traps.mtvec.csrReadData[27] ;
 wire \core.csr.traps.mtvec.csrReadData[28] ;
 wire \core.csr.traps.mtvec.csrReadData[29] ;
 wire \core.csr.traps.mtvec.csrReadData[2] ;
 wire \core.csr.traps.mtvec.csrReadData[30] ;
 wire \core.csr.traps.mtvec.csrReadData[31] ;
 wire \core.csr.traps.mtvec.csrReadData[3] ;
 wire \core.csr.traps.mtvec.csrReadData[4] ;
 wire \core.csr.traps.mtvec.csrReadData[5] ;
 wire \core.csr.traps.mtvec.csrReadData[6] ;
 wire \core.csr.traps.mtvec.csrReadData[7] ;
 wire \core.csr.traps.mtvec.csrReadData[8] ;
 wire \core.csr.traps.mtvec.csrReadData[9] ;
 wire \core.fetchProgramCounter[0] ;
 wire \core.fetchProgramCounter[10] ;
 wire \core.fetchProgramCounter[11] ;
 wire \core.fetchProgramCounter[12] ;
 wire \core.fetchProgramCounter[13] ;
 wire \core.fetchProgramCounter[14] ;
 wire \core.fetchProgramCounter[15] ;
 wire \core.fetchProgramCounter[16] ;
 wire \core.fetchProgramCounter[17] ;
 wire \core.fetchProgramCounter[18] ;
 wire \core.fetchProgramCounter[19] ;
 wire \core.fetchProgramCounter[1] ;
 wire \core.fetchProgramCounter[20] ;
 wire \core.fetchProgramCounter[21] ;
 wire \core.fetchProgramCounter[22] ;
 wire \core.fetchProgramCounter[23] ;
 wire \core.fetchProgramCounter[24] ;
 wire \core.fetchProgramCounter[25] ;
 wire \core.fetchProgramCounter[26] ;
 wire \core.fetchProgramCounter[27] ;
 wire \core.fetchProgramCounter[28] ;
 wire \core.fetchProgramCounter[29] ;
 wire \core.fetchProgramCounter[2] ;
 wire \core.fetchProgramCounter[30] ;
 wire \core.fetchProgramCounter[31] ;
 wire \core.fetchProgramCounter[3] ;
 wire \core.fetchProgramCounter[4] ;
 wire \core.fetchProgramCounter[5] ;
 wire \core.fetchProgramCounter[6] ;
 wire \core.fetchProgramCounter[7] ;
 wire \core.fetchProgramCounter[8] ;
 wire \core.fetchProgramCounter[9] ;
 wire \core.management_interruptEnable ;
 wire \core.management_run ;
 wire \core.pipe0_currentInstruction[0] ;
 wire \core.pipe0_currentInstruction[10] ;
 wire \core.pipe0_currentInstruction[11] ;
 wire \core.pipe0_currentInstruction[12] ;
 wire \core.pipe0_currentInstruction[13] ;
 wire \core.pipe0_currentInstruction[14] ;
 wire \core.pipe0_currentInstruction[15] ;
 wire \core.pipe0_currentInstruction[16] ;
 wire \core.pipe0_currentInstruction[17] ;
 wire \core.pipe0_currentInstruction[18] ;
 wire \core.pipe0_currentInstruction[19] ;
 wire \core.pipe0_currentInstruction[1] ;
 wire \core.pipe0_currentInstruction[20] ;
 wire \core.pipe0_currentInstruction[21] ;
 wire \core.pipe0_currentInstruction[22] ;
 wire \core.pipe0_currentInstruction[23] ;
 wire \core.pipe0_currentInstruction[24] ;
 wire \core.pipe0_currentInstruction[25] ;
 wire \core.pipe0_currentInstruction[26] ;
 wire \core.pipe0_currentInstruction[27] ;
 wire \core.pipe0_currentInstruction[28] ;
 wire \core.pipe0_currentInstruction[29] ;
 wire \core.pipe0_currentInstruction[2] ;
 wire \core.pipe0_currentInstruction[30] ;
 wire \core.pipe0_currentInstruction[31] ;
 wire \core.pipe0_currentInstruction[3] ;
 wire \core.pipe0_currentInstruction[4] ;
 wire \core.pipe0_currentInstruction[5] ;
 wire \core.pipe0_currentInstruction[6] ;
 wire \core.pipe0_currentInstruction[7] ;
 wire \core.pipe0_currentInstruction[8] ;
 wire \core.pipe0_currentInstruction[9] ;
 wire \core.pipe0_fetch.currentPipeStall ;
 wire \core.pipe0_fetch.lastProgramCounter[0] ;
 wire \core.pipe0_fetch.lastProgramCounter[10] ;
 wire \core.pipe0_fetch.lastProgramCounter[11] ;
 wire \core.pipe0_fetch.lastProgramCounter[12] ;
 wire \core.pipe0_fetch.lastProgramCounter[13] ;
 wire \core.pipe0_fetch.lastProgramCounter[14] ;
 wire \core.pipe0_fetch.lastProgramCounter[15] ;
 wire \core.pipe0_fetch.lastProgramCounter[16] ;
 wire \core.pipe0_fetch.lastProgramCounter[17] ;
 wire \core.pipe0_fetch.lastProgramCounter[18] ;
 wire \core.pipe0_fetch.lastProgramCounter[19] ;
 wire \core.pipe0_fetch.lastProgramCounter[1] ;
 wire \core.pipe0_fetch.lastProgramCounter[20] ;
 wire \core.pipe0_fetch.lastProgramCounter[21] ;
 wire \core.pipe0_fetch.lastProgramCounter[22] ;
 wire \core.pipe0_fetch.lastProgramCounter[23] ;
 wire \core.pipe0_fetch.lastProgramCounter[24] ;
 wire \core.pipe0_fetch.lastProgramCounter[25] ;
 wire \core.pipe0_fetch.lastProgramCounter[26] ;
 wire \core.pipe0_fetch.lastProgramCounter[27] ;
 wire \core.pipe0_fetch.lastProgramCounter[28] ;
 wire \core.pipe0_fetch.lastProgramCounter[29] ;
 wire \core.pipe0_fetch.lastProgramCounter[2] ;
 wire \core.pipe0_fetch.lastProgramCounter[30] ;
 wire \core.pipe0_fetch.lastProgramCounter[31] ;
 wire \core.pipe0_fetch.lastProgramCounter[3] ;
 wire \core.pipe0_fetch.lastProgramCounter[4] ;
 wire \core.pipe0_fetch.lastProgramCounter[5] ;
 wire \core.pipe0_fetch.lastProgramCounter[6] ;
 wire \core.pipe0_fetch.lastProgramCounter[7] ;
 wire \core.pipe0_fetch.lastProgramCounter[8] ;
 wire \core.pipe0_fetch.lastProgramCounter[9] ;
 wire \core.pipe1_csrData[0] ;
 wire \core.pipe1_csrData[10] ;
 wire \core.pipe1_csrData[11] ;
 wire \core.pipe1_csrData[12] ;
 wire \core.pipe1_csrData[13] ;
 wire \core.pipe1_csrData[14] ;
 wire \core.pipe1_csrData[15] ;
 wire \core.pipe1_csrData[16] ;
 wire \core.pipe1_csrData[17] ;
 wire \core.pipe1_csrData[18] ;
 wire \core.pipe1_csrData[19] ;
 wire \core.pipe1_csrData[1] ;
 wire \core.pipe1_csrData[20] ;
 wire \core.pipe1_csrData[21] ;
 wire \core.pipe1_csrData[22] ;
 wire \core.pipe1_csrData[23] ;
 wire \core.pipe1_csrData[24] ;
 wire \core.pipe1_csrData[25] ;
 wire \core.pipe1_csrData[26] ;
 wire \core.pipe1_csrData[27] ;
 wire \core.pipe1_csrData[28] ;
 wire \core.pipe1_csrData[29] ;
 wire \core.pipe1_csrData[2] ;
 wire \core.pipe1_csrData[30] ;
 wire \core.pipe1_csrData[31] ;
 wire \core.pipe1_csrData[3] ;
 wire \core.pipe1_csrData[4] ;
 wire \core.pipe1_csrData[5] ;
 wire \core.pipe1_csrData[6] ;
 wire \core.pipe1_csrData[7] ;
 wire \core.pipe1_csrData[8] ;
 wire \core.pipe1_csrData[9] ;
 wire \core.pipe1_operation.currentPipeStall ;
 wire \core.pipe1_resultRegister[0] ;
 wire \core.pipe1_resultRegister[10] ;
 wire \core.pipe1_resultRegister[11] ;
 wire \core.pipe1_resultRegister[12] ;
 wire \core.pipe1_resultRegister[13] ;
 wire \core.pipe1_resultRegister[14] ;
 wire \core.pipe1_resultRegister[15] ;
 wire \core.pipe1_resultRegister[16] ;
 wire \core.pipe1_resultRegister[17] ;
 wire \core.pipe1_resultRegister[18] ;
 wire \core.pipe1_resultRegister[19] ;
 wire \core.pipe1_resultRegister[1] ;
 wire \core.pipe1_resultRegister[20] ;
 wire \core.pipe1_resultRegister[21] ;
 wire \core.pipe1_resultRegister[22] ;
 wire \core.pipe1_resultRegister[23] ;
 wire \core.pipe1_resultRegister[24] ;
 wire \core.pipe1_resultRegister[25] ;
 wire \core.pipe1_resultRegister[26] ;
 wire \core.pipe1_resultRegister[27] ;
 wire \core.pipe1_resultRegister[28] ;
 wire \core.pipe1_resultRegister[29] ;
 wire \core.pipe1_resultRegister[2] ;
 wire \core.pipe1_resultRegister[30] ;
 wire \core.pipe1_resultRegister[31] ;
 wire \core.pipe1_resultRegister[3] ;
 wire \core.pipe1_resultRegister[4] ;
 wire \core.pipe1_resultRegister[5] ;
 wire \core.pipe1_resultRegister[6] ;
 wire \core.pipe1_resultRegister[7] ;
 wire \core.pipe1_resultRegister[8] ;
 wire \core.pipe1_resultRegister[9] ;
 wire \core.pipe2_stall ;
 wire \core.registers[0][0] ;
 wire \core.registers[0][10] ;
 wire \core.registers[0][11] ;
 wire \core.registers[0][12] ;
 wire \core.registers[0][13] ;
 wire \core.registers[0][14] ;
 wire \core.registers[0][15] ;
 wire \core.registers[0][16] ;
 wire \core.registers[0][17] ;
 wire \core.registers[0][18] ;
 wire \core.registers[0][19] ;
 wire \core.registers[0][1] ;
 wire \core.registers[0][20] ;
 wire \core.registers[0][21] ;
 wire \core.registers[0][22] ;
 wire \core.registers[0][23] ;
 wire \core.registers[0][24] ;
 wire \core.registers[0][25] ;
 wire \core.registers[0][26] ;
 wire \core.registers[0][27] ;
 wire \core.registers[0][28] ;
 wire \core.registers[0][29] ;
 wire \core.registers[0][2] ;
 wire \core.registers[0][30] ;
 wire \core.registers[0][31] ;
 wire \core.registers[0][3] ;
 wire \core.registers[0][4] ;
 wire \core.registers[0][5] ;
 wire \core.registers[0][6] ;
 wire \core.registers[0][7] ;
 wire \core.registers[0][8] ;
 wire \core.registers[0][9] ;
 wire \core.registers[10][0] ;
 wire \core.registers[10][10] ;
 wire \core.registers[10][11] ;
 wire \core.registers[10][12] ;
 wire \core.registers[10][13] ;
 wire \core.registers[10][14] ;
 wire \core.registers[10][15] ;
 wire \core.registers[10][16] ;
 wire \core.registers[10][17] ;
 wire \core.registers[10][18] ;
 wire \core.registers[10][19] ;
 wire \core.registers[10][1] ;
 wire \core.registers[10][20] ;
 wire \core.registers[10][21] ;
 wire \core.registers[10][22] ;
 wire \core.registers[10][23] ;
 wire \core.registers[10][24] ;
 wire \core.registers[10][25] ;
 wire \core.registers[10][26] ;
 wire \core.registers[10][27] ;
 wire \core.registers[10][28] ;
 wire \core.registers[10][29] ;
 wire \core.registers[10][2] ;
 wire \core.registers[10][30] ;
 wire \core.registers[10][31] ;
 wire \core.registers[10][3] ;
 wire \core.registers[10][4] ;
 wire \core.registers[10][5] ;
 wire \core.registers[10][6] ;
 wire \core.registers[10][7] ;
 wire \core.registers[10][8] ;
 wire \core.registers[10][9] ;
 wire \core.registers[11][0] ;
 wire \core.registers[11][10] ;
 wire \core.registers[11][11] ;
 wire \core.registers[11][12] ;
 wire \core.registers[11][13] ;
 wire \core.registers[11][14] ;
 wire \core.registers[11][15] ;
 wire \core.registers[11][16] ;
 wire \core.registers[11][17] ;
 wire \core.registers[11][18] ;
 wire \core.registers[11][19] ;
 wire \core.registers[11][1] ;
 wire \core.registers[11][20] ;
 wire \core.registers[11][21] ;
 wire \core.registers[11][22] ;
 wire \core.registers[11][23] ;
 wire \core.registers[11][24] ;
 wire \core.registers[11][25] ;
 wire \core.registers[11][26] ;
 wire \core.registers[11][27] ;
 wire \core.registers[11][28] ;
 wire \core.registers[11][29] ;
 wire \core.registers[11][2] ;
 wire \core.registers[11][30] ;
 wire \core.registers[11][31] ;
 wire \core.registers[11][3] ;
 wire \core.registers[11][4] ;
 wire \core.registers[11][5] ;
 wire \core.registers[11][6] ;
 wire \core.registers[11][7] ;
 wire \core.registers[11][8] ;
 wire \core.registers[11][9] ;
 wire \core.registers[12][0] ;
 wire \core.registers[12][10] ;
 wire \core.registers[12][11] ;
 wire \core.registers[12][12] ;
 wire \core.registers[12][13] ;
 wire \core.registers[12][14] ;
 wire \core.registers[12][15] ;
 wire \core.registers[12][16] ;
 wire \core.registers[12][17] ;
 wire \core.registers[12][18] ;
 wire \core.registers[12][19] ;
 wire \core.registers[12][1] ;
 wire \core.registers[12][20] ;
 wire \core.registers[12][21] ;
 wire \core.registers[12][22] ;
 wire \core.registers[12][23] ;
 wire \core.registers[12][24] ;
 wire \core.registers[12][25] ;
 wire \core.registers[12][26] ;
 wire \core.registers[12][27] ;
 wire \core.registers[12][28] ;
 wire \core.registers[12][29] ;
 wire \core.registers[12][2] ;
 wire \core.registers[12][30] ;
 wire \core.registers[12][31] ;
 wire \core.registers[12][3] ;
 wire \core.registers[12][4] ;
 wire \core.registers[12][5] ;
 wire \core.registers[12][6] ;
 wire \core.registers[12][7] ;
 wire \core.registers[12][8] ;
 wire \core.registers[12][9] ;
 wire \core.registers[13][0] ;
 wire \core.registers[13][10] ;
 wire \core.registers[13][11] ;
 wire \core.registers[13][12] ;
 wire \core.registers[13][13] ;
 wire \core.registers[13][14] ;
 wire \core.registers[13][15] ;
 wire \core.registers[13][16] ;
 wire \core.registers[13][17] ;
 wire \core.registers[13][18] ;
 wire \core.registers[13][19] ;
 wire \core.registers[13][1] ;
 wire \core.registers[13][20] ;
 wire \core.registers[13][21] ;
 wire \core.registers[13][22] ;
 wire \core.registers[13][23] ;
 wire \core.registers[13][24] ;
 wire \core.registers[13][25] ;
 wire \core.registers[13][26] ;
 wire \core.registers[13][27] ;
 wire \core.registers[13][28] ;
 wire \core.registers[13][29] ;
 wire \core.registers[13][2] ;
 wire \core.registers[13][30] ;
 wire \core.registers[13][31] ;
 wire \core.registers[13][3] ;
 wire \core.registers[13][4] ;
 wire \core.registers[13][5] ;
 wire \core.registers[13][6] ;
 wire \core.registers[13][7] ;
 wire \core.registers[13][8] ;
 wire \core.registers[13][9] ;
 wire \core.registers[14][0] ;
 wire \core.registers[14][10] ;
 wire \core.registers[14][11] ;
 wire \core.registers[14][12] ;
 wire \core.registers[14][13] ;
 wire \core.registers[14][14] ;
 wire \core.registers[14][15] ;
 wire \core.registers[14][16] ;
 wire \core.registers[14][17] ;
 wire \core.registers[14][18] ;
 wire \core.registers[14][19] ;
 wire \core.registers[14][1] ;
 wire \core.registers[14][20] ;
 wire \core.registers[14][21] ;
 wire \core.registers[14][22] ;
 wire \core.registers[14][23] ;
 wire \core.registers[14][24] ;
 wire \core.registers[14][25] ;
 wire \core.registers[14][26] ;
 wire \core.registers[14][27] ;
 wire \core.registers[14][28] ;
 wire \core.registers[14][29] ;
 wire \core.registers[14][2] ;
 wire \core.registers[14][30] ;
 wire \core.registers[14][31] ;
 wire \core.registers[14][3] ;
 wire \core.registers[14][4] ;
 wire \core.registers[14][5] ;
 wire \core.registers[14][6] ;
 wire \core.registers[14][7] ;
 wire \core.registers[14][8] ;
 wire \core.registers[14][9] ;
 wire \core.registers[15][0] ;
 wire \core.registers[15][10] ;
 wire \core.registers[15][11] ;
 wire \core.registers[15][12] ;
 wire \core.registers[15][13] ;
 wire \core.registers[15][14] ;
 wire \core.registers[15][15] ;
 wire \core.registers[15][16] ;
 wire \core.registers[15][17] ;
 wire \core.registers[15][18] ;
 wire \core.registers[15][19] ;
 wire \core.registers[15][1] ;
 wire \core.registers[15][20] ;
 wire \core.registers[15][21] ;
 wire \core.registers[15][22] ;
 wire \core.registers[15][23] ;
 wire \core.registers[15][24] ;
 wire \core.registers[15][25] ;
 wire \core.registers[15][26] ;
 wire \core.registers[15][27] ;
 wire \core.registers[15][28] ;
 wire \core.registers[15][29] ;
 wire \core.registers[15][2] ;
 wire \core.registers[15][30] ;
 wire \core.registers[15][31] ;
 wire \core.registers[15][3] ;
 wire \core.registers[15][4] ;
 wire \core.registers[15][5] ;
 wire \core.registers[15][6] ;
 wire \core.registers[15][7] ;
 wire \core.registers[15][8] ;
 wire \core.registers[15][9] ;
 wire \core.registers[16][0] ;
 wire \core.registers[16][10] ;
 wire \core.registers[16][11] ;
 wire \core.registers[16][12] ;
 wire \core.registers[16][13] ;
 wire \core.registers[16][14] ;
 wire \core.registers[16][15] ;
 wire \core.registers[16][16] ;
 wire \core.registers[16][17] ;
 wire \core.registers[16][18] ;
 wire \core.registers[16][19] ;
 wire \core.registers[16][1] ;
 wire \core.registers[16][20] ;
 wire \core.registers[16][21] ;
 wire \core.registers[16][22] ;
 wire \core.registers[16][23] ;
 wire \core.registers[16][24] ;
 wire \core.registers[16][25] ;
 wire \core.registers[16][26] ;
 wire \core.registers[16][27] ;
 wire \core.registers[16][28] ;
 wire \core.registers[16][29] ;
 wire \core.registers[16][2] ;
 wire \core.registers[16][30] ;
 wire \core.registers[16][31] ;
 wire \core.registers[16][3] ;
 wire \core.registers[16][4] ;
 wire \core.registers[16][5] ;
 wire \core.registers[16][6] ;
 wire \core.registers[16][7] ;
 wire \core.registers[16][8] ;
 wire \core.registers[16][9] ;
 wire \core.registers[17][0] ;
 wire \core.registers[17][10] ;
 wire \core.registers[17][11] ;
 wire \core.registers[17][12] ;
 wire \core.registers[17][13] ;
 wire \core.registers[17][14] ;
 wire \core.registers[17][15] ;
 wire \core.registers[17][16] ;
 wire \core.registers[17][17] ;
 wire \core.registers[17][18] ;
 wire \core.registers[17][19] ;
 wire \core.registers[17][1] ;
 wire \core.registers[17][20] ;
 wire \core.registers[17][21] ;
 wire \core.registers[17][22] ;
 wire \core.registers[17][23] ;
 wire \core.registers[17][24] ;
 wire \core.registers[17][25] ;
 wire \core.registers[17][26] ;
 wire \core.registers[17][27] ;
 wire \core.registers[17][28] ;
 wire \core.registers[17][29] ;
 wire \core.registers[17][2] ;
 wire \core.registers[17][30] ;
 wire \core.registers[17][31] ;
 wire \core.registers[17][3] ;
 wire \core.registers[17][4] ;
 wire \core.registers[17][5] ;
 wire \core.registers[17][6] ;
 wire \core.registers[17][7] ;
 wire \core.registers[17][8] ;
 wire \core.registers[17][9] ;
 wire \core.registers[18][0] ;
 wire \core.registers[18][10] ;
 wire \core.registers[18][11] ;
 wire \core.registers[18][12] ;
 wire \core.registers[18][13] ;
 wire \core.registers[18][14] ;
 wire \core.registers[18][15] ;
 wire \core.registers[18][16] ;
 wire \core.registers[18][17] ;
 wire \core.registers[18][18] ;
 wire \core.registers[18][19] ;
 wire \core.registers[18][1] ;
 wire \core.registers[18][20] ;
 wire \core.registers[18][21] ;
 wire \core.registers[18][22] ;
 wire \core.registers[18][23] ;
 wire \core.registers[18][24] ;
 wire \core.registers[18][25] ;
 wire \core.registers[18][26] ;
 wire \core.registers[18][27] ;
 wire \core.registers[18][28] ;
 wire \core.registers[18][29] ;
 wire \core.registers[18][2] ;
 wire \core.registers[18][30] ;
 wire \core.registers[18][31] ;
 wire \core.registers[18][3] ;
 wire \core.registers[18][4] ;
 wire \core.registers[18][5] ;
 wire \core.registers[18][6] ;
 wire \core.registers[18][7] ;
 wire \core.registers[18][8] ;
 wire \core.registers[18][9] ;
 wire \core.registers[19][0] ;
 wire \core.registers[19][10] ;
 wire \core.registers[19][11] ;
 wire \core.registers[19][12] ;
 wire \core.registers[19][13] ;
 wire \core.registers[19][14] ;
 wire \core.registers[19][15] ;
 wire \core.registers[19][16] ;
 wire \core.registers[19][17] ;
 wire \core.registers[19][18] ;
 wire \core.registers[19][19] ;
 wire \core.registers[19][1] ;
 wire \core.registers[19][20] ;
 wire \core.registers[19][21] ;
 wire \core.registers[19][22] ;
 wire \core.registers[19][23] ;
 wire \core.registers[19][24] ;
 wire \core.registers[19][25] ;
 wire \core.registers[19][26] ;
 wire \core.registers[19][27] ;
 wire \core.registers[19][28] ;
 wire \core.registers[19][29] ;
 wire \core.registers[19][2] ;
 wire \core.registers[19][30] ;
 wire \core.registers[19][31] ;
 wire \core.registers[19][3] ;
 wire \core.registers[19][4] ;
 wire \core.registers[19][5] ;
 wire \core.registers[19][6] ;
 wire \core.registers[19][7] ;
 wire \core.registers[19][8] ;
 wire \core.registers[19][9] ;
 wire \core.registers[1][0] ;
 wire \core.registers[1][10] ;
 wire \core.registers[1][11] ;
 wire \core.registers[1][12] ;
 wire \core.registers[1][13] ;
 wire \core.registers[1][14] ;
 wire \core.registers[1][15] ;
 wire \core.registers[1][16] ;
 wire \core.registers[1][17] ;
 wire \core.registers[1][18] ;
 wire \core.registers[1][19] ;
 wire \core.registers[1][1] ;
 wire \core.registers[1][20] ;
 wire \core.registers[1][21] ;
 wire \core.registers[1][22] ;
 wire \core.registers[1][23] ;
 wire \core.registers[1][24] ;
 wire \core.registers[1][25] ;
 wire \core.registers[1][26] ;
 wire \core.registers[1][27] ;
 wire \core.registers[1][28] ;
 wire \core.registers[1][29] ;
 wire \core.registers[1][2] ;
 wire \core.registers[1][30] ;
 wire \core.registers[1][31] ;
 wire \core.registers[1][3] ;
 wire \core.registers[1][4] ;
 wire \core.registers[1][5] ;
 wire \core.registers[1][6] ;
 wire \core.registers[1][7] ;
 wire \core.registers[1][8] ;
 wire \core.registers[1][9] ;
 wire \core.registers[20][0] ;
 wire \core.registers[20][10] ;
 wire \core.registers[20][11] ;
 wire \core.registers[20][12] ;
 wire \core.registers[20][13] ;
 wire \core.registers[20][14] ;
 wire \core.registers[20][15] ;
 wire \core.registers[20][16] ;
 wire \core.registers[20][17] ;
 wire \core.registers[20][18] ;
 wire \core.registers[20][19] ;
 wire \core.registers[20][1] ;
 wire \core.registers[20][20] ;
 wire \core.registers[20][21] ;
 wire \core.registers[20][22] ;
 wire \core.registers[20][23] ;
 wire \core.registers[20][24] ;
 wire \core.registers[20][25] ;
 wire \core.registers[20][26] ;
 wire \core.registers[20][27] ;
 wire \core.registers[20][28] ;
 wire \core.registers[20][29] ;
 wire \core.registers[20][2] ;
 wire \core.registers[20][30] ;
 wire \core.registers[20][31] ;
 wire \core.registers[20][3] ;
 wire \core.registers[20][4] ;
 wire \core.registers[20][5] ;
 wire \core.registers[20][6] ;
 wire \core.registers[20][7] ;
 wire \core.registers[20][8] ;
 wire \core.registers[20][9] ;
 wire \core.registers[21][0] ;
 wire \core.registers[21][10] ;
 wire \core.registers[21][11] ;
 wire \core.registers[21][12] ;
 wire \core.registers[21][13] ;
 wire \core.registers[21][14] ;
 wire \core.registers[21][15] ;
 wire \core.registers[21][16] ;
 wire \core.registers[21][17] ;
 wire \core.registers[21][18] ;
 wire \core.registers[21][19] ;
 wire \core.registers[21][1] ;
 wire \core.registers[21][20] ;
 wire \core.registers[21][21] ;
 wire \core.registers[21][22] ;
 wire \core.registers[21][23] ;
 wire \core.registers[21][24] ;
 wire \core.registers[21][25] ;
 wire \core.registers[21][26] ;
 wire \core.registers[21][27] ;
 wire \core.registers[21][28] ;
 wire \core.registers[21][29] ;
 wire \core.registers[21][2] ;
 wire \core.registers[21][30] ;
 wire \core.registers[21][31] ;
 wire \core.registers[21][3] ;
 wire \core.registers[21][4] ;
 wire \core.registers[21][5] ;
 wire \core.registers[21][6] ;
 wire \core.registers[21][7] ;
 wire \core.registers[21][8] ;
 wire \core.registers[21][9] ;
 wire \core.registers[22][0] ;
 wire \core.registers[22][10] ;
 wire \core.registers[22][11] ;
 wire \core.registers[22][12] ;
 wire \core.registers[22][13] ;
 wire \core.registers[22][14] ;
 wire \core.registers[22][15] ;
 wire \core.registers[22][16] ;
 wire \core.registers[22][17] ;
 wire \core.registers[22][18] ;
 wire \core.registers[22][19] ;
 wire \core.registers[22][1] ;
 wire \core.registers[22][20] ;
 wire \core.registers[22][21] ;
 wire \core.registers[22][22] ;
 wire \core.registers[22][23] ;
 wire \core.registers[22][24] ;
 wire \core.registers[22][25] ;
 wire \core.registers[22][26] ;
 wire \core.registers[22][27] ;
 wire \core.registers[22][28] ;
 wire \core.registers[22][29] ;
 wire \core.registers[22][2] ;
 wire \core.registers[22][30] ;
 wire \core.registers[22][31] ;
 wire \core.registers[22][3] ;
 wire \core.registers[22][4] ;
 wire \core.registers[22][5] ;
 wire \core.registers[22][6] ;
 wire \core.registers[22][7] ;
 wire \core.registers[22][8] ;
 wire \core.registers[22][9] ;
 wire \core.registers[23][0] ;
 wire \core.registers[23][10] ;
 wire \core.registers[23][11] ;
 wire \core.registers[23][12] ;
 wire \core.registers[23][13] ;
 wire \core.registers[23][14] ;
 wire \core.registers[23][15] ;
 wire \core.registers[23][16] ;
 wire \core.registers[23][17] ;
 wire \core.registers[23][18] ;
 wire \core.registers[23][19] ;
 wire \core.registers[23][1] ;
 wire \core.registers[23][20] ;
 wire \core.registers[23][21] ;
 wire \core.registers[23][22] ;
 wire \core.registers[23][23] ;
 wire \core.registers[23][24] ;
 wire \core.registers[23][25] ;
 wire \core.registers[23][26] ;
 wire \core.registers[23][27] ;
 wire \core.registers[23][28] ;
 wire \core.registers[23][29] ;
 wire \core.registers[23][2] ;
 wire \core.registers[23][30] ;
 wire \core.registers[23][31] ;
 wire \core.registers[23][3] ;
 wire \core.registers[23][4] ;
 wire \core.registers[23][5] ;
 wire \core.registers[23][6] ;
 wire \core.registers[23][7] ;
 wire \core.registers[23][8] ;
 wire \core.registers[23][9] ;
 wire \core.registers[24][0] ;
 wire \core.registers[24][10] ;
 wire \core.registers[24][11] ;
 wire \core.registers[24][12] ;
 wire \core.registers[24][13] ;
 wire \core.registers[24][14] ;
 wire \core.registers[24][15] ;
 wire \core.registers[24][16] ;
 wire \core.registers[24][17] ;
 wire \core.registers[24][18] ;
 wire \core.registers[24][19] ;
 wire \core.registers[24][1] ;
 wire \core.registers[24][20] ;
 wire \core.registers[24][21] ;
 wire \core.registers[24][22] ;
 wire \core.registers[24][23] ;
 wire \core.registers[24][24] ;
 wire \core.registers[24][25] ;
 wire \core.registers[24][26] ;
 wire \core.registers[24][27] ;
 wire \core.registers[24][28] ;
 wire \core.registers[24][29] ;
 wire \core.registers[24][2] ;
 wire \core.registers[24][30] ;
 wire \core.registers[24][31] ;
 wire \core.registers[24][3] ;
 wire \core.registers[24][4] ;
 wire \core.registers[24][5] ;
 wire \core.registers[24][6] ;
 wire \core.registers[24][7] ;
 wire \core.registers[24][8] ;
 wire \core.registers[24][9] ;
 wire \core.registers[25][0] ;
 wire \core.registers[25][10] ;
 wire \core.registers[25][11] ;
 wire \core.registers[25][12] ;
 wire \core.registers[25][13] ;
 wire \core.registers[25][14] ;
 wire \core.registers[25][15] ;
 wire \core.registers[25][16] ;
 wire \core.registers[25][17] ;
 wire \core.registers[25][18] ;
 wire \core.registers[25][19] ;
 wire \core.registers[25][1] ;
 wire \core.registers[25][20] ;
 wire \core.registers[25][21] ;
 wire \core.registers[25][22] ;
 wire \core.registers[25][23] ;
 wire \core.registers[25][24] ;
 wire \core.registers[25][25] ;
 wire \core.registers[25][26] ;
 wire \core.registers[25][27] ;
 wire \core.registers[25][28] ;
 wire \core.registers[25][29] ;
 wire \core.registers[25][2] ;
 wire \core.registers[25][30] ;
 wire \core.registers[25][31] ;
 wire \core.registers[25][3] ;
 wire \core.registers[25][4] ;
 wire \core.registers[25][5] ;
 wire \core.registers[25][6] ;
 wire \core.registers[25][7] ;
 wire \core.registers[25][8] ;
 wire \core.registers[25][9] ;
 wire \core.registers[26][0] ;
 wire \core.registers[26][10] ;
 wire \core.registers[26][11] ;
 wire \core.registers[26][12] ;
 wire \core.registers[26][13] ;
 wire \core.registers[26][14] ;
 wire \core.registers[26][15] ;
 wire \core.registers[26][16] ;
 wire \core.registers[26][17] ;
 wire \core.registers[26][18] ;
 wire \core.registers[26][19] ;
 wire \core.registers[26][1] ;
 wire \core.registers[26][20] ;
 wire \core.registers[26][21] ;
 wire \core.registers[26][22] ;
 wire \core.registers[26][23] ;
 wire \core.registers[26][24] ;
 wire \core.registers[26][25] ;
 wire \core.registers[26][26] ;
 wire \core.registers[26][27] ;
 wire \core.registers[26][28] ;
 wire \core.registers[26][29] ;
 wire \core.registers[26][2] ;
 wire \core.registers[26][30] ;
 wire \core.registers[26][31] ;
 wire \core.registers[26][3] ;
 wire \core.registers[26][4] ;
 wire \core.registers[26][5] ;
 wire \core.registers[26][6] ;
 wire \core.registers[26][7] ;
 wire \core.registers[26][8] ;
 wire \core.registers[26][9] ;
 wire \core.registers[27][0] ;
 wire \core.registers[27][10] ;
 wire \core.registers[27][11] ;
 wire \core.registers[27][12] ;
 wire \core.registers[27][13] ;
 wire \core.registers[27][14] ;
 wire \core.registers[27][15] ;
 wire \core.registers[27][16] ;
 wire \core.registers[27][17] ;
 wire \core.registers[27][18] ;
 wire \core.registers[27][19] ;
 wire \core.registers[27][1] ;
 wire \core.registers[27][20] ;
 wire \core.registers[27][21] ;
 wire \core.registers[27][22] ;
 wire \core.registers[27][23] ;
 wire \core.registers[27][24] ;
 wire \core.registers[27][25] ;
 wire \core.registers[27][26] ;
 wire \core.registers[27][27] ;
 wire \core.registers[27][28] ;
 wire \core.registers[27][29] ;
 wire \core.registers[27][2] ;
 wire \core.registers[27][30] ;
 wire \core.registers[27][31] ;
 wire \core.registers[27][3] ;
 wire \core.registers[27][4] ;
 wire \core.registers[27][5] ;
 wire \core.registers[27][6] ;
 wire \core.registers[27][7] ;
 wire \core.registers[27][8] ;
 wire \core.registers[27][9] ;
 wire \core.registers[28][0] ;
 wire \core.registers[28][10] ;
 wire \core.registers[28][11] ;
 wire \core.registers[28][12] ;
 wire \core.registers[28][13] ;
 wire \core.registers[28][14] ;
 wire \core.registers[28][15] ;
 wire \core.registers[28][16] ;
 wire \core.registers[28][17] ;
 wire \core.registers[28][18] ;
 wire \core.registers[28][19] ;
 wire \core.registers[28][1] ;
 wire \core.registers[28][20] ;
 wire \core.registers[28][21] ;
 wire \core.registers[28][22] ;
 wire \core.registers[28][23] ;
 wire \core.registers[28][24] ;
 wire \core.registers[28][25] ;
 wire \core.registers[28][26] ;
 wire \core.registers[28][27] ;
 wire \core.registers[28][28] ;
 wire \core.registers[28][29] ;
 wire \core.registers[28][2] ;
 wire \core.registers[28][30] ;
 wire \core.registers[28][31] ;
 wire \core.registers[28][3] ;
 wire \core.registers[28][4] ;
 wire \core.registers[28][5] ;
 wire \core.registers[28][6] ;
 wire \core.registers[28][7] ;
 wire \core.registers[28][8] ;
 wire \core.registers[28][9] ;
 wire \core.registers[29][0] ;
 wire \core.registers[29][10] ;
 wire \core.registers[29][11] ;
 wire \core.registers[29][12] ;
 wire \core.registers[29][13] ;
 wire \core.registers[29][14] ;
 wire \core.registers[29][15] ;
 wire \core.registers[29][16] ;
 wire \core.registers[29][17] ;
 wire \core.registers[29][18] ;
 wire \core.registers[29][19] ;
 wire \core.registers[29][1] ;
 wire \core.registers[29][20] ;
 wire \core.registers[29][21] ;
 wire \core.registers[29][22] ;
 wire \core.registers[29][23] ;
 wire \core.registers[29][24] ;
 wire \core.registers[29][25] ;
 wire \core.registers[29][26] ;
 wire \core.registers[29][27] ;
 wire \core.registers[29][28] ;
 wire \core.registers[29][29] ;
 wire \core.registers[29][2] ;
 wire \core.registers[29][30] ;
 wire \core.registers[29][31] ;
 wire \core.registers[29][3] ;
 wire \core.registers[29][4] ;
 wire \core.registers[29][5] ;
 wire \core.registers[29][6] ;
 wire \core.registers[29][7] ;
 wire \core.registers[29][8] ;
 wire \core.registers[29][9] ;
 wire \core.registers[2][0] ;
 wire \core.registers[2][10] ;
 wire \core.registers[2][11] ;
 wire \core.registers[2][12] ;
 wire \core.registers[2][13] ;
 wire \core.registers[2][14] ;
 wire \core.registers[2][15] ;
 wire \core.registers[2][16] ;
 wire \core.registers[2][17] ;
 wire \core.registers[2][18] ;
 wire \core.registers[2][19] ;
 wire \core.registers[2][1] ;
 wire \core.registers[2][20] ;
 wire \core.registers[2][21] ;
 wire \core.registers[2][22] ;
 wire \core.registers[2][23] ;
 wire \core.registers[2][24] ;
 wire \core.registers[2][25] ;
 wire \core.registers[2][26] ;
 wire \core.registers[2][27] ;
 wire \core.registers[2][28] ;
 wire \core.registers[2][29] ;
 wire \core.registers[2][2] ;
 wire \core.registers[2][30] ;
 wire \core.registers[2][31] ;
 wire \core.registers[2][3] ;
 wire \core.registers[2][4] ;
 wire \core.registers[2][5] ;
 wire \core.registers[2][6] ;
 wire \core.registers[2][7] ;
 wire \core.registers[2][8] ;
 wire \core.registers[2][9] ;
 wire \core.registers[30][0] ;
 wire \core.registers[30][10] ;
 wire \core.registers[30][11] ;
 wire \core.registers[30][12] ;
 wire \core.registers[30][13] ;
 wire \core.registers[30][14] ;
 wire \core.registers[30][15] ;
 wire \core.registers[30][16] ;
 wire \core.registers[30][17] ;
 wire \core.registers[30][18] ;
 wire \core.registers[30][19] ;
 wire \core.registers[30][1] ;
 wire \core.registers[30][20] ;
 wire \core.registers[30][21] ;
 wire \core.registers[30][22] ;
 wire \core.registers[30][23] ;
 wire \core.registers[30][24] ;
 wire \core.registers[30][25] ;
 wire \core.registers[30][26] ;
 wire \core.registers[30][27] ;
 wire \core.registers[30][28] ;
 wire \core.registers[30][29] ;
 wire \core.registers[30][2] ;
 wire \core.registers[30][30] ;
 wire \core.registers[30][31] ;
 wire \core.registers[30][3] ;
 wire \core.registers[30][4] ;
 wire \core.registers[30][5] ;
 wire \core.registers[30][6] ;
 wire \core.registers[30][7] ;
 wire \core.registers[30][8] ;
 wire \core.registers[30][9] ;
 wire \core.registers[31][0] ;
 wire \core.registers[31][10] ;
 wire \core.registers[31][11] ;
 wire \core.registers[31][12] ;
 wire \core.registers[31][13] ;
 wire \core.registers[31][14] ;
 wire \core.registers[31][15] ;
 wire \core.registers[31][16] ;
 wire \core.registers[31][17] ;
 wire \core.registers[31][18] ;
 wire \core.registers[31][19] ;
 wire \core.registers[31][1] ;
 wire \core.registers[31][20] ;
 wire \core.registers[31][21] ;
 wire \core.registers[31][22] ;
 wire \core.registers[31][23] ;
 wire \core.registers[31][24] ;
 wire \core.registers[31][25] ;
 wire \core.registers[31][26] ;
 wire \core.registers[31][27] ;
 wire \core.registers[31][28] ;
 wire \core.registers[31][29] ;
 wire \core.registers[31][2] ;
 wire \core.registers[31][30] ;
 wire \core.registers[31][31] ;
 wire \core.registers[31][3] ;
 wire \core.registers[31][4] ;
 wire \core.registers[31][5] ;
 wire \core.registers[31][6] ;
 wire \core.registers[31][7] ;
 wire \core.registers[31][8] ;
 wire \core.registers[31][9] ;
 wire \core.registers[3][0] ;
 wire \core.registers[3][10] ;
 wire \core.registers[3][11] ;
 wire \core.registers[3][12] ;
 wire \core.registers[3][13] ;
 wire \core.registers[3][14] ;
 wire \core.registers[3][15] ;
 wire \core.registers[3][16] ;
 wire \core.registers[3][17] ;
 wire \core.registers[3][18] ;
 wire \core.registers[3][19] ;
 wire \core.registers[3][1] ;
 wire \core.registers[3][20] ;
 wire \core.registers[3][21] ;
 wire \core.registers[3][22] ;
 wire \core.registers[3][23] ;
 wire \core.registers[3][24] ;
 wire \core.registers[3][25] ;
 wire \core.registers[3][26] ;
 wire \core.registers[3][27] ;
 wire \core.registers[3][28] ;
 wire \core.registers[3][29] ;
 wire \core.registers[3][2] ;
 wire \core.registers[3][30] ;
 wire \core.registers[3][31] ;
 wire \core.registers[3][3] ;
 wire \core.registers[3][4] ;
 wire \core.registers[3][5] ;
 wire \core.registers[3][6] ;
 wire \core.registers[3][7] ;
 wire \core.registers[3][8] ;
 wire \core.registers[3][9] ;
 wire \core.registers[4][0] ;
 wire \core.registers[4][10] ;
 wire \core.registers[4][11] ;
 wire \core.registers[4][12] ;
 wire \core.registers[4][13] ;
 wire \core.registers[4][14] ;
 wire \core.registers[4][15] ;
 wire \core.registers[4][16] ;
 wire \core.registers[4][17] ;
 wire \core.registers[4][18] ;
 wire \core.registers[4][19] ;
 wire \core.registers[4][1] ;
 wire \core.registers[4][20] ;
 wire \core.registers[4][21] ;
 wire \core.registers[4][22] ;
 wire \core.registers[4][23] ;
 wire \core.registers[4][24] ;
 wire \core.registers[4][25] ;
 wire \core.registers[4][26] ;
 wire \core.registers[4][27] ;
 wire \core.registers[4][28] ;
 wire \core.registers[4][29] ;
 wire \core.registers[4][2] ;
 wire \core.registers[4][30] ;
 wire \core.registers[4][31] ;
 wire \core.registers[4][3] ;
 wire \core.registers[4][4] ;
 wire \core.registers[4][5] ;
 wire \core.registers[4][6] ;
 wire \core.registers[4][7] ;
 wire \core.registers[4][8] ;
 wire \core.registers[4][9] ;
 wire \core.registers[5][0] ;
 wire \core.registers[5][10] ;
 wire \core.registers[5][11] ;
 wire \core.registers[5][12] ;
 wire \core.registers[5][13] ;
 wire \core.registers[5][14] ;
 wire \core.registers[5][15] ;
 wire \core.registers[5][16] ;
 wire \core.registers[5][17] ;
 wire \core.registers[5][18] ;
 wire \core.registers[5][19] ;
 wire \core.registers[5][1] ;
 wire \core.registers[5][20] ;
 wire \core.registers[5][21] ;
 wire \core.registers[5][22] ;
 wire \core.registers[5][23] ;
 wire \core.registers[5][24] ;
 wire \core.registers[5][25] ;
 wire \core.registers[5][26] ;
 wire \core.registers[5][27] ;
 wire \core.registers[5][28] ;
 wire \core.registers[5][29] ;
 wire \core.registers[5][2] ;
 wire \core.registers[5][30] ;
 wire \core.registers[5][31] ;
 wire \core.registers[5][3] ;
 wire \core.registers[5][4] ;
 wire \core.registers[5][5] ;
 wire \core.registers[5][6] ;
 wire \core.registers[5][7] ;
 wire \core.registers[5][8] ;
 wire \core.registers[5][9] ;
 wire \core.registers[6][0] ;
 wire \core.registers[6][10] ;
 wire \core.registers[6][11] ;
 wire \core.registers[6][12] ;
 wire \core.registers[6][13] ;
 wire \core.registers[6][14] ;
 wire \core.registers[6][15] ;
 wire \core.registers[6][16] ;
 wire \core.registers[6][17] ;
 wire \core.registers[6][18] ;
 wire \core.registers[6][19] ;
 wire \core.registers[6][1] ;
 wire \core.registers[6][20] ;
 wire \core.registers[6][21] ;
 wire \core.registers[6][22] ;
 wire \core.registers[6][23] ;
 wire \core.registers[6][24] ;
 wire \core.registers[6][25] ;
 wire \core.registers[6][26] ;
 wire \core.registers[6][27] ;
 wire \core.registers[6][28] ;
 wire \core.registers[6][29] ;
 wire \core.registers[6][2] ;
 wire \core.registers[6][30] ;
 wire \core.registers[6][31] ;
 wire \core.registers[6][3] ;
 wire \core.registers[6][4] ;
 wire \core.registers[6][5] ;
 wire \core.registers[6][6] ;
 wire \core.registers[6][7] ;
 wire \core.registers[6][8] ;
 wire \core.registers[6][9] ;
 wire \core.registers[7][0] ;
 wire \core.registers[7][10] ;
 wire \core.registers[7][11] ;
 wire \core.registers[7][12] ;
 wire \core.registers[7][13] ;
 wire \core.registers[7][14] ;
 wire \core.registers[7][15] ;
 wire \core.registers[7][16] ;
 wire \core.registers[7][17] ;
 wire \core.registers[7][18] ;
 wire \core.registers[7][19] ;
 wire \core.registers[7][1] ;
 wire \core.registers[7][20] ;
 wire \core.registers[7][21] ;
 wire \core.registers[7][22] ;
 wire \core.registers[7][23] ;
 wire \core.registers[7][24] ;
 wire \core.registers[7][25] ;
 wire \core.registers[7][26] ;
 wire \core.registers[7][27] ;
 wire \core.registers[7][28] ;
 wire \core.registers[7][29] ;
 wire \core.registers[7][2] ;
 wire \core.registers[7][30] ;
 wire \core.registers[7][31] ;
 wire \core.registers[7][3] ;
 wire \core.registers[7][4] ;
 wire \core.registers[7][5] ;
 wire \core.registers[7][6] ;
 wire \core.registers[7][7] ;
 wire \core.registers[7][8] ;
 wire \core.registers[7][9] ;
 wire \core.registers[8][0] ;
 wire \core.registers[8][10] ;
 wire \core.registers[8][11] ;
 wire \core.registers[8][12] ;
 wire \core.registers[8][13] ;
 wire \core.registers[8][14] ;
 wire \core.registers[8][15] ;
 wire \core.registers[8][16] ;
 wire \core.registers[8][17] ;
 wire \core.registers[8][18] ;
 wire \core.registers[8][19] ;
 wire \core.registers[8][1] ;
 wire \core.registers[8][20] ;
 wire \core.registers[8][21] ;
 wire \core.registers[8][22] ;
 wire \core.registers[8][23] ;
 wire \core.registers[8][24] ;
 wire \core.registers[8][25] ;
 wire \core.registers[8][26] ;
 wire \core.registers[8][27] ;
 wire \core.registers[8][28] ;
 wire \core.registers[8][29] ;
 wire \core.registers[8][2] ;
 wire \core.registers[8][30] ;
 wire \core.registers[8][31] ;
 wire \core.registers[8][3] ;
 wire \core.registers[8][4] ;
 wire \core.registers[8][5] ;
 wire \core.registers[8][6] ;
 wire \core.registers[8][7] ;
 wire \core.registers[8][8] ;
 wire \core.registers[8][9] ;
 wire \core.registers[9][0] ;
 wire \core.registers[9][10] ;
 wire \core.registers[9][11] ;
 wire \core.registers[9][12] ;
 wire \core.registers[9][13] ;
 wire \core.registers[9][14] ;
 wire \core.registers[9][15] ;
 wire \core.registers[9][16] ;
 wire \core.registers[9][17] ;
 wire \core.registers[9][18] ;
 wire \core.registers[9][19] ;
 wire \core.registers[9][1] ;
 wire \core.registers[9][20] ;
 wire \core.registers[9][21] ;
 wire \core.registers[9][22] ;
 wire \core.registers[9][23] ;
 wire \core.registers[9][24] ;
 wire \core.registers[9][25] ;
 wire \core.registers[9][26] ;
 wire \core.registers[9][27] ;
 wire \core.registers[9][28] ;
 wire \core.registers[9][29] ;
 wire \core.registers[9][2] ;
 wire \core.registers[9][30] ;
 wire \core.registers[9][31] ;
 wire \core.registers[9][3] ;
 wire \core.registers[9][4] ;
 wire \core.registers[9][5] ;
 wire \core.registers[9][6] ;
 wire \core.registers[9][7] ;
 wire \core.registers[9][8] ;
 wire \core.registers[9][9] ;
 wire \coreManagement.control[1] ;
 wire \coreWBInterface.readDataBuffered[0] ;
 wire \coreWBInterface.readDataBuffered[10] ;
 wire \coreWBInterface.readDataBuffered[11] ;
 wire \coreWBInterface.readDataBuffered[12] ;
 wire \coreWBInterface.readDataBuffered[13] ;
 wire \coreWBInterface.readDataBuffered[14] ;
 wire \coreWBInterface.readDataBuffered[15] ;
 wire \coreWBInterface.readDataBuffered[16] ;
 wire \coreWBInterface.readDataBuffered[17] ;
 wire \coreWBInterface.readDataBuffered[18] ;
 wire \coreWBInterface.readDataBuffered[19] ;
 wire \coreWBInterface.readDataBuffered[1] ;
 wire \coreWBInterface.readDataBuffered[20] ;
 wire \coreWBInterface.readDataBuffered[21] ;
 wire \coreWBInterface.readDataBuffered[22] ;
 wire \coreWBInterface.readDataBuffered[23] ;
 wire \coreWBInterface.readDataBuffered[24] ;
 wire \coreWBInterface.readDataBuffered[25] ;
 wire \coreWBInterface.readDataBuffered[26] ;
 wire \coreWBInterface.readDataBuffered[27] ;
 wire \coreWBInterface.readDataBuffered[28] ;
 wire \coreWBInterface.readDataBuffered[29] ;
 wire \coreWBInterface.readDataBuffered[2] ;
 wire \coreWBInterface.readDataBuffered[30] ;
 wire \coreWBInterface.readDataBuffered[31] ;
 wire \coreWBInterface.readDataBuffered[3] ;
 wire \coreWBInterface.readDataBuffered[4] ;
 wire \coreWBInterface.readDataBuffered[5] ;
 wire \coreWBInterface.readDataBuffered[6] ;
 wire \coreWBInterface.readDataBuffered[7] ;
 wire \coreWBInterface.readDataBuffered[8] ;
 wire \coreWBInterface.readDataBuffered[9] ;
 wire \coreWBInterface.state[0] ;
 wire \coreWBInterface.state[1] ;
 wire \jtag.dataBSRRegister.data[0] ;
 wire \jtag.dataBSRRegister.data[10] ;
 wire \jtag.dataBSRRegister.data[11] ;
 wire \jtag.dataBSRRegister.data[12] ;
 wire \jtag.dataBSRRegister.data[13] ;
 wire \jtag.dataBSRRegister.data[14] ;
 wire \jtag.dataBSRRegister.data[15] ;
 wire \jtag.dataBSRRegister.data[16] ;
 wire \jtag.dataBSRRegister.data[17] ;
 wire \jtag.dataBSRRegister.data[18] ;
 wire \jtag.dataBSRRegister.data[19] ;
 wire \jtag.dataBSRRegister.data[1] ;
 wire \jtag.dataBSRRegister.data[20] ;
 wire \jtag.dataBSRRegister.data[21] ;
 wire \jtag.dataBSRRegister.data[22] ;
 wire \jtag.dataBSRRegister.data[23] ;
 wire \jtag.dataBSRRegister.data[24] ;
 wire \jtag.dataBSRRegister.data[25] ;
 wire \jtag.dataBSRRegister.data[26] ;
 wire \jtag.dataBSRRegister.data[27] ;
 wire \jtag.dataBSRRegister.data[28] ;
 wire \jtag.dataBSRRegister.data[29] ;
 wire \jtag.dataBSRRegister.data[2] ;
 wire \jtag.dataBSRRegister.data[30] ;
 wire \jtag.dataBSRRegister.data[31] ;
 wire \jtag.dataBSRRegister.data[3] ;
 wire \jtag.dataBSRRegister.data[4] ;
 wire \jtag.dataBSRRegister.data[5] ;
 wire \jtag.dataBSRRegister.data[6] ;
 wire \jtag.dataBSRRegister.data[7] ;
 wire \jtag.dataBSRRegister.data[8] ;
 wire \jtag.dataBSRRegister.data[9] ;
 wire \jtag.dataBypassRegister.data ;
 wire \jtag.dataIDRegister.data[0] ;
 wire \jtag.dataIDRegister.data[10] ;
 wire \jtag.dataIDRegister.data[11] ;
 wire \jtag.dataIDRegister.data[12] ;
 wire \jtag.dataIDRegister.data[13] ;
 wire \jtag.dataIDRegister.data[14] ;
 wire \jtag.dataIDRegister.data[15] ;
 wire \jtag.dataIDRegister.data[16] ;
 wire \jtag.dataIDRegister.data[17] ;
 wire \jtag.dataIDRegister.data[18] ;
 wire \jtag.dataIDRegister.data[19] ;
 wire \jtag.dataIDRegister.data[1] ;
 wire \jtag.dataIDRegister.data[20] ;
 wire \jtag.dataIDRegister.data[21] ;
 wire \jtag.dataIDRegister.data[22] ;
 wire \jtag.dataIDRegister.data[23] ;
 wire \jtag.dataIDRegister.data[24] ;
 wire \jtag.dataIDRegister.data[25] ;
 wire \jtag.dataIDRegister.data[26] ;
 wire \jtag.dataIDRegister.data[27] ;
 wire \jtag.dataIDRegister.data[28] ;
 wire \jtag.dataIDRegister.data[29] ;
 wire \jtag.dataIDRegister.data[2] ;
 wire \jtag.dataIDRegister.data[30] ;
 wire \jtag.dataIDRegister.data[31] ;
 wire \jtag.dataIDRegister.data[3] ;
 wire \jtag.dataIDRegister.data[4] ;
 wire \jtag.dataIDRegister.data[5] ;
 wire \jtag.dataIDRegister.data[6] ;
 wire \jtag.dataIDRegister.data[7] ;
 wire \jtag.dataIDRegister.data[8] ;
 wire \jtag.dataIDRegister.data[9] ;
 wire \jtag.instructionRegister.data[0] ;
 wire \jtag.instructionRegister.data[1] ;
 wire \jtag.instructionRegister.data[2] ;
 wire \jtag.instructionRegister.data[3] ;
 wire \jtag.instructionRegister.data[4] ;
 wire \jtag.managementAddress[0] ;
 wire \jtag.managementAddress[10] ;
 wire \jtag.managementAddress[11] ;
 wire \jtag.managementAddress[12] ;
 wire \jtag.managementAddress[13] ;
 wire \jtag.managementAddress[14] ;
 wire \jtag.managementAddress[15] ;
 wire \jtag.managementAddress[16] ;
 wire \jtag.managementAddress[17] ;
 wire \jtag.managementAddress[18] ;
 wire \jtag.managementAddress[19] ;
 wire \jtag.managementAddress[1] ;
 wire \jtag.managementAddress[2] ;
 wire \jtag.managementAddress[3] ;
 wire \jtag.managementAddress[4] ;
 wire \jtag.managementAddress[5] ;
 wire \jtag.managementAddress[6] ;
 wire \jtag.managementAddress[7] ;
 wire \jtag.managementAddress[8] ;
 wire \jtag.managementAddress[9] ;
 wire \jtag.managementReadData[0] ;
 wire \jtag.managementReadData[10] ;
 wire \jtag.managementReadData[11] ;
 wire \jtag.managementReadData[12] ;
 wire \jtag.managementReadData[13] ;
 wire \jtag.managementReadData[14] ;
 wire \jtag.managementReadData[15] ;
 wire \jtag.managementReadData[16] ;
 wire \jtag.managementReadData[17] ;
 wire \jtag.managementReadData[18] ;
 wire \jtag.managementReadData[19] ;
 wire \jtag.managementReadData[1] ;
 wire \jtag.managementReadData[20] ;
 wire \jtag.managementReadData[21] ;
 wire \jtag.managementReadData[22] ;
 wire \jtag.managementReadData[23] ;
 wire \jtag.managementReadData[24] ;
 wire \jtag.managementReadData[25] ;
 wire \jtag.managementReadData[26] ;
 wire \jtag.managementReadData[27] ;
 wire \jtag.managementReadData[28] ;
 wire \jtag.managementReadData[29] ;
 wire \jtag.managementReadData[2] ;
 wire \jtag.managementReadData[30] ;
 wire \jtag.managementReadData[31] ;
 wire \jtag.managementReadData[3] ;
 wire \jtag.managementReadData[4] ;
 wire \jtag.managementReadData[5] ;
 wire \jtag.managementReadData[6] ;
 wire \jtag.managementReadData[7] ;
 wire \jtag.managementReadData[8] ;
 wire \jtag.managementReadData[9] ;
 wire \jtag.managementState[0] ;
 wire \jtag.managementState[1] ;
 wire \jtag.managementState[2] ;
 wire \jtag.state[0] ;
 wire \jtag.state[1] ;
 wire \jtag.state[2] ;
 wire \jtag.state[3] ;
 wire \jtag.tckRisingEdge ;
 wire \jtag.tckState ;
 wire \localMemoryInterface.coreReadReady ;
 wire \localMemoryInterface.lastCoreByteSelect[0] ;
 wire \localMemoryInterface.lastCoreByteSelect[1] ;
 wire \localMemoryInterface.lastCoreByteSelect[2] ;
 wire \localMemoryInterface.lastCoreByteSelect[3] ;
 wire \localMemoryInterface.lastRBankSelect ;
 wire \localMemoryInterface.lastRWBankSelect ;
 wire \localMemoryInterface.lastWBByteSelect[0] ;
 wire \localMemoryInterface.lastWBByteSelect[1] ;
 wire \localMemoryInterface.lastWBByteSelect[2] ;
 wire \localMemoryInterface.lastWBByteSelect[3] ;
 wire \localMemoryInterface.wbReadReady ;
 wire \memoryController.last_data_enableLocalMemory ;
 wire \memoryController.last_data_enableWB ;
 wire \memoryController.last_instruction_enableLocalMemory ;
 wire \memoryController.last_instruction_enableWB ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \wbSRAMInterface.currentAddress[0] ;
 wire \wbSRAMInterface.currentAddress[10] ;
 wire \wbSRAMInterface.currentAddress[11] ;
 wire \wbSRAMInterface.currentAddress[12] ;
 wire \wbSRAMInterface.currentAddress[13] ;
 wire \wbSRAMInterface.currentAddress[14] ;
 wire \wbSRAMInterface.currentAddress[15] ;
 wire \wbSRAMInterface.currentAddress[16] ;
 wire \wbSRAMInterface.currentAddress[17] ;
 wire \wbSRAMInterface.currentAddress[18] ;
 wire \wbSRAMInterface.currentAddress[19] ;
 wire \wbSRAMInterface.currentAddress[1] ;
 wire \wbSRAMInterface.currentAddress[20] ;
 wire \wbSRAMInterface.currentAddress[21] ;
 wire \wbSRAMInterface.currentAddress[22] ;
 wire \wbSRAMInterface.currentAddress[23] ;
 wire \wbSRAMInterface.currentAddress[2] ;
 wire \wbSRAMInterface.currentAddress[3] ;
 wire \wbSRAMInterface.currentAddress[4] ;
 wire \wbSRAMInterface.currentAddress[5] ;
 wire \wbSRAMInterface.currentAddress[6] ;
 wire \wbSRAMInterface.currentAddress[7] ;
 wire \wbSRAMInterface.currentAddress[8] ;
 wire \wbSRAMInterface.currentAddress[9] ;
 wire \wbSRAMInterface.currentByteSelect[0] ;
 wire \wbSRAMInterface.currentByteSelect[1] ;
 wire \wbSRAMInterface.currentByteSelect[2] ;
 wire \wbSRAMInterface.currentByteSelect[3] ;
 wire \wbSRAMInterface.state[0] ;
 wire \wbSRAMInterface.state[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_00770_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_06704_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_06704_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_06716_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_01944_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_06732_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_06740_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_06740_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_06740_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_02052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(_06740_));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_06740_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_06740_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_02061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(_06771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_06771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_06771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_02081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_06771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_06787_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(_06796_));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(_06796_));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(_06796_));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(_06796_));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(_06796_));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_06796_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_06796_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_06796_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(_06837_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(_06837_));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(_07163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(_07163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(_07484_));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(_07648_));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(_07721_));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(_07746_));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(_07812_));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(_07836_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(_07939_));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(_07977_));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(_08021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(_08034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(_08069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(_08069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(_08131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(_08198_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(_08211_));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(_08230_));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(_08243_));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(_08275_));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(_08294_));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(_08339_));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(_08339_));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(_08357_));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(_08388_));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(_08401_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(_08401_));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(_08419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(_08463_));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(_08529_));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(_08546_));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(_08559_));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(_08559_));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_02163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(_08624_));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(_08624_));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(_08702_));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(_08702_));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(\core.csr.currentInstruction[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(\core.fetchProgramCounter[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(\core.fetchProgramCounter[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(\core.fetchProgramCounter[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(\core.fetchProgramCounter[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(\core.fetchProgramCounter[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(\core.fetchProgramCounter[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(\core.fetchProgramCounter[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(\core.pipe0_currentInstruction[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(\core.pipe0_currentInstruction[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(\core.pipe0_currentInstruction[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(\core.pipe0_currentInstruction[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(\core.pipe0_currentInstruction[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(\core.pipe0_currentInstruction[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(\core.pipe0_currentInstruction[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(\core.registers[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(\core.registers[0][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(\core.registers[0][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(\core.registers[0][29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(\coreWBInterface.readDataBuffered[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(\coreWBInterface.readDataBuffered[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(\coreWBInterface.readDataBuffered[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(\coreWBInterface.readDataBuffered[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(\coreWBInterface.readDataBuffered[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(\coreWBInterface.readDataBuffered[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(\coreWBInterface.readDataBuffered[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_02199_));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(\coreWBInterface.readDataBuffered[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(\coreWBInterface.readDataBuffered[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(\coreWBInterface.readDataBuffered[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(\coreWBInterface.readDataBuffered[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(\coreWBInterface.readDataBuffered[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(\coreWBInterface.readDataBuffered[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(\coreWBInterface.readDataBuffered[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(\coreWBInterface.readDataBuffered[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(\coreWBInterface.readDataBuffered[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(\coreWBInterface.readDataBuffered[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(\coreWBInterface.readDataBuffered[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(\coreWBInterface.readDataBuffered[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(\coreWBInterface.readDataBuffered[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(\coreWBInterface.readDataBuffered[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(\coreWBInterface.readDataBuffered[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(\jtag.dataBSRRegister.data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(\jtag.dataBSRRegister.data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(\jtag.tckRisingEdge ));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(\jtag.tckRisingEdge ));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(\wbSRAMInterface.currentAddress[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(\wbSRAMInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(\wbSRAMInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_03333_));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_00440_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_03375_));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_03421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(net1592));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(net1669));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(net1684));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(net1705));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(net1709));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(net1711));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(net1719));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(net1719));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(net1719));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(net1719));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(net1751));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(net1755));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(net1767));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(net1771));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(net1780));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(net1780));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(net1782));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(net1784));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(net1799));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(net1904));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(net1906));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(_01935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(_02025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(_02099_));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(_02179_));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(_02208_));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(_03369_));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(_03369_));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(_03420_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(_03592_));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(_04720_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_00441_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(_04720_));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(_04726_));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_407 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_408 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_409 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA_410 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_411 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_412 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_413 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_414 (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA_415 (.DIODE(_05737_));
 sky130_fd_sc_hd__diode_2 ANTENNA_416 (.DIODE(_05737_));
 sky130_fd_sc_hd__diode_2 ANTENNA_417 (.DIODE(_06012_));
 sky130_fd_sc_hd__diode_2 ANTENNA_418 (.DIODE(_06506_));
 sky130_fd_sc_hd__diode_2 ANTENNA_419 (.DIODE(_06506_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA_420 (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_421 (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_422 (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA_423 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_424 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_425 (.DIODE(_06760_));
 sky130_fd_sc_hd__diode_2 ANTENNA_426 (.DIODE(_06760_));
 sky130_fd_sc_hd__diode_2 ANTENNA_427 (.DIODE(_06760_));
 sky130_fd_sc_hd__diode_2 ANTENNA_428 (.DIODE(_06771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_429 (.DIODE(_06771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA_430 (.DIODE(_06771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_431 (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA_432 (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA_433 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA_434 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA_435 (.DIODE(_07252_));
 sky130_fd_sc_hd__diode_2 ANTENNA_436 (.DIODE(_07564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_437 (.DIODE(_07716_));
 sky130_fd_sc_hd__diode_2 ANTENNA_438 (.DIODE(_07771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_439 (.DIODE(_07792_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA_440 (.DIODE(_07851_));
 sky130_fd_sc_hd__diode_2 ANTENNA_441 (.DIODE(_07977_));
 sky130_fd_sc_hd__diode_2 ANTENNA_442 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA_443 (.DIODE(_08034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_444 (.DIODE(_08163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_445 (.DIODE(_08189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_446 (.DIODE(_08189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_447 (.DIODE(_08211_));
 sky130_fd_sc_hd__diode_2 ANTENNA_448 (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA_449 (.DIODE(_08434_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA_450 (.DIODE(_08463_));
 sky130_fd_sc_hd__diode_2 ANTENNA_451 (.DIODE(_08484_));
 sky130_fd_sc_hd__diode_2 ANTENNA_452 (.DIODE(_08814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_453 (.DIODE(\core.csr.currentInstruction[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_454 (.DIODE(\core.csr.traps.mie.currentValue[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_455 (.DIODE(\core.fetchProgramCounter[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_456 (.DIODE(\core.fetchProgramCounter[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_457 (.DIODE(\core.fetchProgramCounter[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_458 (.DIODE(\core.fetchProgramCounter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_459 (.DIODE(\core.registers[0][20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA_460 (.DIODE(\coreWBInterface.readDataBuffered[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_461 (.DIODE(\coreWBInterface.readDataBuffered[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_462 (.DIODE(\coreWBInterface.readDataBuffered[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_463 (.DIODE(\coreWBInterface.readDataBuffered[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_464 (.DIODE(\coreWBInterface.readDataBuffered[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_465 (.DIODE(\coreWBInterface.readDataBuffered[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_466 (.DIODE(\coreWBInterface.readDataBuffered[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_467 (.DIODE(\coreWBInterface.readDataBuffered[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_468 (.DIODE(\coreWBInterface.readDataBuffered[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_469 (.DIODE(\coreWBInterface.readDataBuffered[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA_470 (.DIODE(\coreWBInterface.readDataBuffered[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_471 (.DIODE(\jtag.tckRisingEdge ));
 sky130_fd_sc_hd__diode_2 ANTENNA_472 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_473 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_474 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_475 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_476 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_477 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_478 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_479 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA_480 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_481 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_482 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_483 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_484 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_485 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_486 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_487 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_488 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_489 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA_490 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_491 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_492 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_493 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_494 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_495 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_496 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_497 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_498 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_499 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA_500 (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA_501 (.DIODE(net1764));
 sky130_fd_sc_hd__diode_2 ANTENNA_502 (.DIODE(net1767));
 sky130_fd_sc_hd__diode_2 ANTENNA_503 (.DIODE(net1776));
 sky130_fd_sc_hd__diode_2 ANTENNA_504 (.DIODE(net1776));
 sky130_fd_sc_hd__diode_2 ANTENNA_505 (.DIODE(net1784));
 sky130_fd_sc_hd__diode_2 ANTENNA_506 (.DIODE(net1879));
 sky130_fd_sc_hd__diode_2 ANTENNA_507 (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA_508 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_509 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA_510 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_511 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_512 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_513 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_514 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_515 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_516 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_517 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_518 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_519 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_520 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_521 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_522 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_523 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_524 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_525 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_526 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_527 (.DIODE(_06120_));
 sky130_fd_sc_hd__diode_2 ANTENNA_528 (.DIODE(_06704_));
 sky130_fd_sc_hd__diode_2 ANTENNA_529 (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_04730_));
 sky130_fd_sc_hd__diode_2 ANTENNA_530 (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA_531 (.DIODE(\core.fetchProgramCounter[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_532 (.DIODE(\coreWBInterface.readDataBuffered[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_533 (.DIODE(\coreWBInterface.readDataBuffered[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_534 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_535 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_536 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_537 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_538 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_539 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_04730_));
 sky130_fd_sc_hd__diode_2 ANTENNA_540 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_541 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_542 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_543 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_544 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_545 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_546 (.DIODE(net1669));
 sky130_fd_sc_hd__diode_2 ANTENNA_547 (.DIODE(net1762));
 sky130_fd_sc_hd__diode_2 ANTENNA_548 (.DIODE(net1764));
 sky130_fd_sc_hd__diode_2 ANTENNA_549 (.DIODE(net1764));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_04730_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_04852_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_05108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_05108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_05217_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_05447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_05447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_05748_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_05901_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_06012_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_06043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_06043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_06055_));
 sky130_fd_sc_hd__conb_1 ExperiarCore_1911 (.LO(net1911));
 sky130_fd_sc_hd__decap_6 FILLER_0_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_954 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_6 _08815_ (.A(\core.pipe2_stall ),
    .Y(_03807_));
 sky130_fd_sc_hd__inv_6 _08816_ (.A(net1798),
    .Y(_03808_));
 sky130_fd_sc_hd__inv_2 _08817_ (.A(\core.csr.traps.mtval.csrReadData[0] ),
    .Y(_03809_));
 sky130_fd_sc_hd__inv_2 _08818_ (.A(\core.csr.traps.mtvec.csrReadData[6] ),
    .Y(_03810_));
 sky130_fd_sc_hd__inv_2 _08819_ (.A(\core.csr.trapReturnVector[24] ),
    .Y(_03811_));
 sky130_fd_sc_hd__inv_2 _08820_ (.A(\core.csr.trapReturnVector[3] ),
    .Y(_03812_));
 sky130_fd_sc_hd__inv_2 _08821_ (.A(\core.csr.instretTimer.currentValue[63] ),
    .Y(_03813_));
 sky130_fd_sc_hd__inv_2 _08822_ (.A(\core.fetchProgramCounter[1] ),
    .Y(_03814_));
 sky130_fd_sc_hd__inv_2 _08823_ (.A(\core.fetchProgramCounter[0] ),
    .Y(_03815_));
 sky130_fd_sc_hd__inv_2 _08824_ (.A(\jtag.managementState[0] ),
    .Y(_03816_));
 sky130_fd_sc_hd__inv_4 _08825_ (.A(net1723),
    .Y(_03817_));
 sky130_fd_sc_hd__inv_2 _08826_ (.A(\jtag.state[2] ),
    .Y(_03818_));
 sky130_fd_sc_hd__inv_2 _08827_ (.A(net1721),
    .Y(_03819_));
 sky130_fd_sc_hd__inv_2 _08828_ (.A(net1730),
    .Y(_03820_));
 sky130_fd_sc_hd__inv_2 _08829_ (.A(\core.fetchProgramCounter[28] ),
    .Y(_03821_));
 sky130_fd_sc_hd__inv_2 _08830_ (.A(net409),
    .Y(_03822_));
 sky130_fd_sc_hd__clkinv_4 _08831_ (.A(net474),
    .Y(_03823_));
 sky130_fd_sc_hd__inv_2 _08832_ (.A(net465),
    .Y(_03824_));
 sky130_fd_sc_hd__inv_2 _08833_ (.A(net481),
    .Y(_03825_));
 sky130_fd_sc_hd__clkinv_4 _08834_ (.A(net479),
    .Y(_03826_));
 sky130_fd_sc_hd__inv_6 _08835_ (.A(net472),
    .Y(_03827_));
 sky130_fd_sc_hd__inv_6 _08836_ (.A(net1719),
    .Y(_03828_));
 sky130_fd_sc_hd__clkinv_2 _08837_ (.A(net1749),
    .Y(_03829_));
 sky130_fd_sc_hd__clkinv_4 _08838_ (.A(net1750),
    .Y(_03830_));
 sky130_fd_sc_hd__inv_2 _08839_ (.A(net1752),
    .Y(_03831_));
 sky130_fd_sc_hd__inv_2 _08840_ (.A(\core.pipe0_currentInstruction[27] ),
    .Y(_03832_));
 sky130_fd_sc_hd__inv_2 _08841_ (.A(\core.pipe0_currentInstruction[26] ),
    .Y(_03833_));
 sky130_fd_sc_hd__clkinv_2 _08842_ (.A(net1756),
    .Y(_03834_));
 sky130_fd_sc_hd__inv_8 _08843_ (.A(net1765),
    .Y(_03835_));
 sky130_fd_sc_hd__inv_2 _08844_ (.A(net1773),
    .Y(_03836_));
 sky130_fd_sc_hd__inv_6 _08845_ (.A(net1776),
    .Y(_03837_));
 sky130_fd_sc_hd__inv_2 _08846_ (.A(net1781),
    .Y(_03838_));
 sky130_fd_sc_hd__inv_2 _08847_ (.A(\core.pipe0_currentInstruction[18] ),
    .Y(_03839_));
 sky130_fd_sc_hd__clkinv_2 _08848_ (.A(net1786),
    .Y(_03840_));
 sky130_fd_sc_hd__inv_2 _08849_ (.A(net1788),
    .Y(_03841_));
 sky130_fd_sc_hd__inv_2 _08850_ (.A(net1793),
    .Y(_03842_));
 sky130_fd_sc_hd__clkinv_2 _08851_ (.A(\core.pipe0_currentInstruction[12] ),
    .Y(_03843_));
 sky130_fd_sc_hd__clkinv_2 _08852_ (.A(\core.pipe0_currentInstruction[10] ),
    .Y(_03844_));
 sky130_fd_sc_hd__inv_2 _08853_ (.A(\core.pipe0_currentInstruction[8] ),
    .Y(_03845_));
 sky130_fd_sc_hd__inv_2 _08854_ (.A(\core.pipe0_currentInstruction[6] ),
    .Y(_03846_));
 sky130_fd_sc_hd__inv_2 _08855_ (.A(\core.csr.currentInstruction[5] ),
    .Y(_03847_));
 sky130_fd_sc_hd__inv_2 _08856_ (.A(\core.csr.currentInstruction[2] ),
    .Y(_03848_));
 sky130_fd_sc_hd__inv_2 _08857_ (.A(net1745),
    .Y(_03849_));
 sky130_fd_sc_hd__inv_2 _08858_ (.A(net1746),
    .Y(_03850_));
 sky130_fd_sc_hd__inv_2 _08859_ (.A(net1902),
    .Y(_03851_));
 sky130_fd_sc_hd__inv_2 _08860_ (.A(net9),
    .Y(_03852_));
 sky130_fd_sc_hd__inv_2 _08861_ (.A(net189),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2b_4 _08862_ (.A_N(\coreWBInterface.state[1] ),
    .B(\coreWBInterface.state[0] ),
    .Y(_03854_));
 sky130_fd_sc_hd__inv_2 _08863_ (.A(_03854_),
    .Y(net371));
 sky130_fd_sc_hd__and2b_1 _08864_ (.A_N(\core.cancelStall ),
    .B(\core.pipe0_fetch.currentPipeStall ),
    .X(_03855_));
 sky130_fd_sc_hd__nand2b_1 _08865_ (.A_N(\core.cancelStall ),
    .B(\core.pipe0_fetch.currentPipeStall ),
    .Y(_03856_));
 sky130_fd_sc_hd__nand3_2 _08866_ (.A(\core.pipe0_currentInstruction[1] ),
    .B(\core.pipe0_currentInstruction[0] ),
    .C(net1630),
    .Y(_03857_));
 sky130_fd_sc_hd__or3_4 _08867_ (.A(\core.pipe0_currentInstruction[3] ),
    .B(\core.pipe0_currentInstruction[2] ),
    .C(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__nand2_2 _08868_ (.A(\core.pipe0_currentInstruction[4] ),
    .B(net1630),
    .Y(_03859_));
 sky130_fd_sc_hd__nand3_2 _08869_ (.A(\core.pipe0_currentInstruction[5] ),
    .B(\core.pipe0_currentInstruction[4] ),
    .C(net1630),
    .Y(_03860_));
 sky130_fd_sc_hd__or3_4 _08870_ (.A(_03846_),
    .B(_03858_),
    .C(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__or4_1 _08871_ (.A(\core.pipe0_currentInstruction[10] ),
    .B(\core.pipe0_currentInstruction[9] ),
    .C(\core.pipe0_currentInstruction[8] ),
    .D(\core.pipe0_currentInstruction[7] ),
    .X(_03862_));
 sky130_fd_sc_hd__or3_2 _08872_ (.A(\core.pipe0_currentInstruction[13] ),
    .B(\core.pipe0_currentInstruction[11] ),
    .C(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__or4_1 _08873_ (.A(net1789),
    .B(net1793),
    .C(net1795),
    .D(\core.pipe0_currentInstruction[12] ),
    .X(_03864_));
 sky130_fd_sc_hd__or4_1 _08874_ (.A(net1755),
    .B(net1762),
    .C(\core.pipe0_currentInstruction[18] ),
    .D(net1784),
    .X(_03865_));
 sky130_fd_sc_hd__or4_1 _08875_ (.A(\core.pipe0_currentInstruction[26] ),
    .B(\core.pipe0_currentInstruction[25] ),
    .C(_03864_),
    .D(_03865_),
    .X(_03866_));
 sky130_fd_sc_hd__or3_4 _08876_ (.A(_03861_),
    .B(_03863_),
    .C(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__or3_4 _08877_ (.A(\core.pipe0_currentInstruction[29] ),
    .B(\core.pipe0_currentInstruction[28] ),
    .C(\core.pipe0_currentInstruction[27] ),
    .X(_03868_));
 sky130_fd_sc_hd__or2_2 _08878_ (.A(net1751),
    .B(net1752),
    .X(_03869_));
 sky130_fd_sc_hd__or4_2 _08879_ (.A(_03828_),
    .B(net1764),
    .C(net1771),
    .D(net1780),
    .X(_03870_));
 sky130_fd_sc_hd__nor4_4 _08880_ (.A(_03867_),
    .B(_03868_),
    .C(_03869_),
    .D(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__and2_4 _08881_ (.A(net1684),
    .B(_03871_),
    .X(net444));
 sky130_fd_sc_hd__nand2_2 _08882_ (.A(net1776),
    .B(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__inv_6 _08883_ (.A(net1098),
    .Y(net443));
 sky130_fd_sc_hd__or2_4 _08884_ (.A(\coreWBInterface.state[1] ),
    .B(\coreWBInterface.state[0] ),
    .X(net333));
 sky130_fd_sc_hd__or3_4 _08885_ (.A(\core.fetchProgramCounter[31] ),
    .B(\core.fetchProgramCounter[30] ),
    .C(\core.fetchProgramCounter[29] ),
    .X(_03873_));
 sky130_fd_sc_hd__or4_4 _08886_ (.A(\core.fetchProgramCounter[27] ),
    .B(\core.fetchProgramCounter[26] ),
    .C(\core.fetchProgramCounter[25] ),
    .D(\core.fetchProgramCounter[24] ),
    .X(_03874_));
 sky130_fd_sc_hd__nor3_4 _08887_ (.A(\core.fetchProgramCounter[28] ),
    .B(_03873_),
    .C(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__clkinv_4 _08888_ (.A(net1601),
    .Y(_03876_));
 sky130_fd_sc_hd__or3b_4 _08889_ (.A(_03857_),
    .B(\core.pipe0_currentInstruction[3] ),
    .C_N(\core.pipe0_currentInstruction[2] ),
    .X(_03877_));
 sky130_fd_sc_hd__nor4_4 _08890_ (.A(\core.pipe0_currentInstruction[6] ),
    .B(\core.pipe0_currentInstruction[5] ),
    .C(_03859_),
    .D(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__or4_4 _08891_ (.A(\core.pipe0_currentInstruction[6] ),
    .B(\core.pipe0_currentInstruction[5] ),
    .C(_03859_),
    .D(_03877_),
    .X(_03879_));
 sky130_fd_sc_hd__or2_2 _08892_ (.A(net452),
    .B(net1258),
    .X(_03880_));
 sky130_fd_sc_hd__nor2_8 _08893_ (.A(net1674),
    .B(net1633),
    .Y(_03881_));
 sky130_fd_sc_hd__nand2_8 _08894_ (.A(net1782),
    .B(net1631),
    .Y(_03882_));
 sky130_fd_sc_hd__nor2_2 _08895_ (.A(net1670),
    .B(net1633),
    .Y(_03883_));
 sky130_fd_sc_hd__nand2_2 _08896_ (.A(net1786),
    .B(net1631),
    .Y(_03884_));
 sky130_fd_sc_hd__nor2_2 _08897_ (.A(_03839_),
    .B(net1634),
    .Y(_03885_));
 sky130_fd_sc_hd__nand2_8 _08898_ (.A(\core.pipe0_currentInstruction[18] ),
    .B(net1630),
    .Y(_03886_));
 sky130_fd_sc_hd__nor2_8 _08899_ (.A(net1663),
    .B(net1633),
    .Y(_03887_));
 sky130_fd_sc_hd__nand2_2 _08900_ (.A(net1787),
    .B(net1629),
    .Y(_03888_));
 sky130_fd_sc_hd__nor2_2 _08901_ (.A(net1650),
    .B(net1633),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2_2 _08902_ (.A(net1793),
    .B(net1632),
    .Y(_03890_));
 sky130_fd_sc_hd__and3_1 _08903_ (.A(net1563),
    .B(net1534),
    .C(net1460),
    .X(_03891_));
 sky130_fd_sc_hd__and3_2 _08904_ (.A(net1596),
    .B(net1576),
    .C(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__or3b_1 _08905_ (.A(net1796),
    .B(net1799),
    .C_N(net1800),
    .X(_03893_));
 sky130_fd_sc_hd__or4b_4 _08906_ (.A(net1796),
    .B(net1799),
    .C(\core.csr.currentInstruction[12] ),
    .D_N(net1800),
    .X(_03894_));
 sky130_fd_sc_hd__o31ai_2 _08907_ (.A1(net1796),
    .A2(net1799),
    .A3(\core.csr.currentInstruction[12] ),
    .B1(net1800),
    .Y(_03895_));
 sky130_fd_sc_hd__nand3b_4 _08908_ (.A_N(net1798),
    .B(\core.csr.currentInstruction[1] ),
    .C(\core.csr.currentInstruction[0] ),
    .Y(_03896_));
 sky130_fd_sc_hd__or2_4 _08909_ (.A(\core.csr.currentInstruction[3] ),
    .B(\core.csr.currentInstruction[2] ),
    .X(_03897_));
 sky130_fd_sc_hd__nor2_8 _08910_ (.A(_03896_),
    .B(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__nand2b_2 _08911_ (.A_N(net1796),
    .B(\core.csr.currentInstruction[5] ),
    .Y(_03899_));
 sky130_fd_sc_hd__nor2_1 _08912_ (.A(\core.csr.currentInstruction[6] ),
    .B(\core.csr.currentInstruction[4] ),
    .Y(_03900_));
 sky130_fd_sc_hd__a31o_4 _08913_ (.A1(_03847_),
    .A2(_03895_),
    .A3(_03900_),
    .B1(net1797),
    .X(_03901_));
 sky130_fd_sc_hd__or3b_4 _08914_ (.A(net1796),
    .B(net1800),
    .C_N(\core.csr.currentInstruction[12] ),
    .X(_03902_));
 sky130_fd_sc_hd__nand2b_4 _08915_ (.A_N(net1798),
    .B(net1801),
    .Y(_03903_));
 sky130_fd_sc_hd__and2_4 _08916_ (.A(_03808_),
    .B(\core.csr.currentInstruction[11] ),
    .X(_03904_));
 sky130_fd_sc_hd__nand2b_1 _08917_ (.A_N(net1798),
    .B(\core.csr.currentInstruction[11] ),
    .Y(_03905_));
 sky130_fd_sc_hd__and2_2 _08918_ (.A(_03808_),
    .B(\core.csr.currentInstruction[10] ),
    .X(_03906_));
 sky130_fd_sc_hd__nand2b_2 _08919_ (.A_N(net1798),
    .B(\core.csr.currentInstruction[10] ),
    .Y(_03907_));
 sky130_fd_sc_hd__and3_4 _08920_ (.A(_03903_),
    .B(_03905_),
    .C(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__and2_4 _08921_ (.A(_03808_),
    .B(\core.csr.currentInstruction[7] ),
    .X(_03909_));
 sky130_fd_sc_hd__nand2_8 _08922_ (.A(_03808_),
    .B(\core.csr.currentInstruction[7] ),
    .Y(_03910_));
 sky130_fd_sc_hd__nand2_4 _08923_ (.A(_03808_),
    .B(\core.csr.currentInstruction[8] ),
    .Y(_03911_));
 sky130_fd_sc_hd__and3_2 _08924_ (.A(_03908_),
    .B(_03910_),
    .C(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__o21ba_4 _08925_ (.A1(net1800),
    .A2(\core.csr.currentInstruction[12] ),
    .B1_N(net1796),
    .X(_03913_));
 sky130_fd_sc_hd__o21bai_2 _08926_ (.A1(net1800),
    .A2(\core.csr.currentInstruction[12] ),
    .B1_N(net1796),
    .Y(_03914_));
 sky130_fd_sc_hd__a21oi_4 _08927_ (.A1(_03808_),
    .A2(net1799),
    .B1(_03913_),
    .Y(_03915_));
 sky130_fd_sc_hd__nand2_1 _08928_ (.A(\core.csr.currentInstruction[6] ),
    .B(\core.csr.currentInstruction[4] ),
    .Y(_03916_));
 sky130_fd_sc_hd__or4_4 _08929_ (.A(_03896_),
    .B(_03897_),
    .C(_03899_),
    .D(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__a211oi_4 _08930_ (.A1(_03902_),
    .A2(_03912_),
    .B1(_03915_),
    .C1(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__a21oi_4 _08931_ (.A1(_03898_),
    .A2(_03901_),
    .B1(net1247),
    .Y(_03919_));
 sky130_fd_sc_hd__or4bb_1 _08932_ (.A(net1796),
    .B(net1800),
    .C_N(\core.csr.currentInstruction[12] ),
    .D_N(net1799),
    .X(_03920_));
 sky130_fd_sc_hd__o211a_1 _08933_ (.A1(net1799),
    .A2(_03913_),
    .B1(_03920_),
    .C1(\core.csr.currentInstruction[30] ),
    .X(_03921_));
 sky130_fd_sc_hd__or4_1 _08934_ (.A(\core.csr.currentInstruction[29] ),
    .B(\core.csr.currentInstruction[28] ),
    .C(\core.csr.currentInstruction[27] ),
    .D(\core.csr.currentInstruction[26] ),
    .X(_03922_));
 sky130_fd_sc_hd__or3_1 _08935_ (.A(\core.csr.currentInstruction[31] ),
    .B(\core.csr.currentInstruction[25] ),
    .C(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__a2bb2o_2 _08936_ (.A1_N(_03921_),
    .A2_N(_03923_),
    .B1(_03899_),
    .B2(_03902_),
    .X(_03924_));
 sky130_fd_sc_hd__or3b_2 _08937_ (.A(net1797),
    .B(\core.csr.currentInstruction[6] ),
    .C_N(\core.csr.currentInstruction[4] ),
    .X(_03925_));
 sky130_fd_sc_hd__inv_2 _08938_ (.A(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__and3_4 _08939_ (.A(_03898_),
    .B(_03924_),
    .C(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__or2_4 _08940_ (.A(_03848_),
    .B(_03896_),
    .X(_03928_));
 sky130_fd_sc_hd__or2_2 _08941_ (.A(\core.csr.currentInstruction[3] ),
    .B(_03925_),
    .X(_03929_));
 sky130_fd_sc_hd__nor2_2 _08942_ (.A(\core.csr.currentInstruction[4] ),
    .B(_03899_),
    .Y(_03930_));
 sky130_fd_sc_hd__o211ai_4 _08943_ (.A1(\core.csr.currentInstruction[3] ),
    .A2(_03915_),
    .B1(_03930_),
    .C1(\core.csr.currentInstruction[6] ),
    .Y(_03931_));
 sky130_fd_sc_hd__a21oi_4 _08944_ (.A1(_03929_),
    .A2(_03931_),
    .B1(_03928_),
    .Y(_03932_));
 sky130_fd_sc_hd__a21o_4 _08945_ (.A1(_03929_),
    .A2(_03931_),
    .B1(_03928_),
    .X(_03933_));
 sky130_fd_sc_hd__nor2_8 _08946_ (.A(_03927_),
    .B(net1244),
    .Y(_03934_));
 sky130_fd_sc_hd__or2_4 _08947_ (.A(_03927_),
    .B(net1246),
    .X(_03935_));
 sky130_fd_sc_hd__nand2_1 _08948_ (.A(_03919_),
    .B(net1189),
    .Y(_03936_));
 sky130_fd_sc_hd__xnor2_1 _08949_ (.A(net1534),
    .B(_03911_),
    .Y(_03937_));
 sky130_fd_sc_hd__xnor2_1 _08950_ (.A(net1598),
    .B(_03904_),
    .Y(_03938_));
 sky130_fd_sc_hd__xnor2_1 _08951_ (.A(net1575),
    .B(_03903_),
    .Y(_03939_));
 sky130_fd_sc_hd__o221a_1 _08952_ (.A1(net1570),
    .A2(_03907_),
    .B1(_03909_),
    .B2(net1461),
    .C1(_03938_),
    .X(_03940_));
 sky130_fd_sc_hd__o221a_1 _08953_ (.A1(net1563),
    .A2(_03906_),
    .B1(_03910_),
    .B2(net1502),
    .C1(_03937_),
    .X(_03941_));
 sky130_fd_sc_hd__and3_1 _08954_ (.A(_03939_),
    .B(_03940_),
    .C(_03941_),
    .X(_03942_));
 sky130_fd_sc_hd__o221a_1 _08955_ (.A1(net1563),
    .A2(_03906_),
    .B1(_03910_),
    .B2(net1502),
    .C1(_03939_),
    .X(_03943_));
 sky130_fd_sc_hd__and4_2 _08956_ (.A(_03936_),
    .B(_03937_),
    .C(_03940_),
    .D(_03943_),
    .X(_03944_));
 sky130_fd_sc_hd__nor2_4 _08957_ (.A(_03892_),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__or2_4 _08958_ (.A(_03892_),
    .B(_03944_),
    .X(_03946_));
 sky130_fd_sc_hd__mux4_1 _08959_ (.A0(\core.registers[16][11] ),
    .A1(\core.registers[17][11] ),
    .A2(\core.registers[20][11] ),
    .A3(\core.registers[21][11] ),
    .S0(net1522),
    .S1(net1590),
    .X(_03947_));
 sky130_fd_sc_hd__a22o_1 _08960_ (.A1(net1659),
    .A2(\core.registers[22][11] ),
    .B1(\core.registers[23][11] ),
    .B2(net1522),
    .X(_03948_));
 sky130_fd_sc_hd__a22o_1 _08961_ (.A1(net1659),
    .A2(\core.registers[18][11] ),
    .B1(\core.registers[19][11] ),
    .B2(net1522),
    .X(_03949_));
 sky130_fd_sc_hd__mux2_1 _08962_ (.A0(_03948_),
    .A1(_03949_),
    .S(net1578),
    .X(_03950_));
 sky130_fd_sc_hd__a21o_1 _08963_ (.A1(net1558),
    .A2(_03950_),
    .B1(net1568),
    .X(_03951_));
 sky130_fd_sc_hd__a21oi_1 _08964_ (.A1(net1538),
    .A2(_03947_),
    .B1(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__a22o_1 _08965_ (.A1(net1654),
    .A2(\core.registers[30][11] ),
    .B1(\core.registers[31][11] ),
    .B2(net1503),
    .X(_03953_));
 sky130_fd_sc_hd__a22o_1 _08966_ (.A1(net1654),
    .A2(\core.registers[26][11] ),
    .B1(\core.registers[27][11] ),
    .B2(net1505),
    .X(_03954_));
 sky130_fd_sc_hd__mux2_2 _08967_ (.A0(_03953_),
    .A1(_03954_),
    .S(net1577),
    .X(_03955_));
 sky130_fd_sc_hd__mux4_1 _08968_ (.A0(\core.registers[24][11] ),
    .A1(\core.registers[25][11] ),
    .A2(\core.registers[28][11] ),
    .A3(\core.registers[29][11] ),
    .S0(net1505),
    .S1(net1588),
    .X(_03956_));
 sky130_fd_sc_hd__a21o_1 _08969_ (.A1(net1535),
    .A2(_03956_),
    .B1(net1565),
    .X(_03957_));
 sky130_fd_sc_hd__a21oi_4 _08970_ (.A1(net1552),
    .A2(_03955_),
    .B1(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__mux4_1 _08971_ (.A0(\core.registers[0][11] ),
    .A1(\core.registers[1][11] ),
    .A2(\core.registers[4][11] ),
    .A3(\core.registers[5][11] ),
    .S0(net1517),
    .S1(net1590),
    .X(_03959_));
 sky130_fd_sc_hd__and2_1 _08972_ (.A(net1539),
    .B(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__a22o_1 _08973_ (.A1(net1659),
    .A2(\core.registers[6][11] ),
    .B1(\core.registers[7][11] ),
    .B2(net1522),
    .X(_03961_));
 sky130_fd_sc_hd__a22o_1 _08974_ (.A1(net1659),
    .A2(\core.registers[2][11] ),
    .B1(\core.registers[3][11] ),
    .B2(net1522),
    .X(_03962_));
 sky130_fd_sc_hd__mux2_1 _08975_ (.A0(_03961_),
    .A1(_03962_),
    .S(net1579),
    .X(_03963_));
 sky130_fd_sc_hd__a21o_1 _08976_ (.A1(net1558),
    .A2(_03963_),
    .B1(net1568),
    .X(_03964_));
 sky130_fd_sc_hd__nor2_1 _08977_ (.A(_03960_),
    .B(_03964_),
    .Y(_03965_));
 sky130_fd_sc_hd__mux4_1 _08978_ (.A0(\core.registers[8][11] ),
    .A1(\core.registers[9][11] ),
    .A2(\core.registers[12][11] ),
    .A3(\core.registers[13][11] ),
    .S0(net1517),
    .S1(net1590),
    .X(_03966_));
 sky130_fd_sc_hd__nand2_1 _08979_ (.A(net1539),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__a22o_1 _08980_ (.A1(net1659),
    .A2(\core.registers[14][11] ),
    .B1(\core.registers[15][11] ),
    .B2(net1522),
    .X(_03968_));
 sky130_fd_sc_hd__a22o_1 _08981_ (.A1(net1659),
    .A2(\core.registers[10][11] ),
    .B1(\core.registers[11][11] ),
    .B2(net1522),
    .X(_03969_));
 sky130_fd_sc_hd__mux2_1 _08982_ (.A0(_03968_),
    .A1(_03969_),
    .S(net1578),
    .X(_03970_));
 sky130_fd_sc_hd__a21oi_1 _08983_ (.A1(net1557),
    .A2(_03970_),
    .B1(net1564),
    .Y(_03971_));
 sky130_fd_sc_hd__a21o_1 _08984_ (.A1(_03967_),
    .A2(_03971_),
    .B1(net1599),
    .X(_03972_));
 sky130_fd_sc_hd__o32a_4 _08985_ (.A1(net1595),
    .A2(_03952_),
    .A3(_03958_),
    .B1(_03965_),
    .B2(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__nand2b_1 _08986_ (.A_N(net1745),
    .B(\memoryController.last_data_enableWB ),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _08987_ (.A(\localMemoryInterface.coreReadReady ),
    .B(\localMemoryInterface.lastCoreByteSelect[3] ),
    .Y(_03975_));
 sky130_fd_sc_hd__mux2_8 _08988_ (.A0(net126),
    .A1(net161),
    .S(net1736),
    .X(_03976_));
 sky130_fd_sc_hd__o32a_1 _08989_ (.A1(net1638),
    .A2(net1624),
    .A3(_03976_),
    .B1(net1625),
    .B2(\coreWBInterface.readDataBuffered[27] ),
    .X(_03977_));
 sky130_fd_sc_hd__o21ba_2 _08990_ (.A1(net1799),
    .A2(net1800),
    .B1_N(net1796),
    .X(_03978_));
 sky130_fd_sc_hd__or4b_2 _08991_ (.A(net1797),
    .B(\core.csr.currentInstruction[6] ),
    .C(\core.csr.currentInstruction[4] ),
    .D_N(\core.csr.currentInstruction[5] ),
    .X(_03979_));
 sky130_fd_sc_hd__a2111oi_4 _08992_ (.A1(_03894_),
    .A2(_03978_),
    .B1(_03979_),
    .C1(_03896_),
    .D1(_03897_),
    .Y(_03980_));
 sky130_fd_sc_hd__a21oi_4 _08993_ (.A1(_03898_),
    .A2(_03901_),
    .B1(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__a21o_4 _08994_ (.A1(_03898_),
    .A2(_03901_),
    .B1(_03980_),
    .X(_03982_));
 sky130_fd_sc_hd__nor2_2 _08995_ (.A(\core.pipe1_resultRegister[0] ),
    .B(_03913_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _08996_ (.A(_03830_),
    .B(_03914_),
    .Y(_03984_));
 sky130_fd_sc_hd__or3_1 _08997_ (.A(net1712),
    .B(_03981_),
    .C(_03983_),
    .X(_03985_));
 sky130_fd_sc_hd__o31a_4 _08998_ (.A1(net1749),
    .A2(_03894_),
    .A3(_03981_),
    .B1(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__nor2_1 _08999_ (.A(_03977_),
    .B(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__nor2_2 _09000_ (.A(net1712),
    .B(net1750),
    .Y(_03988_));
 sky130_fd_sc_hd__nand2_8 _09001_ (.A(\localMemoryInterface.coreReadReady ),
    .B(\localMemoryInterface.lastCoreByteSelect[1] ),
    .Y(_03989_));
 sky130_fd_sc_hd__mux2_8 _09002_ (.A0(net113),
    .A1(net148),
    .S(net1735),
    .X(_03990_));
 sky130_fd_sc_hd__o32a_1 _09003_ (.A1(net1638),
    .A2(_03989_),
    .A3(_03990_),
    .B1(net1625),
    .B2(\coreWBInterface.readDataBuffered[15] ),
    .X(_03991_));
 sky130_fd_sc_hd__mux2_8 _09004_ (.A0(net131),
    .A1(net166),
    .S(net1736),
    .X(_03992_));
 sky130_fd_sc_hd__o32a_2 _09005_ (.A1(net1638),
    .A2(net1624),
    .A3(_03992_),
    .B1(net1628),
    .B2(\coreWBInterface.readDataBuffered[31] ),
    .X(_03993_));
 sky130_fd_sc_hd__mux2_1 _09006_ (.A0(_03991_),
    .A1(_03993_),
    .S(net1749),
    .X(_03994_));
 sky130_fd_sc_hd__nand2_1 _09007_ (.A(\localMemoryInterface.coreReadReady ),
    .B(\localMemoryInterface.lastCoreByteSelect[2] ),
    .Y(_03995_));
 sky130_fd_sc_hd__mux2_8 _09008_ (.A0(net122),
    .A1(net157),
    .S(net1737),
    .X(_03996_));
 sky130_fd_sc_hd__o32a_2 _09009_ (.A1(net1638),
    .A2(net1622),
    .A3(_03996_),
    .B1(net1628),
    .B2(\coreWBInterface.readDataBuffered[23] ),
    .X(_03997_));
 sky130_fd_sc_hd__nand2_2 _09010_ (.A(\localMemoryInterface.lastCoreByteSelect[0] ),
    .B(\localMemoryInterface.coreReadReady ),
    .Y(_03998_));
 sky130_fd_sc_hd__mux2_8 _09011_ (.A0(net168),
    .A1(net139),
    .S(net1734),
    .X(_03999_));
 sky130_fd_sc_hd__or3_1 _09012_ (.A(net1640),
    .B(net1619),
    .C(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__nor2_2 _09013_ (.A(net1749),
    .B(net1750),
    .Y(_04001_));
 sky130_fd_sc_hd__or2_4 _09014_ (.A(net1749),
    .B(net1750),
    .X(_04002_));
 sky130_fd_sc_hd__o21a_1 _09015_ (.A1(\coreWBInterface.readDataBuffered[7] ),
    .A2(net1628),
    .B1(net1617),
    .X(_04003_));
 sky130_fd_sc_hd__a22o_1 _09016_ (.A1(net1458),
    .A2(_03997_),
    .B1(_04000_),
    .B2(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__a21o_1 _09017_ (.A1(net1750),
    .A2(_03994_),
    .B1(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__a211o_4 _09018_ (.A1(net1750),
    .A2(_03994_),
    .B1(_04004_),
    .C1(_03913_),
    .X(_04006_));
 sky130_fd_sc_hd__nor2_2 _09019_ (.A(net1749),
    .B(_03830_),
    .Y(_04007_));
 sky130_fd_sc_hd__nand2_4 _09020_ (.A(net1712),
    .B(net1750),
    .Y(_04008_));
 sky130_fd_sc_hd__or2_1 _09021_ (.A(_03991_),
    .B(net1616),
    .X(_04009_));
 sky130_fd_sc_hd__a21o_1 _09022_ (.A1(net1712),
    .A2(_03997_),
    .B1(_03830_),
    .X(_04010_));
 sky130_fd_sc_hd__o21ba_1 _09023_ (.A1(net1712),
    .A2(_03993_),
    .B1_N(_03978_),
    .X(_04011_));
 sky130_fd_sc_hd__a31o_2 _09024_ (.A1(_04009_),
    .A2(_04010_),
    .A3(_04011_),
    .B1(_03915_),
    .X(_04012_));
 sky130_fd_sc_hd__nand2_4 _09025_ (.A(_04006_),
    .B(_04012_),
    .Y(_04013_));
 sky130_fd_sc_hd__nand2_4 _09026_ (.A(_03986_),
    .B(_04013_),
    .Y(_04014_));
 sky130_fd_sc_hd__nand2_2 _09027_ (.A(net1458),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__nor2_2 _09028_ (.A(net1712),
    .B(_03830_),
    .Y(_04016_));
 sky130_fd_sc_hd__nand2_2 _09029_ (.A(\core.pipe1_resultRegister[1] ),
    .B(net1750),
    .Y(_04017_));
 sky130_fd_sc_hd__a31o_4 _09030_ (.A1(_04006_),
    .A2(_04012_),
    .A3(_04016_),
    .B1(net1617),
    .X(_04018_));
 sky130_fd_sc_hd__mux2_1 _09031_ (.A0(_03894_),
    .A1(_03914_),
    .S(net1750),
    .X(_04019_));
 sky130_fd_sc_hd__nand2_1 _09032_ (.A(net1712),
    .B(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__and3_1 _09033_ (.A(_03982_),
    .B(_04017_),
    .C(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__nor2_4 _09034_ (.A(_04013_),
    .B(net1243),
    .Y(_04022_));
 sky130_fd_sc_hd__mux2_8 _09035_ (.A0(net117),
    .A1(net153),
    .S(net1736),
    .X(_04023_));
 sky130_fd_sc_hd__o32a_1 _09036_ (.A1(net1638),
    .A2(net1622),
    .A3(_04023_),
    .B1(net1625),
    .B2(\coreWBInterface.readDataBuffered[19] ),
    .X(_04024_));
 sky130_fd_sc_hd__a21o_1 _09037_ (.A1(net1243),
    .A2(_04024_),
    .B1(_04022_),
    .X(_04025_));
 sky130_fd_sc_hd__a2bb2o_1 _09038_ (.A1_N(_03987_),
    .A2_N(_04015_),
    .B1(_04025_),
    .B2(_04007_),
    .X(_04026_));
 sky130_fd_sc_hd__or2_2 _09039_ (.A(_03894_),
    .B(_04008_),
    .X(_04027_));
 sky130_fd_sc_hd__o211a_2 _09040_ (.A1(net1712),
    .A2(_04019_),
    .B1(_03901_),
    .C1(_03898_),
    .X(_04028_));
 sky130_fd_sc_hd__and2_4 _09041_ (.A(_04027_),
    .B(_04028_),
    .X(_04029_));
 sky130_fd_sc_hd__nand2_2 _09042_ (.A(_04027_),
    .B(_04028_),
    .Y(_04030_));
 sky130_fd_sc_hd__and3_4 _09043_ (.A(net1712),
    .B(_03982_),
    .C(_03984_),
    .X(_04031_));
 sky130_fd_sc_hd__mux2_4 _09044_ (.A0(net109),
    .A1(net144),
    .S(net1735),
    .X(_04032_));
 sky130_fd_sc_hd__nor2_1 _09045_ (.A(_03989_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__nand2_1 _09046_ (.A(\memoryController.last_data_enableLocalMemory ),
    .B(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__o211a_1 _09047_ (.A1(\coreWBInterface.readDataBuffered[11] ),
    .A2(net1625),
    .B1(_04031_),
    .C1(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__nor2_1 _09048_ (.A(_04013_),
    .B(_04031_),
    .Y(_04036_));
 sky130_fd_sc_hd__nor2_1 _09049_ (.A(_04002_),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__or2_4 _09050_ (.A(_04002_),
    .B(_04036_),
    .X(_04038_));
 sky130_fd_sc_hd__o22a_1 _09051_ (.A1(_04018_),
    .A2(_04026_),
    .B1(_04035_),
    .B2(_04038_),
    .X(_04039_));
 sky130_fd_sc_hd__nand2_1 _09052_ (.A(_04029_),
    .B(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__a221oi_1 _09053_ (.A1(\core.pipe1_csrData[11] ),
    .A2(net1249),
    .B1(_03927_),
    .B2(\core.pipe1_resultRegister[11] ),
    .C1(net1244),
    .Y(_04041_));
 sky130_fd_sc_hd__o2bb2a_2 _09054_ (.A1_N(_04041_),
    .A2_N(_04040_),
    .B1(_03933_),
    .B2(\core.pipe1_resultRegister[11] ),
    .X(_04042_));
 sky130_fd_sc_hd__and3b_1 _09055_ (.A_N(_03892_),
    .B(_03936_),
    .C(_03942_),
    .X(_04043_));
 sky130_fd_sc_hd__a2bb2o_4 _09056_ (.A1_N(net1044),
    .A2_N(_03973_),
    .B1(net764),
    .B2(net1095),
    .X(_04044_));
 sky130_fd_sc_hd__o21ai_4 _09057_ (.A1(net1263),
    .A2(_04044_),
    .B1(_03880_),
    .Y(_04045_));
 sky130_fd_sc_hd__clkinv_2 _09058_ (.A(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2_8 _09059_ (.A(\core.pipe0_currentInstruction[13] ),
    .B(net1629),
    .Y(_04047_));
 sky130_fd_sc_hd__nand2_8 _09060_ (.A(\core.pipe0_currentInstruction[12] ),
    .B(net1629),
    .Y(_04048_));
 sky130_fd_sc_hd__nor2_4 _09061_ (.A(_03843_),
    .B(_04047_),
    .Y(_04049_));
 sky130_fd_sc_hd__and3b_1 _09062_ (.A_N(\core.pipe0_currentInstruction[4] ),
    .B(net1630),
    .C(\core.pipe0_currentInstruction[5] ),
    .X(_04050_));
 sky130_fd_sc_hd__nor2_2 _09063_ (.A(\core.pipe0_currentInstruction[12] ),
    .B(_04047_),
    .Y(_04051_));
 sky130_fd_sc_hd__or2_2 _09064_ (.A(net1794),
    .B(_04047_),
    .X(_04052_));
 sky130_fd_sc_hd__or2_4 _09065_ (.A(\core.pipe0_currentInstruction[12] ),
    .B(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__and3_4 _09066_ (.A(\core.pipe0_currentInstruction[13] ),
    .B(net1629),
    .C(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__or2_1 _09067_ (.A(\core.pipe0_currentInstruction[6] ),
    .B(_03858_),
    .X(_04055_));
 sky130_fd_sc_hd__or4b_4 _09068_ (.A(net1794),
    .B(_04054_),
    .C(_04055_),
    .D_N(_04050_),
    .X(_04056_));
 sky130_fd_sc_hd__inv_8 _09069_ (.A(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__or4_2 _09070_ (.A(\core.pipe0_currentInstruction[6] ),
    .B(\core.pipe0_currentInstruction[5] ),
    .C(_03858_),
    .D(_03859_),
    .X(_04058_));
 sky130_fd_sc_hd__nor2_4 _09071_ (.A(\core.pipe0_currentInstruction[13] ),
    .B(_04048_),
    .Y(_04059_));
 sky130_fd_sc_hd__or2_4 _09072_ (.A(\core.pipe0_currentInstruction[13] ),
    .B(_04048_),
    .X(_04060_));
 sky130_fd_sc_hd__or4_4 _09073_ (.A(net1751),
    .B(\core.pipe0_currentInstruction[26] ),
    .C(\core.pipe0_currentInstruction[25] ),
    .D(_03868_),
    .X(_04061_));
 sky130_fd_sc_hd__nand2_8 _09074_ (.A(net1794),
    .B(net1629),
    .Y(_04062_));
 sky130_fd_sc_hd__or3_2 _09075_ (.A(_03831_),
    .B(net1634),
    .C(_04061_),
    .X(_04063_));
 sky130_fd_sc_hd__a21o_1 _09076_ (.A1(net1752),
    .A2(_04062_),
    .B1(_04061_),
    .X(_04064_));
 sky130_fd_sc_hd__a21o_4 _09077_ (.A1(_04059_),
    .A2(_04064_),
    .B1(_04058_),
    .X(_04065_));
 sky130_fd_sc_hd__o31a_2 _09078_ (.A1(\core.pipe0_currentInstruction[6] ),
    .A2(\core.pipe0_currentInstruction[5] ),
    .A3(\core.pipe0_currentInstruction[4] ),
    .B1(net1630),
    .X(_04066_));
 sky130_fd_sc_hd__nor3_4 _09079_ (.A(_03858_),
    .B(_04054_),
    .C(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__or3_4 _09080_ (.A(_03858_),
    .B(_04054_),
    .C(_04066_),
    .X(_04068_));
 sky130_fd_sc_hd__nand2_4 _09081_ (.A(_04065_),
    .B(net1150),
    .Y(_04069_));
 sky130_fd_sc_hd__nor2_8 _09082_ (.A(_04057_),
    .B(net1153),
    .Y(_04070_));
 sky130_fd_sc_hd__nand2_8 _09083_ (.A(_04056_),
    .B(_04068_),
    .Y(_04071_));
 sky130_fd_sc_hd__nor2_4 _09084_ (.A(_04057_),
    .B(net1093),
    .Y(_04072_));
 sky130_fd_sc_hd__or2_1 _09085_ (.A(_04057_),
    .B(net1093),
    .X(_04073_));
 sky130_fd_sc_hd__nor2_8 _09086_ (.A(net1705),
    .B(net1633),
    .Y(_04074_));
 sky130_fd_sc_hd__nand2_4 _09087_ (.A(net1763),
    .B(net1629),
    .Y(_04075_));
 sky130_fd_sc_hd__and2_4 _09088_ (.A(net1761),
    .B(net1631),
    .X(_04076_));
 sky130_fd_sc_hd__nand2_8 _09089_ (.A(net1761),
    .B(net1631),
    .Y(_04077_));
 sky130_fd_sc_hd__nor2_1 _09090_ (.A(_03906_),
    .B(net1427),
    .Y(_04078_));
 sky130_fd_sc_hd__nor2_1 _09091_ (.A(_03907_),
    .B(net1431),
    .Y(_04079_));
 sky130_fd_sc_hd__nor2_8 _09092_ (.A(net1684),
    .B(net1633),
    .Y(_04080_));
 sky130_fd_sc_hd__nand2_4 _09093_ (.A(net1777),
    .B(net1631),
    .Y(_04081_));
 sky130_fd_sc_hd__xnor2_1 _09094_ (.A(_03910_),
    .B(net1403),
    .Y(_04082_));
 sky130_fd_sc_hd__nor2_1 _09095_ (.A(net1700),
    .B(net1633),
    .Y(_04083_));
 sky130_fd_sc_hd__nand2_1 _09096_ (.A(net1770),
    .B(net1629),
    .Y(_04084_));
 sky130_fd_sc_hd__xnor2_1 _09097_ (.A(_03911_),
    .B(net1333),
    .Y(_04085_));
 sky130_fd_sc_hd__nor2_8 _09098_ (.A(net1709),
    .B(net1633),
    .Y(_04086_));
 sky130_fd_sc_hd__nand2_8 _09099_ (.A(net1760),
    .B(net1631),
    .Y(_04087_));
 sky130_fd_sc_hd__a221o_1 _09100_ (.A1(_03903_),
    .A2(net1452),
    .B1(net1321),
    .B2(_03904_),
    .C1(_04082_),
    .X(_04088_));
 sky130_fd_sc_hd__o221a_1 _09101_ (.A1(_03903_),
    .A2(net1452),
    .B1(_04087_),
    .B2(_03904_),
    .C1(_04085_),
    .X(_04089_));
 sky130_fd_sc_hd__or4b_4 _09102_ (.A(_04078_),
    .B(_04079_),
    .C(_04088_),
    .D_N(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__a21oi_4 _09103_ (.A1(_03919_),
    .A2(net1189),
    .B1(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__a21o_1 _09104_ (.A1(_03919_),
    .A2(net1189),
    .B1(_04090_),
    .X(_04092_));
 sky130_fd_sc_hd__or2_1 _09105_ (.A(net764),
    .B(net1144),
    .X(_04093_));
 sky130_fd_sc_hd__nand2_1 _09106_ (.A(net1437),
    .B(net1321),
    .Y(_04094_));
 sky130_fd_sc_hd__and4b_4 _09107_ (.A_N(_04094_),
    .B(net1329),
    .C(net1358),
    .D(net1427),
    .X(_04095_));
 sky130_fd_sc_hd__or4_4 _09108_ (.A(net1430),
    .B(net1375),
    .C(net1346),
    .D(_04094_),
    .X(_04096_));
 sky130_fd_sc_hd__a221o_1 _09109_ (.A1(net1690),
    .A2(\core.registers[26][11] ),
    .B1(\core.registers[27][11] ),
    .B2(net1406),
    .C1(net1333),
    .X(_04097_));
 sky130_fd_sc_hd__and3_1 _09110_ (.A(net1777),
    .B(\core.registers[25][11] ),
    .C(net1631),
    .X(_04098_));
 sky130_fd_sc_hd__a211o_1 _09111_ (.A1(\core.registers[24][11] ),
    .A2(net1362),
    .B1(net1349),
    .C1(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__a21bo_1 _09112_ (.A1(_04097_),
    .A2(_04099_),
    .B1_N(net1761),
    .X(_04100_));
 sky130_fd_sc_hd__or2_1 _09113_ (.A(\core.registers[16][11] ),
    .B(net1424),
    .X(_04101_));
 sky130_fd_sc_hd__o211a_1 _09114_ (.A1(\core.registers[17][11] ),
    .A2(net1360),
    .B1(net1337),
    .C1(_04101_),
    .X(_04102_));
 sky130_fd_sc_hd__o221a_1 _09115_ (.A1(net1696),
    .A2(\core.registers[19][11] ),
    .B1(net1424),
    .B2(\core.registers[18][11] ),
    .C1(net1353),
    .X(_04103_));
 sky130_fd_sc_hd__o311a_1 _09116_ (.A1(net1761),
    .A2(_04102_),
    .A3(_04103_),
    .B1(net1706),
    .C1(_04100_),
    .X(_04104_));
 sky130_fd_sc_hd__a221o_1 _09117_ (.A1(net1690),
    .A2(\core.registers[30][11] ),
    .B1(\core.registers[31][11] ),
    .B2(net1404),
    .C1(net1333),
    .X(_04105_));
 sky130_fd_sc_hd__and3_1 _09118_ (.A(net1777),
    .B(\core.registers[29][11] ),
    .C(net1631),
    .X(_04106_));
 sky130_fd_sc_hd__a211o_1 _09119_ (.A1(\core.registers[28][11] ),
    .A2(net1362),
    .B1(net1355),
    .C1(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__a21bo_1 _09120_ (.A1(_04105_),
    .A2(_04107_),
    .B1_N(net1761),
    .X(_04108_));
 sky130_fd_sc_hd__mux2_1 _09121_ (.A0(\core.registers[20][11] ),
    .A1(\core.registers[21][11] ),
    .S(net1424),
    .X(_04109_));
 sky130_fd_sc_hd__o221a_1 _09122_ (.A1(net1696),
    .A2(\core.registers[23][11] ),
    .B1(net1424),
    .B2(\core.registers[22][11] ),
    .C1(net1353),
    .X(_04110_));
 sky130_fd_sc_hd__a211o_1 _09123_ (.A1(net1337),
    .A2(_04109_),
    .B1(_04110_),
    .C1(net1761),
    .X(_04111_));
 sky130_fd_sc_hd__a31o_1 _09124_ (.A1(net1766),
    .A2(_04108_),
    .A3(_04111_),
    .B1(net1322),
    .X(_04112_));
 sky130_fd_sc_hd__a22o_1 _09125_ (.A1(net1696),
    .A2(\core.registers[14][11] ),
    .B1(\core.registers[15][11] ),
    .B2(net1424),
    .X(_04113_));
 sky130_fd_sc_hd__a22o_1 _09126_ (.A1(net1696),
    .A2(\core.registers[10][11] ),
    .B1(\core.registers[11][11] ),
    .B2(net1424),
    .X(_04114_));
 sky130_fd_sc_hd__mux2_1 _09127_ (.A0(_04113_),
    .A1(_04114_),
    .S(net1706),
    .X(_04115_));
 sky130_fd_sc_hd__mux4_1 _09128_ (.A0(\core.registers[8][11] ),
    .A1(\core.registers[9][11] ),
    .A2(\core.registers[12][11] ),
    .A3(\core.registers[13][11] ),
    .S0(net1418),
    .S1(net1766),
    .X(_04116_));
 sky130_fd_sc_hd__mux2_1 _09129_ (.A0(_04115_),
    .A1(_04116_),
    .S(net1337),
    .X(_04117_));
 sky130_fd_sc_hd__mux2_1 _09130_ (.A0(\core.registers[0][11] ),
    .A1(\core.registers[1][11] ),
    .S(net1418),
    .X(_04118_));
 sky130_fd_sc_hd__mux2_1 _09131_ (.A0(\core.registers[4][11] ),
    .A1(\core.registers[5][11] ),
    .S(net1418),
    .X(_04119_));
 sky130_fd_sc_hd__mux2_1 _09132_ (.A0(\core.registers[2][11] ),
    .A1(\core.registers[3][11] ),
    .S(net1424),
    .X(_04120_));
 sky130_fd_sc_hd__mux2_1 _09133_ (.A0(_04118_),
    .A1(_04120_),
    .S(net1353),
    .X(_04121_));
 sky130_fd_sc_hd__mux2_1 _09134_ (.A0(\core.registers[6][11] ),
    .A1(\core.registers[7][11] ),
    .S(net1424),
    .X(_04122_));
 sky130_fd_sc_hd__mux2_1 _09135_ (.A0(_04119_),
    .A1(_04122_),
    .S(net1353),
    .X(_04123_));
 sky130_fd_sc_hd__mux2_1 _09136_ (.A0(_04121_),
    .A1(_04123_),
    .S(net1456),
    .X(_04124_));
 sky130_fd_sc_hd__mux2_1 _09137_ (.A0(_04117_),
    .A1(_04124_),
    .S(net1428),
    .X(_04125_));
 sky130_fd_sc_hd__o22a_2 _09138_ (.A1(_04104_),
    .A2(_04112_),
    .B1(_04125_),
    .B2(net1327),
    .X(_04126_));
 sky130_fd_sc_hd__o211a_4 _09139_ (.A1(net1149),
    .A2(_04126_),
    .B1(net1240),
    .C1(_04093_),
    .X(_04127_));
 sky130_fd_sc_hd__mux2_1 _09140_ (.A0(net1751),
    .A1(_04127_),
    .S(_04072_),
    .X(_04128_));
 sky130_fd_sc_hd__nor2_1 _09141_ (.A(net1263),
    .B(net1039),
    .Y(_04129_));
 sky130_fd_sc_hd__and2_1 _09142_ (.A(net1257),
    .B(_04128_),
    .X(_04130_));
 sky130_fd_sc_hd__nor2_2 _09143_ (.A(_04046_),
    .B(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__and3_2 _09144_ (.A(net1257),
    .B(_04044_),
    .C(_04128_),
    .X(_04132_));
 sky130_fd_sc_hd__nor2_4 _09145_ (.A(_04131_),
    .B(_04132_),
    .Y(_04133_));
 sky130_fd_sc_hd__mux2_8 _09146_ (.A0(net125),
    .A1(net160),
    .S(net1736),
    .X(_04134_));
 sky130_fd_sc_hd__o32a_1 _09147_ (.A1(net1639),
    .A2(net1623),
    .A3(_04134_),
    .B1(net1627),
    .B2(\coreWBInterface.readDataBuffered[26] ),
    .X(_04135_));
 sky130_fd_sc_hd__or2_1 _09148_ (.A(_03986_),
    .B(_04135_),
    .X(_04136_));
 sky130_fd_sc_hd__mux2_8 _09149_ (.A0(net116),
    .A1(net152),
    .S(net1736),
    .X(_04137_));
 sky130_fd_sc_hd__o32a_1 _09150_ (.A1(net1639),
    .A2(net1621),
    .A3(_04137_),
    .B1(net1627),
    .B2(\coreWBInterface.readDataBuffered[18] ),
    .X(_04138_));
 sky130_fd_sc_hd__a21o_1 _09151_ (.A1(net1243),
    .A2(_04138_),
    .B1(_04022_),
    .X(_04139_));
 sky130_fd_sc_hd__a32o_1 _09152_ (.A1(net1458),
    .A2(_04014_),
    .A3(_04136_),
    .B1(_04139_),
    .B2(_04007_),
    .X(_04140_));
 sky130_fd_sc_hd__mux2_4 _09153_ (.A0(net108),
    .A1(net143),
    .S(net1735),
    .X(_04141_));
 sky130_fd_sc_hd__nor2_1 _09154_ (.A(_03989_),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__a2bb2o_1 _09155_ (.A1_N(\coreWBInterface.readDataBuffered[10] ),
    .A2_N(net1627),
    .B1(_04142_),
    .B2(net1745),
    .X(_04143_));
 sky130_fd_sc_hd__or4_1 _09156_ (.A(net1749),
    .B(_03981_),
    .C(_03983_),
    .D(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__o2bb2a_1 _09157_ (.A1_N(_04037_),
    .A2_N(_04144_),
    .B1(_04140_),
    .B2(_04018_),
    .X(_04145_));
 sky130_fd_sc_hd__a221o_1 _09158_ (.A1(\core.pipe1_csrData[10] ),
    .A2(net1249),
    .B1(_03927_),
    .B2(\core.pipe1_resultRegister[10] ),
    .C1(net1244),
    .X(_04146_));
 sky130_fd_sc_hd__a21o_1 _09159_ (.A1(_04029_),
    .A2(_04145_),
    .B1(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__o21a_4 _09160_ (.A1(\core.pipe1_resultRegister[10] ),
    .A2(_03933_),
    .B1(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__mux2_1 _09161_ (.A0(\core.registers[26][10] ),
    .A1(\core.registers[27][10] ),
    .S(net1410),
    .X(_04149_));
 sky130_fd_sc_hd__mux2_1 _09162_ (.A0(\core.registers[24][10] ),
    .A1(\core.registers[25][10] ),
    .S(net1410),
    .X(_04150_));
 sky130_fd_sc_hd__mux2_1 _09163_ (.A0(_04149_),
    .A1(_04150_),
    .S(net1335),
    .X(_04151_));
 sky130_fd_sc_hd__mux2_1 _09164_ (.A0(\core.registers[16][10] ),
    .A1(\core.registers[17][10] ),
    .S(net1412),
    .X(_04152_));
 sky130_fd_sc_hd__o221a_1 _09165_ (.A1(net1692),
    .A2(\core.registers[19][10] ),
    .B1(net1412),
    .B2(\core.registers[18][10] ),
    .C1(net1351),
    .X(_04153_));
 sky130_fd_sc_hd__a21o_1 _09166_ (.A1(net1335),
    .A2(_04152_),
    .B1(_04153_),
    .X(_04154_));
 sky130_fd_sc_hd__mux2_1 _09167_ (.A0(\core.registers[30][10] ),
    .A1(\core.registers[31][10] ),
    .S(net1411),
    .X(_04155_));
 sky130_fd_sc_hd__mux2_1 _09168_ (.A0(\core.registers[28][10] ),
    .A1(\core.registers[29][10] ),
    .S(net1410),
    .X(_04156_));
 sky130_fd_sc_hd__mux2_1 _09169_ (.A0(_04155_),
    .A1(_04156_),
    .S(net1335),
    .X(_04157_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(\core.registers[20][10] ),
    .A1(\core.registers[21][10] ),
    .S(net1413),
    .X(_04158_));
 sky130_fd_sc_hd__o221a_1 _09171_ (.A1(net1692),
    .A2(\core.registers[23][10] ),
    .B1(net1412),
    .B2(\core.registers[22][10] ),
    .C1(net1351),
    .X(_04159_));
 sky130_fd_sc_hd__a21o_1 _09172_ (.A1(net1335),
    .A2(_04158_),
    .B1(_04159_),
    .X(_04160_));
 sky130_fd_sc_hd__mux4_2 _09173_ (.A0(_04154_),
    .A1(_04160_),
    .A2(_04151_),
    .A3(_04157_),
    .S0(net1766),
    .S1(net1761),
    .X(_04161_));
 sky130_fd_sc_hd__a22o_1 _09174_ (.A1(net1691),
    .A2(\core.registers[14][10] ),
    .B1(\core.registers[15][10] ),
    .B2(net1411),
    .X(_04162_));
 sky130_fd_sc_hd__a22o_1 _09175_ (.A1(net1691),
    .A2(\core.registers[10][10] ),
    .B1(\core.registers[11][10] ),
    .B2(net1410),
    .X(_04163_));
 sky130_fd_sc_hd__mux2_1 _09176_ (.A0(_04162_),
    .A1(_04163_),
    .S(net1706),
    .X(_04164_));
 sky130_fd_sc_hd__mux4_1 _09177_ (.A0(\core.registers[8][10] ),
    .A1(\core.registers[9][10] ),
    .A2(\core.registers[12][10] ),
    .A3(\core.registers[13][10] ),
    .S0(net1411),
    .S1(net1765),
    .X(_04165_));
 sky130_fd_sc_hd__mux2_1 _09178_ (.A0(_04164_),
    .A1(_04165_),
    .S(net1335),
    .X(_04166_));
 sky130_fd_sc_hd__or2_1 _09179_ (.A(\core.registers[0][10] ),
    .B(net1412),
    .X(_04167_));
 sky130_fd_sc_hd__o211a_1 _09180_ (.A1(\core.registers[1][10] ),
    .A2(net1361),
    .B1(_04167_),
    .C1(net1443),
    .X(_04168_));
 sky130_fd_sc_hd__mux2_1 _09181_ (.A0(\core.registers[4][10] ),
    .A1(\core.registers[5][10] ),
    .S(net1413),
    .X(_04169_));
 sky130_fd_sc_hd__a211o_1 _09182_ (.A1(net1457),
    .A2(_04169_),
    .B1(_04168_),
    .C1(net1351),
    .X(_04170_));
 sky130_fd_sc_hd__o221a_1 _09183_ (.A1(net1693),
    .A2(\core.registers[7][10] ),
    .B1(net1413),
    .B2(\core.registers[6][10] ),
    .C1(net1454),
    .X(_04171_));
 sky130_fd_sc_hd__o221a_1 _09184_ (.A1(net1693),
    .A2(\core.registers[3][10] ),
    .B1(net1413),
    .B2(\core.registers[2][10] ),
    .C1(net1443),
    .X(_04172_));
 sky130_fd_sc_hd__o31a_1 _09185_ (.A1(net1336),
    .A2(_04171_),
    .A3(_04172_),
    .B1(net1428),
    .X(_04173_));
 sky130_fd_sc_hd__and2_1 _09186_ (.A(_04170_),
    .B(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__a21o_1 _09187_ (.A1(net1433),
    .A2(_04166_),
    .B1(net1326),
    .X(_04175_));
 sky130_fd_sc_hd__o22a_4 _09188_ (.A1(net1322),
    .A2(_04161_),
    .B1(_04174_),
    .B2(_04175_),
    .X(_04176_));
 sky130_fd_sc_hd__o21a_1 _09189_ (.A1(net1148),
    .A2(_04176_),
    .B1(net1240),
    .X(_04177_));
 sky130_fd_sc_hd__o21ai_4 _09190_ (.A1(net1144),
    .A2(net758),
    .B1(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__nor2_1 _09191_ (.A(net1752),
    .B(net1042),
    .Y(_04179_));
 sky130_fd_sc_hd__a211o_2 _09192_ (.A1(net1042),
    .A2(_04178_),
    .B1(_04179_),
    .C1(net1265),
    .X(_04180_));
 sky130_fd_sc_hd__or2_4 _09193_ (.A(net451),
    .B(net1261),
    .X(_04181_));
 sky130_fd_sc_hd__a221o_1 _09194_ (.A1(net1656),
    .A2(\core.registers[30][10] ),
    .B1(\core.registers[31][10] ),
    .B2(net1509),
    .C1(net1664),
    .X(_04182_));
 sky130_fd_sc_hd__mux2_1 _09195_ (.A0(\core.registers[28][10] ),
    .A1(\core.registers[29][10] ),
    .S(net1508),
    .X(_04183_));
 sky130_fd_sc_hd__o21a_1 _09196_ (.A1(net1792),
    .A2(_04183_),
    .B1(_04182_),
    .X(_04184_));
 sky130_fd_sc_hd__mux2_1 _09197_ (.A0(\core.registers[8][10] ),
    .A1(\core.registers[9][10] ),
    .S(net1509),
    .X(_04185_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(\core.registers[10][10] ),
    .A1(\core.registers[11][10] ),
    .S(net1508),
    .X(_04186_));
 sky130_fd_sc_hd__mux2_1 _09199_ (.A0(\core.registers[24][10] ),
    .A1(\core.registers[25][10] ),
    .S(net1508),
    .X(_04187_));
 sky130_fd_sc_hd__a221o_1 _09200_ (.A1(net1655),
    .A2(\core.registers[26][10] ),
    .B1(\core.registers[27][10] ),
    .B2(net1508),
    .C1(net1664),
    .X(_04188_));
 sky130_fd_sc_hd__mux2_1 _09201_ (.A0(_04185_),
    .A1(_04186_),
    .S(net1555),
    .X(_04189_));
 sky130_fd_sc_hd__o21ai_1 _09202_ (.A1(net1790),
    .A2(_04187_),
    .B1(_04188_),
    .Y(_04190_));
 sky130_fd_sc_hd__nand2_1 _09203_ (.A(net1781),
    .B(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__o211a_1 _09204_ (.A1(net1781),
    .A2(_04189_),
    .B1(_04191_),
    .C1(net1670),
    .X(_04192_));
 sky130_fd_sc_hd__mux2_1 _09205_ (.A0(\core.registers[12][10] ),
    .A1(\core.registers[13][10] ),
    .S(net1509),
    .X(_04193_));
 sky130_fd_sc_hd__mux2_1 _09206_ (.A0(\core.registers[14][10] ),
    .A1(\core.registers[15][10] ),
    .S(net1509),
    .X(_04194_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(_04193_),
    .A1(_04194_),
    .S(net1555),
    .X(_04195_));
 sky130_fd_sc_hd__mux2_1 _09208_ (.A0(_04184_),
    .A1(_04195_),
    .S(net1672),
    .X(_04196_));
 sky130_fd_sc_hd__a211o_1 _09209_ (.A1(net1785),
    .A2(_04196_),
    .B1(_04192_),
    .C1(net1564),
    .X(_04197_));
 sky130_fd_sc_hd__mux2_1 _09210_ (.A0(\core.registers[18][10] ),
    .A1(\core.registers[19][10] ),
    .S(net1511),
    .X(_04198_));
 sky130_fd_sc_hd__mux2_1 _09211_ (.A0(\core.registers[16][10] ),
    .A1(\core.registers[17][10] ),
    .S(net1511),
    .X(_04199_));
 sky130_fd_sc_hd__mux2_1 _09212_ (.A0(_04198_),
    .A1(_04199_),
    .S(net1536),
    .X(_04200_));
 sky130_fd_sc_hd__o221a_1 _09213_ (.A1(net1656),
    .A2(\core.registers[23][10] ),
    .B1(net1511),
    .B2(\core.registers[22][10] ),
    .C1(net1556),
    .X(_04201_));
 sky130_fd_sc_hd__mux2_1 _09214_ (.A0(\core.registers[20][10] ),
    .A1(\core.registers[21][10] ),
    .S(net1512),
    .X(_04202_));
 sky130_fd_sc_hd__mux2_1 _09215_ (.A0(\core.registers[0][10] ),
    .A1(\core.registers[1][10] ),
    .S(net1511),
    .X(_04203_));
 sky130_fd_sc_hd__mux2_1 _09216_ (.A0(\core.registers[2][10] ),
    .A1(\core.registers[3][10] ),
    .S(net1512),
    .X(_04204_));
 sky130_fd_sc_hd__mux2_1 _09217_ (.A0(_04203_),
    .A1(_04204_),
    .S(net1556),
    .X(_04205_));
 sky130_fd_sc_hd__mux2_1 _09218_ (.A0(\core.registers[4][10] ),
    .A1(\core.registers[5][10] ),
    .S(net1512),
    .X(_04206_));
 sky130_fd_sc_hd__o221a_1 _09219_ (.A1(net1657),
    .A2(\core.registers[7][10] ),
    .B1(net1512),
    .B2(\core.registers[6][10] ),
    .C1(net1556),
    .X(_04207_));
 sky130_fd_sc_hd__a211o_1 _09220_ (.A1(net1537),
    .A2(_04206_),
    .B1(_04207_),
    .C1(net1580),
    .X(_04208_));
 sky130_fd_sc_hd__a211o_1 _09221_ (.A1(net1536),
    .A2(_04202_),
    .B1(_04201_),
    .C1(net1580),
    .X(_04209_));
 sky130_fd_sc_hd__o211a_1 _09222_ (.A1(net1589),
    .A2(_04200_),
    .B1(_04209_),
    .C1(net1599),
    .X(_04210_));
 sky130_fd_sc_hd__o211a_2 _09223_ (.A1(net1589),
    .A2(_04205_),
    .B1(_04208_),
    .C1(net1595),
    .X(_04211_));
 sky130_fd_sc_hd__o31a_4 _09224_ (.A1(net1568),
    .A2(_04210_),
    .A3(_04211_),
    .B1(_04197_),
    .X(_04212_));
 sky130_fd_sc_hd__a22o_4 _09225_ (.A1(net1095),
    .A2(net758),
    .B1(_04212_),
    .B2(net1046),
    .X(_04213_));
 sky130_fd_sc_hd__o21a_4 _09226_ (.A1(net1265),
    .A2(_04213_),
    .B1(_04181_),
    .X(_04214_));
 sky130_fd_sc_hd__o21ai_4 _09227_ (.A1(net1265),
    .A2(_04213_),
    .B1(_04181_),
    .Y(_04215_));
 sky130_fd_sc_hd__nor2_1 _09228_ (.A(_04180_),
    .B(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__nand2_2 _09229_ (.A(_04180_),
    .B(_04215_),
    .Y(_04217_));
 sky130_fd_sc_hd__nand2b_4 _09230_ (.A_N(_04216_),
    .B(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__mux2_8 _09231_ (.A0(net124),
    .A1(net159),
    .S(net1737),
    .X(_04219_));
 sky130_fd_sc_hd__nor2_1 _09232_ (.A(net1623),
    .B(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__a2bb2o_1 _09233_ (.A1_N(\coreWBInterface.readDataBuffered[25] ),
    .A2_N(net1626),
    .B1(_04220_),
    .B2(net1745),
    .X(_04221_));
 sky130_fd_sc_hd__nand2b_1 _09234_ (.A_N(_03986_),
    .B(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__mux2_4 _09235_ (.A0(net115),
    .A1(net150),
    .S(net1736),
    .X(_04223_));
 sky130_fd_sc_hd__nor2_1 _09236_ (.A(net1621),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__a2bb2o_1 _09237_ (.A1_N(\coreWBInterface.readDataBuffered[17] ),
    .A2_N(net1626),
    .B1(_04224_),
    .B2(net1745),
    .X(_04225_));
 sky130_fd_sc_hd__inv_2 _09238_ (.A(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__a21o_1 _09239_ (.A1(_04021_),
    .A2(_04226_),
    .B1(_04022_),
    .X(_04227_));
 sky130_fd_sc_hd__a31o_1 _09240_ (.A1(net1458),
    .A2(_04014_),
    .A3(_04222_),
    .B1(_04018_),
    .X(_04228_));
 sky130_fd_sc_hd__a21oi_1 _09241_ (.A1(_04007_),
    .A2(_04227_),
    .B1(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__mux2_4 _09242_ (.A0(net170),
    .A1(net142),
    .S(net1734),
    .X(_04230_));
 sky130_fd_sc_hd__nor2_1 _09243_ (.A(_03989_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__a2bb2o_1 _09244_ (.A1_N(\coreWBInterface.readDataBuffered[9] ),
    .A2_N(net1627),
    .B1(_04231_),
    .B2(net1745),
    .X(_04232_));
 sky130_fd_sc_hd__or4_2 _09245_ (.A(net1749),
    .B(_03981_),
    .C(_03983_),
    .D(_04232_),
    .X(_04233_));
 sky130_fd_sc_hd__a211o_1 _09246_ (.A1(_04037_),
    .A2(_04233_),
    .B1(_04229_),
    .C1(net1242),
    .X(_04234_));
 sky130_fd_sc_hd__a221oi_1 _09247_ (.A1(\core.pipe1_csrData[9] ),
    .A2(net1249),
    .B1(_03927_),
    .B2(\core.pipe1_resultRegister[9] ),
    .C1(net1244),
    .Y(_04235_));
 sky130_fd_sc_hd__o2bb2a_1 _09248_ (.A1_N(_04235_),
    .A2_N(_04234_),
    .B1(_03933_),
    .B2(\core.pipe1_resultRegister[9] ),
    .X(_04236_));
 sky130_fd_sc_hd__mux2_1 _09249_ (.A0(\core.registers[26][9] ),
    .A1(\core.registers[27][9] ),
    .S(net1419),
    .X(_04237_));
 sky130_fd_sc_hd__mux2_1 _09250_ (.A0(\core.registers[24][9] ),
    .A1(\core.registers[25][9] ),
    .S(net1418),
    .X(_04238_));
 sky130_fd_sc_hd__mux2_1 _09251_ (.A0(_04237_),
    .A1(_04238_),
    .S(net1338),
    .X(_04239_));
 sky130_fd_sc_hd__mux2_1 _09252_ (.A0(\core.registers[16][9] ),
    .A1(\core.registers[17][9] ),
    .S(net1419),
    .X(_04240_));
 sky130_fd_sc_hd__o221a_1 _09253_ (.A1(net1698),
    .A2(\core.registers[19][9] ),
    .B1(net1418),
    .B2(\core.registers[18][9] ),
    .C1(net1353),
    .X(_04241_));
 sky130_fd_sc_hd__a21o_1 _09254_ (.A1(net1338),
    .A2(_04240_),
    .B1(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__mux2_1 _09255_ (.A0(\core.registers[30][9] ),
    .A1(\core.registers[31][9] ),
    .S(net1416),
    .X(_04243_));
 sky130_fd_sc_hd__mux2_1 _09256_ (.A0(\core.registers[28][9] ),
    .A1(\core.registers[29][9] ),
    .S(net1417),
    .X(_04244_));
 sky130_fd_sc_hd__mux2_1 _09257_ (.A0(_04243_),
    .A1(_04244_),
    .S(net1338),
    .X(_04245_));
 sky130_fd_sc_hd__mux2_1 _09258_ (.A0(\core.registers[20][9] ),
    .A1(\core.registers[21][9] ),
    .S(net1418),
    .X(_04246_));
 sky130_fd_sc_hd__o221a_1 _09259_ (.A1(net1698),
    .A2(\core.registers[23][9] ),
    .B1(net1418),
    .B2(\core.registers[22][9] ),
    .C1(net1354),
    .X(_04247_));
 sky130_fd_sc_hd__a21o_1 _09260_ (.A1(net1338),
    .A2(_04246_),
    .B1(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__mux4_1 _09261_ (.A0(_04242_),
    .A1(_04248_),
    .A2(_04239_),
    .A3(_04245_),
    .S0(net1766),
    .S1(net1761),
    .X(_04249_));
 sky130_fd_sc_hd__a22o_1 _09262_ (.A1(net1698),
    .A2(\core.registers[14][9] ),
    .B1(\core.registers[15][9] ),
    .B2(net1419),
    .X(_04250_));
 sky130_fd_sc_hd__a22o_1 _09263_ (.A1(net1698),
    .A2(\core.registers[10][9] ),
    .B1(\core.registers[11][9] ),
    .B2(net1419),
    .X(_04251_));
 sky130_fd_sc_hd__mux2_1 _09264_ (.A0(_04250_),
    .A1(_04251_),
    .S(net1706),
    .X(_04252_));
 sky130_fd_sc_hd__mux4_1 _09265_ (.A0(\core.registers[8][9] ),
    .A1(\core.registers[9][9] ),
    .A2(\core.registers[12][9] ),
    .A3(\core.registers[13][9] ),
    .S0(net1419),
    .S1(net1766),
    .X(_04253_));
 sky130_fd_sc_hd__mux2_1 _09266_ (.A0(_04252_),
    .A1(_04253_),
    .S(net1338),
    .X(_04254_));
 sky130_fd_sc_hd__or2_1 _09267_ (.A(\core.registers[0][9] ),
    .B(net1418),
    .X(_04255_));
 sky130_fd_sc_hd__o211a_1 _09268_ (.A1(\core.registers[1][9] ),
    .A2(net1360),
    .B1(_04255_),
    .C1(net1445),
    .X(_04256_));
 sky130_fd_sc_hd__mux2_1 _09269_ (.A0(\core.registers[4][9] ),
    .A1(\core.registers[5][9] ),
    .S(net1418),
    .X(_04257_));
 sky130_fd_sc_hd__a211o_1 _09270_ (.A1(net1456),
    .A2(_04257_),
    .B1(_04256_),
    .C1(net1354),
    .X(_04258_));
 sky130_fd_sc_hd__o221a_1 _09271_ (.A1(net1698),
    .A2(\core.registers[7][9] ),
    .B1(net1418),
    .B2(\core.registers[6][9] ),
    .C1(net1456),
    .X(_04259_));
 sky130_fd_sc_hd__o221a_1 _09272_ (.A1(net1698),
    .A2(\core.registers[3][9] ),
    .B1(net1419),
    .B2(\core.registers[2][9] ),
    .C1(net1445),
    .X(_04260_));
 sky130_fd_sc_hd__o31a_1 _09273_ (.A1(net1338),
    .A2(_04259_),
    .A3(_04260_),
    .B1(net1428),
    .X(_04261_));
 sky130_fd_sc_hd__and2_1 _09274_ (.A(_04258_),
    .B(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__a21o_1 _09275_ (.A1(net1433),
    .A2(_04254_),
    .B1(net1326),
    .X(_04263_));
 sky130_fd_sc_hd__o22a_2 _09276_ (.A1(net1322),
    .A2(_04249_),
    .B1(_04262_),
    .B2(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__o21a_1 _09277_ (.A1(net1149),
    .A2(_04264_),
    .B1(net1240),
    .X(_04265_));
 sky130_fd_sc_hd__o21ai_4 _09278_ (.A1(net1144),
    .A2(net903),
    .B1(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__nor2_1 _09279_ (.A(\core.pipe0_currentInstruction[29] ),
    .B(net1042),
    .Y(_04267_));
 sky130_fd_sc_hd__a211o_2 _09280_ (.A1(net1042),
    .A2(_04266_),
    .B1(_04267_),
    .C1(net1265),
    .X(_04268_));
 sky130_fd_sc_hd__nand2_2 _09281_ (.A(_03825_),
    .B(net1266),
    .Y(_04269_));
 sky130_fd_sc_hd__mux2_1 _09282_ (.A0(\core.registers[24][9] ),
    .A1(\core.registers[25][9] ),
    .S(net1517),
    .X(_04270_));
 sky130_fd_sc_hd__a221o_1 _09283_ (.A1(net1661),
    .A2(\core.registers[26][9] ),
    .B1(\core.registers[27][9] ),
    .B2(net1518),
    .C1(net1665),
    .X(_04271_));
 sky130_fd_sc_hd__o211a_1 _09284_ (.A1(net1792),
    .A2(_04270_),
    .B1(_04271_),
    .C1(net1783),
    .X(_04272_));
 sky130_fd_sc_hd__and3_1 _09285_ (.A(net1793),
    .B(\core.registers[9][9] ),
    .C(net1631),
    .X(_04273_));
 sky130_fd_sc_hd__a211o_1 _09286_ (.A1(\core.registers[8][9] ),
    .A2(net1461),
    .B1(_04273_),
    .C1(net1559),
    .X(_04274_));
 sky130_fd_sc_hd__mux2_1 _09287_ (.A0(\core.registers[10][9] ),
    .A1(\core.registers[11][9] ),
    .S(net1518),
    .X(_04275_));
 sky130_fd_sc_hd__o211a_1 _09288_ (.A1(net1540),
    .A2(_04275_),
    .B1(_04274_),
    .C1(net1672),
    .X(_04276_));
 sky130_fd_sc_hd__o21a_1 _09289_ (.A1(_04272_),
    .A2(_04276_),
    .B1(net1671),
    .X(_04277_));
 sky130_fd_sc_hd__mux2_1 _09290_ (.A0(\core.registers[28][9] ),
    .A1(\core.registers[29][9] ),
    .S(net1516),
    .X(_04278_));
 sky130_fd_sc_hd__a221o_1 _09291_ (.A1(net1661),
    .A2(\core.registers[30][9] ),
    .B1(\core.registers[31][9] ),
    .B2(net1516),
    .C1(net1665),
    .X(_04279_));
 sky130_fd_sc_hd__o21a_1 _09292_ (.A1(net1792),
    .A2(_04278_),
    .B1(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__mux2_1 _09293_ (.A0(\core.registers[12][9] ),
    .A1(\core.registers[13][9] ),
    .S(net1518),
    .X(_04281_));
 sky130_fd_sc_hd__mux2_1 _09294_ (.A0(\core.registers[14][9] ),
    .A1(\core.registers[15][9] ),
    .S(net1518),
    .X(_04282_));
 sky130_fd_sc_hd__mux2_1 _09295_ (.A0(_04281_),
    .A1(_04282_),
    .S(net1559),
    .X(_04283_));
 sky130_fd_sc_hd__mux2_1 _09296_ (.A0(_04280_),
    .A1(_04283_),
    .S(net1673),
    .X(_04284_));
 sky130_fd_sc_hd__a211o_1 _09297_ (.A1(net1786),
    .A2(_04284_),
    .B1(_04277_),
    .C1(net1564),
    .X(_04285_));
 sky130_fd_sc_hd__mux2_1 _09298_ (.A0(\core.registers[18][9] ),
    .A1(\core.registers[19][9] ),
    .S(net1517),
    .X(_04286_));
 sky130_fd_sc_hd__mux2_1 _09299_ (.A0(\core.registers[16][9] ),
    .A1(\core.registers[17][9] ),
    .S(net1517),
    .X(_04287_));
 sky130_fd_sc_hd__mux2_1 _09300_ (.A0(_04286_),
    .A1(_04287_),
    .S(net1540),
    .X(_04288_));
 sky130_fd_sc_hd__o221a_1 _09301_ (.A1(net1661),
    .A2(\core.registers[23][9] ),
    .B1(net1517),
    .B2(\core.registers[22][9] ),
    .C1(net1559),
    .X(_04289_));
 sky130_fd_sc_hd__mux2_1 _09302_ (.A0(\core.registers[20][9] ),
    .A1(\core.registers[21][9] ),
    .S(net1518),
    .X(_04290_));
 sky130_fd_sc_hd__mux2_1 _09303_ (.A0(\core.registers[0][9] ),
    .A1(\core.registers[1][9] ),
    .S(net1517),
    .X(_04291_));
 sky130_fd_sc_hd__mux2_1 _09304_ (.A0(\core.registers[2][9] ),
    .A1(\core.registers[3][9] ),
    .S(net1517),
    .X(_04292_));
 sky130_fd_sc_hd__mux2_1 _09305_ (.A0(_04291_),
    .A1(_04292_),
    .S(net1559),
    .X(_04293_));
 sky130_fd_sc_hd__mux2_1 _09306_ (.A0(\core.registers[4][9] ),
    .A1(\core.registers[5][9] ),
    .S(net1517),
    .X(_04294_));
 sky130_fd_sc_hd__o221a_1 _09307_ (.A1(net1661),
    .A2(\core.registers[7][9] ),
    .B1(net1517),
    .B2(\core.registers[6][9] ),
    .C1(net1559),
    .X(_04295_));
 sky130_fd_sc_hd__a211o_1 _09308_ (.A1(net1540),
    .A2(_04294_),
    .B1(_04295_),
    .C1(net1579),
    .X(_04296_));
 sky130_fd_sc_hd__a211o_1 _09309_ (.A1(net1540),
    .A2(_04290_),
    .B1(_04289_),
    .C1(net1579),
    .X(_04297_));
 sky130_fd_sc_hd__o211a_1 _09310_ (.A1(net1591),
    .A2(_04288_),
    .B1(_04297_),
    .C1(net1599),
    .X(_04298_));
 sky130_fd_sc_hd__o211a_1 _09311_ (.A1(net1591),
    .A2(_04293_),
    .B1(_04296_),
    .C1(net1595),
    .X(_04299_));
 sky130_fd_sc_hd__o31a_2 _09312_ (.A1(net1568),
    .A2(_04298_),
    .A3(_04299_),
    .B1(_04285_),
    .X(_04300_));
 sky130_fd_sc_hd__a22o_4 _09313_ (.A1(net1095),
    .A2(net903),
    .B1(_04300_),
    .B2(net1046),
    .X(_04301_));
 sky130_fd_sc_hd__o21ai_4 _09314_ (.A1(net1265),
    .A2(_04301_),
    .B1(_04269_),
    .Y(_04302_));
 sky130_fd_sc_hd__inv_2 _09315_ (.A(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__or2_2 _09316_ (.A(_04268_),
    .B(_04302_),
    .X(_04304_));
 sky130_fd_sc_hd__nand2_2 _09317_ (.A(_04268_),
    .B(_04302_),
    .Y(_04305_));
 sky130_fd_sc_hd__nand2_2 _09318_ (.A(_04304_),
    .B(_04305_),
    .Y(_04306_));
 sky130_fd_sc_hd__inv_2 _09319_ (.A(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__mux2_8 _09320_ (.A0(net123),
    .A1(net158),
    .S(net1737),
    .X(_04308_));
 sky130_fd_sc_hd__o32a_2 _09321_ (.A1(net1639),
    .A2(net1623),
    .A3(_04308_),
    .B1(net1627),
    .B2(\coreWBInterface.readDataBuffered[24] ),
    .X(_04309_));
 sky130_fd_sc_hd__or2_1 _09322_ (.A(_03986_),
    .B(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__mux2_8 _09323_ (.A0(net114),
    .A1(net149),
    .S(net1736),
    .X(_04311_));
 sky130_fd_sc_hd__o32a_1 _09324_ (.A1(net1640),
    .A2(net1621),
    .A3(_04311_),
    .B1(net1626),
    .B2(\coreWBInterface.readDataBuffered[16] ),
    .X(_04312_));
 sky130_fd_sc_hd__and4_1 _09325_ (.A(_03982_),
    .B(_04017_),
    .C(_04020_),
    .D(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__nor2_1 _09326_ (.A(_04022_),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__a31o_1 _09327_ (.A1(net1458),
    .A2(_04014_),
    .A3(_04310_),
    .B1(_04018_),
    .X(_04315_));
 sky130_fd_sc_hd__o21ba_1 _09328_ (.A1(_04008_),
    .A2(_04314_),
    .B1_N(_04315_),
    .X(_04316_));
 sky130_fd_sc_hd__mux2_8 _09329_ (.A0(net169),
    .A1(net141),
    .S(net1734),
    .X(_04317_));
 sky130_fd_sc_hd__o32a_1 _09330_ (.A1(net1639),
    .A2(_03989_),
    .A3(_04317_),
    .B1(net1627),
    .B2(\coreWBInterface.readDataBuffered[8] ),
    .X(_04318_));
 sky130_fd_sc_hd__nand2_1 _09331_ (.A(_04031_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__a211o_1 _09332_ (.A1(_04037_),
    .A2(_04319_),
    .B1(_04316_),
    .C1(net1242),
    .X(_04320_));
 sky130_fd_sc_hd__a221oi_4 _09333_ (.A1(\core.pipe1_csrData[8] ),
    .A2(net1249),
    .B1(_03927_),
    .B2(\core.pipe1_resultRegister[8] ),
    .C1(net1244),
    .Y(_04321_));
 sky130_fd_sc_hd__o2bb2a_4 _09334_ (.A1_N(_04321_),
    .A2_N(_04320_),
    .B1(_03933_),
    .B2(\core.pipe1_resultRegister[8] ),
    .X(_04322_));
 sky130_fd_sc_hd__mux2_1 _09335_ (.A0(\core.registers[26][8] ),
    .A1(\core.registers[27][8] ),
    .S(net1400),
    .X(_04323_));
 sky130_fd_sc_hd__mux2_1 _09336_ (.A0(\core.registers[24][8] ),
    .A1(\core.registers[25][8] ),
    .S(net1400),
    .X(_04324_));
 sky130_fd_sc_hd__mux2_1 _09337_ (.A0(_04323_),
    .A1(_04324_),
    .S(net1334),
    .X(_04325_));
 sky130_fd_sc_hd__mux2_1 _09338_ (.A0(\core.registers[16][8] ),
    .A1(\core.registers[17][8] ),
    .S(net1411),
    .X(_04326_));
 sky130_fd_sc_hd__o221a_1 _09339_ (.A1(net1695),
    .A2(\core.registers[19][8] ),
    .B1(net1411),
    .B2(\core.registers[18][8] ),
    .C1(net1350),
    .X(_04327_));
 sky130_fd_sc_hd__a21o_1 _09340_ (.A1(net1335),
    .A2(_04326_),
    .B1(_04327_),
    .X(_04328_));
 sky130_fd_sc_hd__mux2_1 _09341_ (.A0(\core.registers[30][8] ),
    .A1(\core.registers[31][8] ),
    .S(net1410),
    .X(_04329_));
 sky130_fd_sc_hd__mux2_1 _09342_ (.A0(\core.registers[28][8] ),
    .A1(\core.registers[29][8] ),
    .S(net1410),
    .X(_04330_));
 sky130_fd_sc_hd__mux2_1 _09343_ (.A0(_04329_),
    .A1(_04330_),
    .S(net1335),
    .X(_04331_));
 sky130_fd_sc_hd__mux2_1 _09344_ (.A0(\core.registers[20][8] ),
    .A1(\core.registers[21][8] ),
    .S(net1411),
    .X(_04332_));
 sky130_fd_sc_hd__o221a_1 _09345_ (.A1(net1691),
    .A2(\core.registers[23][8] ),
    .B1(net1411),
    .B2(\core.registers[22][8] ),
    .C1(net1350),
    .X(_04333_));
 sky130_fd_sc_hd__a21o_1 _09346_ (.A1(net1335),
    .A2(_04332_),
    .B1(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__mux4_1 _09347_ (.A0(_04328_),
    .A1(_04334_),
    .A2(_04325_),
    .A3(_04331_),
    .S0(net1765),
    .S1(net1761),
    .X(_04335_));
 sky130_fd_sc_hd__a22o_1 _09348_ (.A1(net1689),
    .A2(\core.registers[14][8] ),
    .B1(\core.registers[15][8] ),
    .B2(net1410),
    .X(_04336_));
 sky130_fd_sc_hd__a22o_1 _09349_ (.A1(net1689),
    .A2(\core.registers[10][8] ),
    .B1(\core.registers[11][8] ),
    .B2(net1417),
    .X(_04337_));
 sky130_fd_sc_hd__mux2_1 _09350_ (.A0(_04336_),
    .A1(_04337_),
    .S(net1707),
    .X(_04338_));
 sky130_fd_sc_hd__mux4_1 _09351_ (.A0(\core.registers[8][8] ),
    .A1(\core.registers[9][8] ),
    .A2(\core.registers[12][8] ),
    .A3(\core.registers[13][8] ),
    .S0(net1410),
    .S1(net1765),
    .X(_04339_));
 sky130_fd_sc_hd__mux2_1 _09352_ (.A0(_04338_),
    .A1(_04339_),
    .S(net1338),
    .X(_04340_));
 sky130_fd_sc_hd__or2_1 _09353_ (.A(\core.registers[0][8] ),
    .B(net1416),
    .X(_04341_));
 sky130_fd_sc_hd__o211a_1 _09354_ (.A1(\core.registers[1][8] ),
    .A2(net1361),
    .B1(_04341_),
    .C1(net1443),
    .X(_04342_));
 sky130_fd_sc_hd__mux2_1 _09355_ (.A0(\core.registers[4][8] ),
    .A1(\core.registers[5][8] ),
    .S(net1416),
    .X(_04343_));
 sky130_fd_sc_hd__a211o_1 _09356_ (.A1(net1454),
    .A2(_04343_),
    .B1(_04342_),
    .C1(net1352),
    .X(_04344_));
 sky130_fd_sc_hd__o221a_1 _09357_ (.A1(net1692),
    .A2(\core.registers[7][8] ),
    .B1(net1412),
    .B2(\core.registers[6][8] ),
    .C1(net1454),
    .X(_04345_));
 sky130_fd_sc_hd__o221a_1 _09358_ (.A1(net1692),
    .A2(\core.registers[3][8] ),
    .B1(net1412),
    .B2(\core.registers[2][8] ),
    .C1(net1443),
    .X(_04346_));
 sky130_fd_sc_hd__o31a_1 _09359_ (.A1(net1336),
    .A2(_04345_),
    .A3(_04346_),
    .B1(net1428),
    .X(_04347_));
 sky130_fd_sc_hd__and2_1 _09360_ (.A(_04344_),
    .B(_04347_),
    .X(_04348_));
 sky130_fd_sc_hd__a21o_1 _09361_ (.A1(net1433),
    .A2(_04340_),
    .B1(net1326),
    .X(_04349_));
 sky130_fd_sc_hd__o22a_2 _09362_ (.A1(net1322),
    .A2(_04335_),
    .B1(_04348_),
    .B2(_04349_),
    .X(_04350_));
 sky130_fd_sc_hd__o21a_1 _09363_ (.A1(net1149),
    .A2(_04350_),
    .B1(net1241),
    .X(_04351_));
 sky130_fd_sc_hd__o21ai_4 _09364_ (.A1(net1144),
    .A2(_04322_),
    .B1(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__and2_2 _09365_ (.A(net1042),
    .B(_04352_),
    .X(_04353_));
 sky130_fd_sc_hd__o21ai_4 _09366_ (.A1(\core.pipe0_currentInstruction[28] ),
    .A2(_04072_),
    .B1(net1261),
    .Y(_04354_));
 sky130_fd_sc_hd__or2_2 _09367_ (.A(net480),
    .B(net1261),
    .X(_04355_));
 sky130_fd_sc_hd__mux2_1 _09368_ (.A0(\core.registers[28][8] ),
    .A1(\core.registers[29][8] ),
    .S(net1508),
    .X(_04356_));
 sky130_fd_sc_hd__a221o_1 _09369_ (.A1(net1656),
    .A2(\core.registers[30][8] ),
    .B1(\core.registers[31][8] ),
    .B2(net1508),
    .C1(net1664),
    .X(_04357_));
 sky130_fd_sc_hd__mux2_1 _09370_ (.A0(\core.registers[24][8] ),
    .A1(\core.registers[25][8] ),
    .S(net1497),
    .X(_04358_));
 sky130_fd_sc_hd__a221o_1 _09371_ (.A1(net1651),
    .A2(\core.registers[26][8] ),
    .B1(\core.registers[27][8] ),
    .B2(net1497),
    .C1(net1664),
    .X(_04359_));
 sky130_fd_sc_hd__mux2_1 _09372_ (.A0(\core.registers[8][8] ),
    .A1(\core.registers[9][8] ),
    .S(net1515),
    .X(_04360_));
 sky130_fd_sc_hd__mux2_1 _09373_ (.A0(\core.registers[10][8] ),
    .A1(\core.registers[11][8] ),
    .S(net1515),
    .X(_04361_));
 sky130_fd_sc_hd__mux2_1 _09374_ (.A0(_04360_),
    .A1(_04361_),
    .S(net1559),
    .X(_04362_));
 sky130_fd_sc_hd__o21ai_1 _09375_ (.A1(net1790),
    .A2(_04358_),
    .B1(_04359_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand2_1 _09376_ (.A(net1781),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__o211a_1 _09377_ (.A1(net1782),
    .A2(_04362_),
    .B1(_04364_),
    .C1(net1671),
    .X(_04365_));
 sky130_fd_sc_hd__o21a_1 _09378_ (.A1(net1790),
    .A2(_04356_),
    .B1(_04357_),
    .X(_04366_));
 sky130_fd_sc_hd__mux2_1 _09379_ (.A0(\core.registers[12][8] ),
    .A1(\core.registers[13][8] ),
    .S(net1508),
    .X(_04367_));
 sky130_fd_sc_hd__mux2_1 _09380_ (.A0(\core.registers[14][8] ),
    .A1(\core.registers[15][8] ),
    .S(net1508),
    .X(_04368_));
 sky130_fd_sc_hd__mux2_1 _09381_ (.A0(_04367_),
    .A1(_04368_),
    .S(net1560),
    .X(_04369_));
 sky130_fd_sc_hd__mux2_1 _09382_ (.A0(_04366_),
    .A1(_04369_),
    .S(net1673),
    .X(_04370_));
 sky130_fd_sc_hd__a211o_1 _09383_ (.A1(net1785),
    .A2(_04370_),
    .B1(_04365_),
    .C1(net1565),
    .X(_04371_));
 sky130_fd_sc_hd__mux2_1 _09384_ (.A0(\core.registers[18][8] ),
    .A1(\core.registers[19][8] ),
    .S(net1509),
    .X(_04372_));
 sky130_fd_sc_hd__mux2_1 _09385_ (.A0(\core.registers[16][8] ),
    .A1(\core.registers[17][8] ),
    .S(net1509),
    .X(_04373_));
 sky130_fd_sc_hd__mux2_1 _09386_ (.A0(_04372_),
    .A1(_04373_),
    .S(net1536),
    .X(_04374_));
 sky130_fd_sc_hd__o221a_1 _09387_ (.A1(net1656),
    .A2(\core.registers[23][8] ),
    .B1(net1509),
    .B2(\core.registers[22][8] ),
    .C1(net1555),
    .X(_04375_));
 sky130_fd_sc_hd__mux2_1 _09388_ (.A0(\core.registers[20][8] ),
    .A1(\core.registers[21][8] ),
    .S(net1509),
    .X(_04376_));
 sky130_fd_sc_hd__mux2_1 _09389_ (.A0(\core.registers[0][8] ),
    .A1(\core.registers[1][8] ),
    .S(net1515),
    .X(_04377_));
 sky130_fd_sc_hd__mux2_1 _09390_ (.A0(\core.registers[2][8] ),
    .A1(\core.registers[3][8] ),
    .S(net1511),
    .X(_04378_));
 sky130_fd_sc_hd__mux2_1 _09391_ (.A0(_04377_),
    .A1(_04378_),
    .S(net1555),
    .X(_04379_));
 sky130_fd_sc_hd__mux2_1 _09392_ (.A0(\core.registers[4][8] ),
    .A1(\core.registers[5][8] ),
    .S(net1509),
    .X(_04380_));
 sky130_fd_sc_hd__o221a_1 _09393_ (.A1(net1657),
    .A2(\core.registers[7][8] ),
    .B1(net1511),
    .B2(\core.registers[6][8] ),
    .C1(net1560),
    .X(_04381_));
 sky130_fd_sc_hd__a211o_1 _09394_ (.A1(net1537),
    .A2(_04380_),
    .B1(_04381_),
    .C1(net1580),
    .X(_04382_));
 sky130_fd_sc_hd__a211o_1 _09395_ (.A1(net1537),
    .A2(_04376_),
    .B1(_04375_),
    .C1(net1580),
    .X(_04383_));
 sky130_fd_sc_hd__o211a_1 _09396_ (.A1(net1589),
    .A2(_04374_),
    .B1(_04383_),
    .C1(net1599),
    .X(_04384_));
 sky130_fd_sc_hd__o211a_1 _09397_ (.A1(net1589),
    .A2(_04379_),
    .B1(_04382_),
    .C1(net1595),
    .X(_04385_));
 sky130_fd_sc_hd__o31a_4 _09398_ (.A1(net1568),
    .A2(_04384_),
    .A3(_04385_),
    .B1(_04371_),
    .X(_04386_));
 sky130_fd_sc_hd__a22o_4 _09399_ (.A1(net1095),
    .A2(_04322_),
    .B1(_04386_),
    .B2(net1046),
    .X(_04387_));
 sky130_fd_sc_hd__o21ai_4 _09400_ (.A1(net1267),
    .A2(_04387_),
    .B1(_04355_),
    .Y(_04388_));
 sky130_fd_sc_hd__or3_4 _09401_ (.A(_04353_),
    .B(_04354_),
    .C(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__o21ai_4 _09402_ (.A1(_04353_),
    .A2(_04354_),
    .B1(_04388_),
    .Y(_04390_));
 sky130_fd_sc_hd__and2_4 _09403_ (.A(_04389_),
    .B(_04390_),
    .X(_04391_));
 sky130_fd_sc_hd__inv_2 _09404_ (.A(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__nand2_2 _09405_ (.A(_03826_),
    .B(net1266),
    .Y(_04393_));
 sky130_fd_sc_hd__mux4_1 _09406_ (.A0(\core.registers[16][7] ),
    .A1(\core.registers[17][7] ),
    .A2(\core.registers[20][7] ),
    .A3(\core.registers[21][7] ),
    .S0(net1496),
    .S1(net1587),
    .X(_04394_));
 sky130_fd_sc_hd__a22o_1 _09407_ (.A1(net1651),
    .A2(\core.registers[22][7] ),
    .B1(\core.registers[23][7] ),
    .B2(net1496),
    .X(_04395_));
 sky130_fd_sc_hd__a22o_1 _09408_ (.A1(net1651),
    .A2(\core.registers[18][7] ),
    .B1(\core.registers[19][7] ),
    .B2(net1496),
    .X(_04396_));
 sky130_fd_sc_hd__mux2_1 _09409_ (.A0(_04395_),
    .A1(_04396_),
    .S(net1576),
    .X(_04397_));
 sky130_fd_sc_hd__a21o_1 _09410_ (.A1(net1550),
    .A2(_04397_),
    .B1(net1569),
    .X(_04398_));
 sky130_fd_sc_hd__a21oi_1 _09411_ (.A1(net1533),
    .A2(_04394_),
    .B1(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__a22o_1 _09412_ (.A1(net1651),
    .A2(\core.registers[30][7] ),
    .B1(\core.registers[31][7] ),
    .B2(net1496),
    .X(_04400_));
 sky130_fd_sc_hd__a22o_1 _09413_ (.A1(net1651),
    .A2(\core.registers[26][7] ),
    .B1(\core.registers[27][7] ),
    .B2(net1496),
    .X(_04401_));
 sky130_fd_sc_hd__mux2_1 _09414_ (.A0(_04400_),
    .A1(_04401_),
    .S(net1576),
    .X(_04402_));
 sky130_fd_sc_hd__mux4_1 _09415_ (.A0(\core.registers[24][7] ),
    .A1(\core.registers[25][7] ),
    .A2(\core.registers[28][7] ),
    .A3(\core.registers[29][7] ),
    .S0(net1496),
    .S1(net1587),
    .X(_04403_));
 sky130_fd_sc_hd__a21o_1 _09416_ (.A1(net1534),
    .A2(_04403_),
    .B1(net1563),
    .X(_04404_));
 sky130_fd_sc_hd__a21oi_2 _09417_ (.A1(net1550),
    .A2(_04402_),
    .B1(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__mux4_1 _09418_ (.A0(\core.registers[0][7] ),
    .A1(\core.registers[1][7] ),
    .A2(\core.registers[4][7] ),
    .A3(\core.registers[5][7] ),
    .S0(net1497),
    .S1(net1587),
    .X(_04406_));
 sky130_fd_sc_hd__and2_1 _09419_ (.A(net1533),
    .B(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__a22o_1 _09420_ (.A1(net1652),
    .A2(\core.registers[6][7] ),
    .B1(\core.registers[7][7] ),
    .B2(net1497),
    .X(_04408_));
 sky130_fd_sc_hd__a22o_1 _09421_ (.A1(net1651),
    .A2(\core.registers[2][7] ),
    .B1(\core.registers[3][7] ),
    .B2(net1497),
    .X(_04409_));
 sky130_fd_sc_hd__mux2_1 _09422_ (.A0(_04408_),
    .A1(_04409_),
    .S(net1576),
    .X(_04410_));
 sky130_fd_sc_hd__a21o_1 _09423_ (.A1(net1550),
    .A2(_04410_),
    .B1(net1569),
    .X(_04411_));
 sky130_fd_sc_hd__nor2_1 _09424_ (.A(_04407_),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__mux4_1 _09425_ (.A0(\core.registers[8][7] ),
    .A1(\core.registers[9][7] ),
    .A2(\core.registers[12][7] ),
    .A3(\core.registers[13][7] ),
    .S0(net1496),
    .S1(net1588),
    .X(_04413_));
 sky130_fd_sc_hd__nand2_1 _09426_ (.A(net1533),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__a22o_1 _09427_ (.A1(net1651),
    .A2(\core.registers[14][7] ),
    .B1(\core.registers[15][7] ),
    .B2(net1496),
    .X(_04415_));
 sky130_fd_sc_hd__a22o_1 _09428_ (.A1(net1652),
    .A2(\core.registers[10][7] ),
    .B1(\core.registers[11][7] ),
    .B2(net1496),
    .X(_04416_));
 sky130_fd_sc_hd__mux2_1 _09429_ (.A0(_04415_),
    .A1(_04416_),
    .S(net1576),
    .X(_04417_));
 sky130_fd_sc_hd__a21oi_1 _09430_ (.A1(net1550),
    .A2(_04417_),
    .B1(net1563),
    .Y(_04418_));
 sky130_fd_sc_hd__a21o_1 _09431_ (.A1(_04414_),
    .A2(_04418_),
    .B1(net1600),
    .X(_04419_));
 sky130_fd_sc_hd__o32a_4 _09432_ (.A1(net1596),
    .A2(_04399_),
    .A3(_04405_),
    .B1(_04412_),
    .B2(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__a22o_1 _09433_ (.A1(\core.pipe1_csrData[7] ),
    .A2(net1247),
    .B1(_04005_),
    .B2(_04029_),
    .X(_04421_));
 sky130_fd_sc_hd__a21o_2 _09434_ (.A1(\core.pipe1_resultRegister[7] ),
    .A2(_03935_),
    .B1(_04421_),
    .X(_04422_));
 sky130_fd_sc_hd__a2bb2o_2 _09435_ (.A1_N(net1044),
    .A2_N(_04420_),
    .B1(net1140),
    .B2(net1096),
    .X(_04423_));
 sky130_fd_sc_hd__o21a_4 _09436_ (.A1(net1267),
    .A2(_04423_),
    .B1(_04393_),
    .X(_04424_));
 sky130_fd_sc_hd__or2_2 _09437_ (.A(net1143),
    .B(net1140),
    .X(_04425_));
 sky130_fd_sc_hd__or2_1 _09438_ (.A(\core.registers[5][7] ),
    .B(net1362),
    .X(_04426_));
 sky130_fd_sc_hd__o211a_1 _09439_ (.A1(\core.registers[4][7] ),
    .A2(net1399),
    .B1(_04426_),
    .C1(net1453),
    .X(_04427_));
 sky130_fd_sc_hd__mux2_1 _09440_ (.A0(\core.registers[0][7] ),
    .A1(\core.registers[1][7] ),
    .S(net1399),
    .X(_04428_));
 sky130_fd_sc_hd__a211o_1 _09441_ (.A1(net1441),
    .A2(_04428_),
    .B1(_04427_),
    .C1(net1348),
    .X(_04429_));
 sky130_fd_sc_hd__o221a_1 _09442_ (.A1(net1688),
    .A2(\core.registers[7][7] ),
    .B1(net1399),
    .B2(\core.registers[6][7] ),
    .C1(net1453),
    .X(_04430_));
 sky130_fd_sc_hd__o221a_1 _09443_ (.A1(net1688),
    .A2(\core.registers[3][7] ),
    .B1(net1399),
    .B2(\core.registers[2][7] ),
    .C1(net1441),
    .X(_04431_));
 sky130_fd_sc_hd__o31a_1 _09444_ (.A1(net1332),
    .A2(_04430_),
    .A3(_04431_),
    .B1(net1323),
    .X(_04432_));
 sky130_fd_sc_hd__or2_1 _09445_ (.A(\core.registers[16][7] ),
    .B(net1398),
    .X(_04433_));
 sky130_fd_sc_hd__o211a_1 _09446_ (.A1(\core.registers[17][7] ),
    .A2(net1362),
    .B1(_04433_),
    .C1(net1441),
    .X(_04434_));
 sky130_fd_sc_hd__mux2_1 _09447_ (.A0(\core.registers[20][7] ),
    .A1(\core.registers[21][7] ),
    .S(net1396),
    .X(_04435_));
 sky130_fd_sc_hd__a211o_1 _09448_ (.A1(net1453),
    .A2(_04435_),
    .B1(_04434_),
    .C1(net1348),
    .X(_04436_));
 sky130_fd_sc_hd__o221a_1 _09449_ (.A1(net1688),
    .A2(\core.registers[23][7] ),
    .B1(net1398),
    .B2(\core.registers[22][7] ),
    .C1(net1453),
    .X(_04437_));
 sky130_fd_sc_hd__o221a_1 _09450_ (.A1(net1688),
    .A2(\core.registers[19][7] ),
    .B1(net1396),
    .B2(\core.registers[18][7] ),
    .C1(net1441),
    .X(_04438_));
 sky130_fd_sc_hd__o31a_1 _09451_ (.A1(net1332),
    .A2(_04437_),
    .A3(_04438_),
    .B1(net1327),
    .X(_04439_));
 sky130_fd_sc_hd__mux2_1 _09452_ (.A0(\core.registers[12][7] ),
    .A1(\core.registers[13][7] ),
    .S(net1396),
    .X(_04440_));
 sky130_fd_sc_hd__mux2_1 _09453_ (.A0(\core.registers[14][7] ),
    .A1(\core.registers[15][7] ),
    .S(net1396),
    .X(_04441_));
 sky130_fd_sc_hd__mux2_1 _09454_ (.A0(_04440_),
    .A1(_04441_),
    .S(net1348),
    .X(_04442_));
 sky130_fd_sc_hd__mux2_1 _09455_ (.A0(\core.registers[28][7] ),
    .A1(\core.registers[29][7] ),
    .S(net1396),
    .X(_04443_));
 sky130_fd_sc_hd__and3_1 _09456_ (.A(net1773),
    .B(\core.registers[31][7] ),
    .C(net1396),
    .X(_04444_));
 sky130_fd_sc_hd__nor2_8 _09457_ (.A(net1703),
    .B(net1777),
    .Y(_04445_));
 sky130_fd_sc_hd__a31o_1 _09458_ (.A1(net1773),
    .A2(net1688),
    .A3(\core.registers[30][7] ),
    .B1(net1710),
    .X(_04446_));
 sky130_fd_sc_hd__a211o_1 _09459_ (.A1(net1701),
    .A2(_04443_),
    .B1(_04444_),
    .C1(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__o211a_1 _09460_ (.A1(net1756),
    .A2(_04442_),
    .B1(_04447_),
    .C1(net1765),
    .X(_04448_));
 sky130_fd_sc_hd__mux2_1 _09461_ (.A0(\core.registers[8][7] ),
    .A1(\core.registers[9][7] ),
    .S(net1396),
    .X(_04449_));
 sky130_fd_sc_hd__mux2_1 _09462_ (.A0(\core.registers[10][7] ),
    .A1(\core.registers[11][7] ),
    .S(net1396),
    .X(_04450_));
 sky130_fd_sc_hd__mux2_1 _09463_ (.A0(_04449_),
    .A1(_04450_),
    .S(net1348),
    .X(_04451_));
 sky130_fd_sc_hd__mux2_1 _09464_ (.A0(\core.registers[24][7] ),
    .A1(\core.registers[25][7] ),
    .S(net1396),
    .X(_04452_));
 sky130_fd_sc_hd__a22o_1 _09465_ (.A1(net1688),
    .A2(\core.registers[26][7] ),
    .B1(\core.registers[27][7] ),
    .B2(net1396),
    .X(_04453_));
 sky130_fd_sc_hd__mux2_1 _09466_ (.A0(_04452_),
    .A1(_04453_),
    .S(net1773),
    .X(_04454_));
 sky130_fd_sc_hd__mux2_1 _09467_ (.A0(_04451_),
    .A1(_04454_),
    .S(net1756),
    .X(_04455_));
 sky130_fd_sc_hd__a21o_1 _09468_ (.A1(_04429_),
    .A2(_04432_),
    .B1(net1432),
    .X(_04456_));
 sky130_fd_sc_hd__a21o_1 _09469_ (.A1(_04436_),
    .A2(_04439_),
    .B1(_04456_),
    .X(_04457_));
 sky130_fd_sc_hd__a211o_1 _09470_ (.A1(net1707),
    .A2(_04455_),
    .B1(_04448_),
    .C1(net1428),
    .X(_04458_));
 sky130_fd_sc_hd__a21o_4 _09471_ (.A1(_04457_),
    .A2(_04458_),
    .B1(net1149),
    .X(_04459_));
 sky130_fd_sc_hd__a31o_1 _09472_ (.A1(net1240),
    .A2(_04425_),
    .A3(_04459_),
    .B1(net1041),
    .X(_04460_));
 sky130_fd_sc_hd__o211a_2 _09473_ (.A1(\core.pipe0_currentInstruction[27] ),
    .A2(net1042),
    .B1(_04460_),
    .C1(net1261),
    .X(_04461_));
 sky130_fd_sc_hd__and2_4 _09474_ (.A(_04424_),
    .B(_04461_),
    .X(_04462_));
 sky130_fd_sc_hd__nor2_4 _09475_ (.A(_04424_),
    .B(_04461_),
    .Y(_04463_));
 sky130_fd_sc_hd__or2_1 _09476_ (.A(net478),
    .B(net1260),
    .X(_04464_));
 sky130_fd_sc_hd__mux2_8 _09477_ (.A0(net167),
    .A1(net138),
    .S(net1734),
    .X(_04465_));
 sky130_fd_sc_hd__o32a_1 _09478_ (.A1(net1638),
    .A2(net1619),
    .A3(_04465_),
    .B1(net1625),
    .B2(\coreWBInterface.readDataBuffered[6] ),
    .X(_04466_));
 sky130_fd_sc_hd__mux2_4 _09479_ (.A0(net112),
    .A1(net147),
    .S(net1735),
    .X(_04467_));
 sky130_fd_sc_hd__nor2_1 _09480_ (.A(_03989_),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__nand2_1 _09481_ (.A(net1745),
    .B(_04468_),
    .Y(_04469_));
 sky130_fd_sc_hd__o211a_1 _09482_ (.A1(\coreWBInterface.readDataBuffered[14] ),
    .A2(net1626),
    .B1(_04031_),
    .C1(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__nor2_2 _09483_ (.A(_03981_),
    .B(_04017_),
    .Y(_04471_));
 sky130_fd_sc_hd__mux2_8 _09484_ (.A0(net130),
    .A1(net165),
    .S(net1737),
    .X(_04472_));
 sky130_fd_sc_hd__o32a_1 _09485_ (.A1(net1639),
    .A2(net1623),
    .A3(_04472_),
    .B1(net1626),
    .B2(\coreWBInterface.readDataBuffered[30] ),
    .X(_04473_));
 sky130_fd_sc_hd__mux2_8 _09486_ (.A0(net121),
    .A1(net156),
    .S(net1736),
    .X(_04474_));
 sky130_fd_sc_hd__o32a_2 _09487_ (.A1(net1639),
    .A2(net1621),
    .A3(_04474_),
    .B1(net1626),
    .B2(\coreWBInterface.readDataBuffered[22] ),
    .X(_04475_));
 sky130_fd_sc_hd__a32o_1 _09488_ (.A1(net1458),
    .A2(net1243),
    .A3(_04475_),
    .B1(_04473_),
    .B2(_04471_),
    .X(_04476_));
 sky130_fd_sc_hd__or3_2 _09489_ (.A(net1618),
    .B(_04470_),
    .C(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__o211a_1 _09490_ (.A1(net1616),
    .A2(_04466_),
    .B1(_04477_),
    .C1(_04029_),
    .X(_04478_));
 sky130_fd_sc_hd__a221o_2 _09491_ (.A1(\core.pipe1_csrData[6] ),
    .A2(net1247),
    .B1(_03935_),
    .B2(\core.pipe1_resultRegister[6] ),
    .C1(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__mux2_1 _09492_ (.A0(\core.registers[28][6] ),
    .A1(\core.registers[29][6] ),
    .S(net1503),
    .X(_04480_));
 sky130_fd_sc_hd__a221o_1 _09493_ (.A1(net1653),
    .A2(\core.registers[30][6] ),
    .B1(\core.registers[31][6] ),
    .B2(net1503),
    .C1(net1666),
    .X(_04481_));
 sky130_fd_sc_hd__and3_1 _09494_ (.A(net1793),
    .B(\core.registers[25][6] ),
    .C(net1632),
    .X(_04482_));
 sky130_fd_sc_hd__a211o_1 _09495_ (.A1(\core.registers[24][6] ),
    .A2(net1460),
    .B1(_04482_),
    .C1(net1792),
    .X(_04483_));
 sky130_fd_sc_hd__a221o_1 _09496_ (.A1(net1653),
    .A2(\core.registers[26][6] ),
    .B1(\core.registers[27][6] ),
    .B2(net1503),
    .C1(net1665),
    .X(_04484_));
 sky130_fd_sc_hd__mux2_1 _09497_ (.A0(\core.registers[8][6] ),
    .A1(\core.registers[9][6] ),
    .S(net1502),
    .X(_04485_));
 sky130_fd_sc_hd__mux2_1 _09498_ (.A0(\core.registers[10][6] ),
    .A1(\core.registers[11][6] ),
    .S(net1502),
    .X(_04486_));
 sky130_fd_sc_hd__mux2_1 _09499_ (.A0(_04485_),
    .A1(_04486_),
    .S(net1552),
    .X(_04487_));
 sky130_fd_sc_hd__a21o_1 _09500_ (.A1(_04483_),
    .A2(_04484_),
    .B1(net1672),
    .X(_04488_));
 sky130_fd_sc_hd__o211a_1 _09501_ (.A1(net1783),
    .A2(_04487_),
    .B1(_04488_),
    .C1(net1670),
    .X(_04489_));
 sky130_fd_sc_hd__mux2_1 _09502_ (.A0(\core.registers[12][6] ),
    .A1(\core.registers[13][6] ),
    .S(net1500),
    .X(_04490_));
 sky130_fd_sc_hd__mux2_1 _09503_ (.A0(\core.registers[14][6] ),
    .A1(\core.registers[15][6] ),
    .S(net1503),
    .X(_04491_));
 sky130_fd_sc_hd__mux2_1 _09504_ (.A0(_04490_),
    .A1(_04491_),
    .S(net1553),
    .X(_04492_));
 sky130_fd_sc_hd__o21a_1 _09505_ (.A1(net1792),
    .A2(_04480_),
    .B1(_04481_),
    .X(_04493_));
 sky130_fd_sc_hd__mux2_1 _09506_ (.A0(_04492_),
    .A1(_04493_),
    .S(net1782),
    .X(_04494_));
 sky130_fd_sc_hd__a211o_1 _09507_ (.A1(net1786),
    .A2(_04494_),
    .B1(_04489_),
    .C1(net1565),
    .X(_04495_));
 sky130_fd_sc_hd__mux2_1 _09508_ (.A0(\core.registers[18][6] ),
    .A1(\core.registers[19][6] ),
    .S(net1501),
    .X(_04496_));
 sky130_fd_sc_hd__mux2_1 _09509_ (.A0(\core.registers[16][6] ),
    .A1(\core.registers[17][6] ),
    .S(net1501),
    .X(_04497_));
 sky130_fd_sc_hd__mux2_1 _09510_ (.A0(_04496_),
    .A1(_04497_),
    .S(net1534),
    .X(_04498_));
 sky130_fd_sc_hd__o221a_1 _09511_ (.A1(net1653),
    .A2(\core.registers[23][6] ),
    .B1(net1501),
    .B2(\core.registers[22][6] ),
    .C1(net1552),
    .X(_04499_));
 sky130_fd_sc_hd__mux2_1 _09512_ (.A0(\core.registers[20][6] ),
    .A1(\core.registers[21][6] ),
    .S(net1501),
    .X(_04500_));
 sky130_fd_sc_hd__or2_1 _09513_ (.A(\core.registers[0][6] ),
    .B(net1500),
    .X(_04501_));
 sky130_fd_sc_hd__o211a_1 _09514_ (.A1(\core.registers[1][6] ),
    .A2(net1460),
    .B1(_04501_),
    .C1(net1535),
    .X(_04502_));
 sky130_fd_sc_hd__mux2_1 _09515_ (.A0(\core.registers[2][6] ),
    .A1(\core.registers[3][6] ),
    .S(net1500),
    .X(_04503_));
 sky130_fd_sc_hd__a211o_1 _09516_ (.A1(net1552),
    .A2(_04503_),
    .B1(_04502_),
    .C1(net1588),
    .X(_04504_));
 sky130_fd_sc_hd__mux2_1 _09517_ (.A0(\core.registers[4][6] ),
    .A1(\core.registers[5][6] ),
    .S(net1500),
    .X(_04505_));
 sky130_fd_sc_hd__o221a_1 _09518_ (.A1(net1653),
    .A2(\core.registers[7][6] ),
    .B1(net1500),
    .B2(\core.registers[6][6] ),
    .C1(net1552),
    .X(_04506_));
 sky130_fd_sc_hd__a211o_1 _09519_ (.A1(net1535),
    .A2(_04505_),
    .B1(_04506_),
    .C1(net1575),
    .X(_04507_));
 sky130_fd_sc_hd__a211o_1 _09520_ (.A1(net1534),
    .A2(_04500_),
    .B1(_04499_),
    .C1(net1577),
    .X(_04508_));
 sky130_fd_sc_hd__o211a_1 _09521_ (.A1(net1588),
    .A2(_04498_),
    .B1(_04508_),
    .C1(net1600),
    .X(_04509_));
 sky130_fd_sc_hd__a311o_1 _09522_ (.A1(net1594),
    .A2(_04504_),
    .A3(_04507_),
    .B1(_04509_),
    .C1(net1569),
    .X(_04510_));
 sky130_fd_sc_hd__and3_2 _09523_ (.A(net1046),
    .B(_04495_),
    .C(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__a21oi_4 _09524_ (.A1(net1096),
    .A2(net1036),
    .B1(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__a21boi_4 _09525_ (.A1(net1260),
    .A2(_04512_),
    .B1_N(_04464_),
    .Y(_04513_));
 sky130_fd_sc_hd__mux4_1 _09526_ (.A0(\core.registers[16][6] ),
    .A1(\core.registers[17][6] ),
    .A2(\core.registers[20][6] ),
    .A3(\core.registers[21][6] ),
    .S0(net1402),
    .S1(net1453),
    .X(_04514_));
 sky130_fd_sc_hd__o22a_1 _09527_ (.A1(net1686),
    .A2(\core.registers[23][6] ),
    .B1(net1402),
    .B2(\core.registers[22][6] ),
    .X(_04515_));
 sky130_fd_sc_hd__o22a_1 _09528_ (.A1(net1686),
    .A2(\core.registers[19][6] ),
    .B1(net1402),
    .B2(\core.registers[18][6] ),
    .X(_04516_));
 sky130_fd_sc_hd__mux2_1 _09529_ (.A0(_04515_),
    .A1(_04516_),
    .S(net1442),
    .X(_04517_));
 sky130_fd_sc_hd__o21a_1 _09530_ (.A1(net1333),
    .A2(_04517_),
    .B1(net1327),
    .X(_04518_));
 sky130_fd_sc_hd__o21ai_1 _09531_ (.A1(net1349),
    .A2(_04514_),
    .B1(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__o22a_1 _09532_ (.A1(net1686),
    .A2(\core.registers[7][6] ),
    .B1(net1401),
    .B2(\core.registers[6][6] ),
    .X(_04520_));
 sky130_fd_sc_hd__o22a_1 _09533_ (.A1(net1683),
    .A2(\core.registers[3][6] ),
    .B1(net1401),
    .B2(\core.registers[2][6] ),
    .X(_04521_));
 sky130_fd_sc_hd__mux2_1 _09534_ (.A0(_04520_),
    .A1(_04521_),
    .S(net1440),
    .X(_04522_));
 sky130_fd_sc_hd__or2_1 _09535_ (.A(net1333),
    .B(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__mux4_1 _09536_ (.A0(\core.registers[0][6] ),
    .A1(\core.registers[1][6] ),
    .A2(\core.registers[4][6] ),
    .A3(\core.registers[5][6] ),
    .S0(net1401),
    .S1(net1452),
    .X(_04524_));
 sky130_fd_sc_hd__o21a_1 _09537_ (.A1(net1349),
    .A2(_04524_),
    .B1(net1321),
    .X(_04525_));
 sky130_fd_sc_hd__a221o_1 _09538_ (.A1(net1690),
    .A2(\core.registers[26][6] ),
    .B1(\core.registers[27][6] ),
    .B2(net1404),
    .C1(net1703),
    .X(_04526_));
 sky130_fd_sc_hd__mux2_1 _09539_ (.A0(\core.registers[24][6] ),
    .A1(\core.registers[25][6] ),
    .S(net1406),
    .X(_04527_));
 sky130_fd_sc_hd__o21ai_1 _09540_ (.A1(net1775),
    .A2(_04527_),
    .B1(_04526_),
    .Y(_04528_));
 sky130_fd_sc_hd__mux2_1 _09541_ (.A0(\core.registers[8][6] ),
    .A1(\core.registers[9][6] ),
    .S(net1403),
    .X(_04529_));
 sky130_fd_sc_hd__mux2_1 _09542_ (.A0(\core.registers[10][6] ),
    .A1(\core.registers[11][6] ),
    .S(net1403),
    .X(_04530_));
 sky130_fd_sc_hd__mux2_1 _09543_ (.A0(_04529_),
    .A1(_04530_),
    .S(net1349),
    .X(_04531_));
 sky130_fd_sc_hd__nor2_1 _09544_ (.A(net1758),
    .B(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__mux2_1 _09545_ (.A0(\core.registers[28][6] ),
    .A1(\core.registers[29][6] ),
    .S(net1404),
    .X(_04533_));
 sky130_fd_sc_hd__a221o_1 _09546_ (.A1(net1686),
    .A2(\core.registers[30][6] ),
    .B1(\core.registers[31][6] ),
    .B2(net1404),
    .C1(net1702),
    .X(_04534_));
 sky130_fd_sc_hd__o21ai_1 _09547_ (.A1(net1775),
    .A2(_04533_),
    .B1(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__a21oi_1 _09548_ (.A1(_04523_),
    .A2(_04525_),
    .B1(net1431),
    .Y(_04536_));
 sky130_fd_sc_hd__a211o_1 _09549_ (.A1(net1758),
    .A2(_04528_),
    .B1(_04532_),
    .C1(net1767),
    .X(_04537_));
 sky130_fd_sc_hd__mux2_1 _09550_ (.A0(\core.registers[12][6] ),
    .A1(\core.registers[13][6] ),
    .S(net1401),
    .X(_04538_));
 sky130_fd_sc_hd__mux2_1 _09551_ (.A0(\core.registers[14][6] ),
    .A1(\core.registers[15][6] ),
    .S(net1404),
    .X(_04539_));
 sky130_fd_sc_hd__mux2_1 _09552_ (.A0(_04538_),
    .A1(_04539_),
    .S(net1349),
    .X(_04540_));
 sky130_fd_sc_hd__nor2_1 _09553_ (.A(net1758),
    .B(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__a211o_1 _09554_ (.A1(net1758),
    .A2(_04535_),
    .B1(_04541_),
    .C1(net1707),
    .X(_04542_));
 sky130_fd_sc_hd__a32o_2 _09555_ (.A1(net1432),
    .A2(_04537_),
    .A3(_04542_),
    .B1(_04519_),
    .B2(_04536_),
    .X(_04543_));
 sky130_fd_sc_hd__a21oi_4 _09556_ (.A1(net1146),
    .A2(_04543_),
    .B1(_04095_),
    .Y(_04544_));
 sky130_fd_sc_hd__o21ai_4 _09557_ (.A1(net1146),
    .A2(net1036),
    .B1(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__nand2_1 _09558_ (.A(net1042),
    .B(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__o211a_1 _09559_ (.A1(\core.pipe0_currentInstruction[26] ),
    .A2(net1042),
    .B1(_04546_),
    .C1(net1261),
    .X(_04547_));
 sky130_fd_sc_hd__and2_2 _09560_ (.A(_04513_),
    .B(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__or2_2 _09561_ (.A(_04513_),
    .B(_04547_),
    .X(_04549_));
 sky130_fd_sc_hd__or2_1 _09562_ (.A(net477),
    .B(net1260),
    .X(_04550_));
 sky130_fd_sc_hd__mux2_8 _09563_ (.A0(net162),
    .A1(net137),
    .S(net1734),
    .X(_04551_));
 sky130_fd_sc_hd__o32a_1 _09564_ (.A1(net1638),
    .A2(net1619),
    .A3(_04551_),
    .B1(net1625),
    .B2(\coreWBInterface.readDataBuffered[5] ),
    .X(_04552_));
 sky130_fd_sc_hd__mux2_4 _09565_ (.A0(net111),
    .A1(net146),
    .S(net1735),
    .X(_04553_));
 sky130_fd_sc_hd__nor2_1 _09566_ (.A(_03989_),
    .B(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__nand2_1 _09567_ (.A(net1745),
    .B(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__o211a_1 _09568_ (.A1(\coreWBInterface.readDataBuffered[13] ),
    .A2(net1626),
    .B1(_04031_),
    .C1(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__mux2_8 _09569_ (.A0(net128),
    .A1(net164),
    .S(net1737),
    .X(_04557_));
 sky130_fd_sc_hd__o32a_1 _09570_ (.A1(net1639),
    .A2(net1623),
    .A3(_04557_),
    .B1(net1627),
    .B2(\coreWBInterface.readDataBuffered[29] ),
    .X(_04558_));
 sky130_fd_sc_hd__mux2_8 _09571_ (.A0(net120),
    .A1(net155),
    .S(net1736),
    .X(_04559_));
 sky130_fd_sc_hd__o32a_1 _09572_ (.A1(net1639),
    .A2(net1621),
    .A3(_04559_),
    .B1(net1626),
    .B2(\coreWBInterface.readDataBuffered[21] ),
    .X(_04560_));
 sky130_fd_sc_hd__a32o_1 _09573_ (.A1(net1458),
    .A2(net1243),
    .A3(_04560_),
    .B1(_04558_),
    .B2(_04471_),
    .X(_04561_));
 sky130_fd_sc_hd__or3_2 _09574_ (.A(net1618),
    .B(_04556_),
    .C(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__o211a_1 _09575_ (.A1(net1616),
    .A2(_04552_),
    .B1(_04562_),
    .C1(_04029_),
    .X(_04563_));
 sky130_fd_sc_hd__a221o_4 _09576_ (.A1(\core.pipe1_csrData[5] ),
    .A2(net1247),
    .B1(_03935_),
    .B2(\core.pipe1_resultRegister[5] ),
    .C1(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__a221o_1 _09577_ (.A1(net1652),
    .A2(\core.registers[30][5] ),
    .B1(\core.registers[31][5] ),
    .B2(net1491),
    .C1(net1666),
    .X(_04565_));
 sky130_fd_sc_hd__mux2_1 _09578_ (.A0(\core.registers[28][5] ),
    .A1(\core.registers[29][5] ),
    .S(net1491),
    .X(_04566_));
 sky130_fd_sc_hd__o21a_1 _09579_ (.A1(net1791),
    .A2(_04566_),
    .B1(_04565_),
    .X(_04567_));
 sky130_fd_sc_hd__mux2_1 _09580_ (.A0(\core.registers[8][5] ),
    .A1(\core.registers[9][5] ),
    .S(net1491),
    .X(_04568_));
 sky130_fd_sc_hd__mux2_1 _09581_ (.A0(\core.registers[10][5] ),
    .A1(\core.registers[11][5] ),
    .S(net1491),
    .X(_04569_));
 sky130_fd_sc_hd__mux2_1 _09582_ (.A0(\core.registers[24][5] ),
    .A1(\core.registers[25][5] ),
    .S(net1491),
    .X(_04570_));
 sky130_fd_sc_hd__a221o_1 _09583_ (.A1(net1652),
    .A2(\core.registers[26][5] ),
    .B1(\core.registers[27][5] ),
    .B2(net1491),
    .C1(net1666),
    .X(_04571_));
 sky130_fd_sc_hd__mux2_1 _09584_ (.A0(_04568_),
    .A1(_04569_),
    .S(net1551),
    .X(_04572_));
 sky130_fd_sc_hd__or2_1 _09585_ (.A(net1782),
    .B(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__o21a_1 _09586_ (.A1(net1791),
    .A2(_04570_),
    .B1(_04571_),
    .X(_04574_));
 sky130_fd_sc_hd__o211a_1 _09587_ (.A1(net1673),
    .A2(_04574_),
    .B1(_04573_),
    .C1(net1670),
    .X(_04575_));
 sky130_fd_sc_hd__mux2_1 _09588_ (.A0(\core.registers[12][5] ),
    .A1(\core.registers[13][5] ),
    .S(net1491),
    .X(_04576_));
 sky130_fd_sc_hd__mux2_1 _09589_ (.A0(\core.registers[14][5] ),
    .A1(\core.registers[15][5] ),
    .S(net1490),
    .X(_04577_));
 sky130_fd_sc_hd__mux2_1 _09590_ (.A0(_04576_),
    .A1(_04577_),
    .S(net1551),
    .X(_04578_));
 sky130_fd_sc_hd__mux2_1 _09591_ (.A0(_04567_),
    .A1(_04578_),
    .S(net1673),
    .X(_04579_));
 sky130_fd_sc_hd__a211o_1 _09592_ (.A1(net1785),
    .A2(_04579_),
    .B1(_04575_),
    .C1(net1563),
    .X(_04580_));
 sky130_fd_sc_hd__mux2_1 _09593_ (.A0(\core.registers[18][5] ),
    .A1(\core.registers[19][5] ),
    .S(net1491),
    .X(_04581_));
 sky130_fd_sc_hd__mux2_1 _09594_ (.A0(\core.registers[16][5] ),
    .A1(\core.registers[17][5] ),
    .S(net1491),
    .X(_04582_));
 sky130_fd_sc_hd__mux2_1 _09595_ (.A0(_04581_),
    .A1(_04582_),
    .S(net1533),
    .X(_04583_));
 sky130_fd_sc_hd__o221a_1 _09596_ (.A1(net1652),
    .A2(\core.registers[23][5] ),
    .B1(net1492),
    .B2(\core.registers[22][5] ),
    .C1(net1551),
    .X(_04584_));
 sky130_fd_sc_hd__mux2_1 _09597_ (.A0(\core.registers[20][5] ),
    .A1(\core.registers[21][5] ),
    .S(net1494),
    .X(_04585_));
 sky130_fd_sc_hd__or2_1 _09598_ (.A(\core.registers[0][5] ),
    .B(net1492),
    .X(_04586_));
 sky130_fd_sc_hd__o211a_1 _09599_ (.A1(\core.registers[1][5] ),
    .A2(net1460),
    .B1(_04586_),
    .C1(net1533),
    .X(_04587_));
 sky130_fd_sc_hd__mux2_1 _09600_ (.A0(\core.registers[2][5] ),
    .A1(\core.registers[3][5] ),
    .S(net1492),
    .X(_04588_));
 sky130_fd_sc_hd__a211o_1 _09601_ (.A1(net1551),
    .A2(_04588_),
    .B1(_04587_),
    .C1(net1587),
    .X(_04589_));
 sky130_fd_sc_hd__mux2_1 _09602_ (.A0(\core.registers[4][5] ),
    .A1(\core.registers[5][5] ),
    .S(net1492),
    .X(_04590_));
 sky130_fd_sc_hd__o221a_1 _09603_ (.A1(net1652),
    .A2(\core.registers[7][5] ),
    .B1(net1493),
    .B2(\core.registers[6][5] ),
    .C1(net1551),
    .X(_04591_));
 sky130_fd_sc_hd__a211o_1 _09604_ (.A1(net1533),
    .A2(_04590_),
    .B1(_04591_),
    .C1(net1576),
    .X(_04592_));
 sky130_fd_sc_hd__a211o_1 _09605_ (.A1(net1533),
    .A2(_04585_),
    .B1(_04584_),
    .C1(net1576),
    .X(_04593_));
 sky130_fd_sc_hd__o211a_1 _09606_ (.A1(net1587),
    .A2(_04583_),
    .B1(_04593_),
    .C1(net1600),
    .X(_04594_));
 sky130_fd_sc_hd__a311o_1 _09607_ (.A1(net1596),
    .A2(_04589_),
    .A3(_04592_),
    .B1(_04594_),
    .C1(net1569),
    .X(_04595_));
 sky130_fd_sc_hd__nand2_2 _09608_ (.A(_04580_),
    .B(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__o2bb2a_4 _09609_ (.A1_N(net1096),
    .A2_N(_04564_),
    .B1(_04596_),
    .B2(net1044),
    .X(_04597_));
 sky130_fd_sc_hd__a21boi_4 _09610_ (.A1(net1260),
    .A2(_04597_),
    .B1_N(_04550_),
    .Y(_04598_));
 sky130_fd_sc_hd__nor2_1 _09611_ (.A(net1146),
    .B(_04564_),
    .Y(_04599_));
 sky130_fd_sc_hd__mux4_1 _09612_ (.A0(\core.registers[16][5] ),
    .A1(\core.registers[17][5] ),
    .A2(\core.registers[20][5] ),
    .A3(\core.registers[21][5] ),
    .S0(net1392),
    .S1(net1453),
    .X(_04600_));
 sky130_fd_sc_hd__o22a_1 _09613_ (.A1(net1687),
    .A2(\core.registers[23][5] ),
    .B1(net1394),
    .B2(\core.registers[22][5] ),
    .X(_04601_));
 sky130_fd_sc_hd__o22a_1 _09614_ (.A1(net1687),
    .A2(\core.registers[19][5] ),
    .B1(net1392),
    .B2(\core.registers[18][5] ),
    .X(_04602_));
 sky130_fd_sc_hd__mux2_1 _09615_ (.A0(_04601_),
    .A1(_04602_),
    .S(net1441),
    .X(_04603_));
 sky130_fd_sc_hd__o21a_1 _09616_ (.A1(net1332),
    .A2(_04603_),
    .B1(net1327),
    .X(_04604_));
 sky130_fd_sc_hd__o21ai_1 _09617_ (.A1(net1347),
    .A2(_04600_),
    .B1(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__o22a_1 _09618_ (.A1(net1687),
    .A2(\core.registers[7][5] ),
    .B1(net1394),
    .B2(\core.registers[6][5] ),
    .X(_04606_));
 sky130_fd_sc_hd__o22a_1 _09619_ (.A1(net1687),
    .A2(\core.registers[3][5] ),
    .B1(net1393),
    .B2(\core.registers[2][5] ),
    .X(_04607_));
 sky130_fd_sc_hd__mux2_1 _09620_ (.A0(_04606_),
    .A1(_04607_),
    .S(net1439),
    .X(_04608_));
 sky130_fd_sc_hd__or2_1 _09621_ (.A(net1332),
    .B(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__mux4_1 _09622_ (.A0(\core.registers[0][5] ),
    .A1(\core.registers[1][5] ),
    .A2(\core.registers[4][5] ),
    .A3(\core.registers[5][5] ),
    .S0(net1393),
    .S1(net1451),
    .X(_04610_));
 sky130_fd_sc_hd__o21a_1 _09623_ (.A1(net1347),
    .A2(_04610_),
    .B1(net1321),
    .X(_04611_));
 sky130_fd_sc_hd__a221o_1 _09624_ (.A1(net1687),
    .A2(\core.registers[26][5] ),
    .B1(\core.registers[27][5] ),
    .B2(net1392),
    .C1(net1702),
    .X(_04612_));
 sky130_fd_sc_hd__mux2_1 _09625_ (.A0(\core.registers[24][5] ),
    .A1(\core.registers[25][5] ),
    .S(net1392),
    .X(_04613_));
 sky130_fd_sc_hd__o21ai_1 _09626_ (.A1(net1772),
    .A2(_04613_),
    .B1(_04612_),
    .Y(_04614_));
 sky130_fd_sc_hd__mux2_1 _09627_ (.A0(\core.registers[8][5] ),
    .A1(\core.registers[9][5] ),
    .S(net1392),
    .X(_04615_));
 sky130_fd_sc_hd__mux2_1 _09628_ (.A0(\core.registers[10][5] ),
    .A1(\core.registers[11][5] ),
    .S(net1392),
    .X(_04616_));
 sky130_fd_sc_hd__mux2_1 _09629_ (.A0(_04615_),
    .A1(_04616_),
    .S(net1347),
    .X(_04617_));
 sky130_fd_sc_hd__nor2_1 _09630_ (.A(net1756),
    .B(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__a221o_1 _09631_ (.A1(net1687),
    .A2(\core.registers[30][5] ),
    .B1(\core.registers[31][5] ),
    .B2(net1392),
    .C1(net1702),
    .X(_04619_));
 sky130_fd_sc_hd__mux2_1 _09632_ (.A0(\core.registers[28][5] ),
    .A1(\core.registers[29][5] ),
    .S(net1395),
    .X(_04620_));
 sky130_fd_sc_hd__o21ai_1 _09633_ (.A1(net1772),
    .A2(_04620_),
    .B1(_04619_),
    .Y(_04621_));
 sky130_fd_sc_hd__a21oi_1 _09634_ (.A1(_04609_),
    .A2(_04611_),
    .B1(net1432),
    .Y(_04622_));
 sky130_fd_sc_hd__a211o_1 _09635_ (.A1(net1756),
    .A2(_04614_),
    .B1(_04618_),
    .C1(net1765),
    .X(_04623_));
 sky130_fd_sc_hd__mux2_1 _09636_ (.A0(\core.registers[12][5] ),
    .A1(\core.registers[13][5] ),
    .S(net1392),
    .X(_04624_));
 sky130_fd_sc_hd__mux2_1 _09637_ (.A0(\core.registers[14][5] ),
    .A1(\core.registers[15][5] ),
    .S(net1391),
    .X(_04625_));
 sky130_fd_sc_hd__mux2_1 _09638_ (.A0(_04624_),
    .A1(_04625_),
    .S(net1347),
    .X(_04626_));
 sky130_fd_sc_hd__nor2_1 _09639_ (.A(net1756),
    .B(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__a211o_1 _09640_ (.A1(net1756),
    .A2(_04621_),
    .B1(_04627_),
    .C1(net1707),
    .X(_04628_));
 sky130_fd_sc_hd__a32o_4 _09641_ (.A1(net1432),
    .A2(_04623_),
    .A3(_04628_),
    .B1(_04605_),
    .B2(_04622_),
    .X(_04629_));
 sky130_fd_sc_hd__a211o_4 _09642_ (.A1(net1146),
    .A2(_04629_),
    .B1(_04599_),
    .C1(_04095_),
    .X(_04630_));
 sky130_fd_sc_hd__nand2_1 _09643_ (.A(net1042),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__o211a_4 _09644_ (.A1(\core.pipe0_currentInstruction[25] ),
    .A2(net1042),
    .B1(_04631_),
    .C1(net1261),
    .X(_04632_));
 sky130_fd_sc_hd__and2_2 _09645_ (.A(_04598_),
    .B(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__nor2_1 _09646_ (.A(_04598_),
    .B(_04632_),
    .Y(_04634_));
 sky130_fd_sc_hd__xor2_4 _09647_ (.A(_04598_),
    .B(_04632_),
    .X(_04635_));
 sky130_fd_sc_hd__or2_1 _09648_ (.A(_04633_),
    .B(_04634_),
    .X(_04636_));
 sky130_fd_sc_hd__mux2_8 _09649_ (.A0(net151),
    .A1(net136),
    .S(net1734),
    .X(_04637_));
 sky130_fd_sc_hd__o32a_1 _09650_ (.A1(net1640),
    .A2(net1620),
    .A3(_04637_),
    .B1(net1628),
    .B2(\coreWBInterface.readDataBuffered[4] ),
    .X(_04638_));
 sky130_fd_sc_hd__mux2_4 _09651_ (.A0(net110),
    .A1(net145),
    .S(net1735),
    .X(_04639_));
 sky130_fd_sc_hd__nor2_1 _09652_ (.A(_03989_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__nand2_1 _09653_ (.A(net1745),
    .B(_04640_),
    .Y(_04641_));
 sky130_fd_sc_hd__o211a_1 _09654_ (.A1(\coreWBInterface.readDataBuffered[12] ),
    .A2(net1626),
    .B1(_04031_),
    .C1(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__mux2_8 _09655_ (.A0(net127),
    .A1(net163),
    .S(net1737),
    .X(_04643_));
 sky130_fd_sc_hd__o32a_1 _09656_ (.A1(net1640),
    .A2(net1623),
    .A3(_04643_),
    .B1(net1626),
    .B2(\coreWBInterface.readDataBuffered[28] ),
    .X(_04644_));
 sky130_fd_sc_hd__mux2_8 _09657_ (.A0(net119),
    .A1(net154),
    .S(net1736),
    .X(_04645_));
 sky130_fd_sc_hd__o32a_1 _09658_ (.A1(net1639),
    .A2(net1621),
    .A3(_04645_),
    .B1(net1627),
    .B2(\coreWBInterface.readDataBuffered[20] ),
    .X(_04646_));
 sky130_fd_sc_hd__a32o_1 _09659_ (.A1(net1458),
    .A2(net1243),
    .A3(_04646_),
    .B1(_04644_),
    .B2(_04471_),
    .X(_04647_));
 sky130_fd_sc_hd__or3_2 _09660_ (.A(net1617),
    .B(_04642_),
    .C(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__o211a_1 _09661_ (.A1(net1616),
    .A2(_04638_),
    .B1(_04648_),
    .C1(_04029_),
    .X(_04649_));
 sky130_fd_sc_hd__a221o_4 _09662_ (.A1(\core.pipe1_csrData[4] ),
    .A2(net1247),
    .B1(_03935_),
    .B2(\core.pipe1_resultRegister[4] ),
    .C1(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__mux2_1 _09663_ (.A0(\core.registers[24][4] ),
    .A1(\core.registers[25][4] ),
    .S(net1399),
    .X(_04651_));
 sky130_fd_sc_hd__a221o_1 _09664_ (.A1(net1689),
    .A2(\core.registers[26][4] ),
    .B1(\core.registers[27][4] ),
    .B2(net1399),
    .C1(net1701),
    .X(_04652_));
 sky130_fd_sc_hd__o21ai_1 _09665_ (.A1(net1774),
    .A2(_04651_),
    .B1(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__mux2_1 _09666_ (.A0(\core.registers[10][4] ),
    .A1(\core.registers[11][4] ),
    .S(net1399),
    .X(_04654_));
 sky130_fd_sc_hd__mux2_1 _09667_ (.A0(\core.registers[8][4] ),
    .A1(\core.registers[9][4] ),
    .S(net1399),
    .X(_04655_));
 sky130_fd_sc_hd__mux2_1 _09668_ (.A0(_04654_),
    .A1(_04655_),
    .S(net1332),
    .X(_04656_));
 sky130_fd_sc_hd__nor2_1 _09669_ (.A(net1757),
    .B(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__a211o_1 _09670_ (.A1(net1756),
    .A2(_04653_),
    .B1(_04657_),
    .C1(net1765),
    .X(_04658_));
 sky130_fd_sc_hd__mux2_1 _09671_ (.A0(\core.registers[28][4] ),
    .A1(\core.registers[29][4] ),
    .S(net1399),
    .X(_04659_));
 sky130_fd_sc_hd__a221o_1 _09672_ (.A1(net1686),
    .A2(\core.registers[30][4] ),
    .B1(\core.registers[31][4] ),
    .B2(net1394),
    .C1(net1702),
    .X(_04660_));
 sky130_fd_sc_hd__o21ai_1 _09673_ (.A1(net1772),
    .A2(_04659_),
    .B1(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__mux4_1 _09674_ (.A0(\core.registers[16][4] ),
    .A1(\core.registers[17][4] ),
    .A2(\core.registers[20][4] ),
    .A3(\core.registers[21][4] ),
    .S0(net1394),
    .S1(net1453),
    .X(_04662_));
 sky130_fd_sc_hd__o22a_1 _09675_ (.A1(net1686),
    .A2(\core.registers[23][4] ),
    .B1(net1394),
    .B2(\core.registers[22][4] ),
    .X(_04663_));
 sky130_fd_sc_hd__o22a_1 _09676_ (.A1(net1686),
    .A2(\core.registers[19][4] ),
    .B1(net1402),
    .B2(\core.registers[18][4] ),
    .X(_04664_));
 sky130_fd_sc_hd__mux2_1 _09677_ (.A0(_04663_),
    .A1(_04664_),
    .S(net1441),
    .X(_04665_));
 sky130_fd_sc_hd__o21a_1 _09678_ (.A1(net1332),
    .A2(_04665_),
    .B1(net1327),
    .X(_04666_));
 sky130_fd_sc_hd__o21ai_1 _09679_ (.A1(net1347),
    .A2(_04662_),
    .B1(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__o22a_1 _09680_ (.A1(net1690),
    .A2(\core.registers[7][4] ),
    .B1(net1402),
    .B2(\core.registers[6][4] ),
    .X(_04668_));
 sky130_fd_sc_hd__o22a_1 _09681_ (.A1(net1687),
    .A2(\core.registers[3][4] ),
    .B1(net1404),
    .B2(\core.registers[2][4] ),
    .X(_04669_));
 sky130_fd_sc_hd__mux2_1 _09682_ (.A0(_04668_),
    .A1(_04669_),
    .S(net1441),
    .X(_04670_));
 sky130_fd_sc_hd__or2_1 _09683_ (.A(net1333),
    .B(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__mux4_1 _09684_ (.A0(\core.registers[0][4] ),
    .A1(\core.registers[1][4] ),
    .A2(\core.registers[4][4] ),
    .A3(\core.registers[5][4] ),
    .S0(net1401),
    .S1(net1457),
    .X(_04672_));
 sky130_fd_sc_hd__o21a_1 _09685_ (.A1(net1349),
    .A2(_04672_),
    .B1(net1323),
    .X(_04673_));
 sky130_fd_sc_hd__a21oi_1 _09686_ (.A1(_04671_),
    .A2(_04673_),
    .B1(net1433),
    .Y(_04674_));
 sky130_fd_sc_hd__mux2_1 _09687_ (.A0(\core.registers[12][4] ),
    .A1(\core.registers[13][4] ),
    .S(net1394),
    .X(_04675_));
 sky130_fd_sc_hd__mux2_1 _09688_ (.A0(\core.registers[14][4] ),
    .A1(\core.registers[15][4] ),
    .S(net1394),
    .X(_04676_));
 sky130_fd_sc_hd__mux2_1 _09689_ (.A0(_04675_),
    .A1(_04676_),
    .S(net1347),
    .X(_04677_));
 sky130_fd_sc_hd__nor2_1 _09690_ (.A(net1756),
    .B(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hd__a211o_1 _09691_ (.A1(net1756),
    .A2(_04661_),
    .B1(_04678_),
    .C1(net1707),
    .X(_04679_));
 sky130_fd_sc_hd__a32o_2 _09692_ (.A1(net1432),
    .A2(_04658_),
    .A3(_04679_),
    .B1(_04674_),
    .B2(_04667_),
    .X(_04680_));
 sky130_fd_sc_hd__a21oi_2 _09693_ (.A1(net1146),
    .A2(_04680_),
    .B1(_04095_),
    .Y(_04681_));
 sky130_fd_sc_hd__o21ai_4 _09694_ (.A1(net1146),
    .A2(_04650_),
    .B1(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__nor2_1 _09695_ (.A(\core.pipe0_currentInstruction[11] ),
    .B(net1154),
    .Y(_04683_));
 sky130_fd_sc_hd__a211o_2 _09696_ (.A1(net1154),
    .A2(_04682_),
    .B1(_04683_),
    .C1(net1093),
    .X(_04684_));
 sky130_fd_sc_hd__nand2_2 _09697_ (.A(net1755),
    .B(_04069_),
    .Y(_04685_));
 sky130_fd_sc_hd__a21oi_4 _09698_ (.A1(_04684_),
    .A2(_04685_),
    .B1(net1265),
    .Y(_04686_));
 sky130_fd_sc_hd__a21o_2 _09699_ (.A1(_04684_),
    .A2(_04685_),
    .B1(net1265),
    .X(_04687_));
 sky130_fd_sc_hd__mux2_1 _09700_ (.A0(\core.registers[24][4] ),
    .A1(\core.registers[25][4] ),
    .S(net1497),
    .X(_04688_));
 sky130_fd_sc_hd__a221o_1 _09701_ (.A1(net1655),
    .A2(\core.registers[26][4] ),
    .B1(\core.registers[27][4] ),
    .B2(net1497),
    .C1(net1664),
    .X(_04689_));
 sky130_fd_sc_hd__mux2_1 _09702_ (.A0(\core.registers[8][4] ),
    .A1(\core.registers[9][4] ),
    .S(net1497),
    .X(_04690_));
 sky130_fd_sc_hd__mux2_1 _09703_ (.A0(\core.registers[10][4] ),
    .A1(\core.registers[11][4] ),
    .S(net1497),
    .X(_04691_));
 sky130_fd_sc_hd__mux2_1 _09704_ (.A0(\core.registers[28][4] ),
    .A1(\core.registers[29][4] ),
    .S(net1497),
    .X(_04692_));
 sky130_fd_sc_hd__a221o_1 _09705_ (.A1(net1652),
    .A2(\core.registers[30][4] ),
    .B1(\core.registers[31][4] ),
    .B2(net1493),
    .C1(net1666),
    .X(_04693_));
 sky130_fd_sc_hd__mux2_1 _09706_ (.A0(_04690_),
    .A1(_04691_),
    .S(net1550),
    .X(_04694_));
 sky130_fd_sc_hd__o21ai_1 _09707_ (.A1(net1790),
    .A2(_04688_),
    .B1(_04689_),
    .Y(_04695_));
 sky130_fd_sc_hd__nand2_1 _09708_ (.A(net1781),
    .B(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__o211a_1 _09709_ (.A1(net1781),
    .A2(_04694_),
    .B1(_04696_),
    .C1(net1671),
    .X(_04697_));
 sky130_fd_sc_hd__o21a_1 _09710_ (.A1(net1791),
    .A2(_04692_),
    .B1(_04693_),
    .X(_04698_));
 sky130_fd_sc_hd__mux2_1 _09711_ (.A0(\core.registers[12][4] ),
    .A1(\core.registers[13][4] ),
    .S(net1493),
    .X(_04699_));
 sky130_fd_sc_hd__mux2_1 _09712_ (.A0(\core.registers[14][4] ),
    .A1(\core.registers[15][4] ),
    .S(net1493),
    .X(_04700_));
 sky130_fd_sc_hd__mux2_1 _09713_ (.A0(_04699_),
    .A1(_04700_),
    .S(net1551),
    .X(_04701_));
 sky130_fd_sc_hd__mux2_1 _09714_ (.A0(_04698_),
    .A1(_04701_),
    .S(net1673),
    .X(_04702_));
 sky130_fd_sc_hd__a211o_1 _09715_ (.A1(net1785),
    .A2(_04702_),
    .B1(_04697_),
    .C1(net1563),
    .X(_04703_));
 sky130_fd_sc_hd__mux2_1 _09716_ (.A0(\core.registers[18][4] ),
    .A1(\core.registers[19][4] ),
    .S(net1501),
    .X(_04704_));
 sky130_fd_sc_hd__mux2_1 _09717_ (.A0(\core.registers[16][4] ),
    .A1(\core.registers[17][4] ),
    .S(net1492),
    .X(_04705_));
 sky130_fd_sc_hd__mux2_1 _09718_ (.A0(_04704_),
    .A1(_04705_),
    .S(net1533),
    .X(_04706_));
 sky130_fd_sc_hd__o221a_1 _09719_ (.A1(net1653),
    .A2(\core.registers[23][4] ),
    .B1(net1493),
    .B2(\core.registers[22][4] ),
    .C1(net1552),
    .X(_04707_));
 sky130_fd_sc_hd__mux2_1 _09720_ (.A0(\core.registers[20][4] ),
    .A1(\core.registers[21][4] ),
    .S(net1493),
    .X(_04708_));
 sky130_fd_sc_hd__mux2_1 _09721_ (.A0(\core.registers[0][4] ),
    .A1(\core.registers[1][4] ),
    .S(net1501),
    .X(_04709_));
 sky130_fd_sc_hd__mux2_1 _09722_ (.A0(\core.registers[2][4] ),
    .A1(\core.registers[3][4] ),
    .S(net1503),
    .X(_04710_));
 sky130_fd_sc_hd__mux2_1 _09723_ (.A0(_04709_),
    .A1(_04710_),
    .S(net1552),
    .X(_04711_));
 sky130_fd_sc_hd__mux2_1 _09724_ (.A0(\core.registers[4][4] ),
    .A1(\core.registers[5][4] ),
    .S(net1501),
    .X(_04712_));
 sky130_fd_sc_hd__o221a_1 _09725_ (.A1(net1653),
    .A2(\core.registers[7][4] ),
    .B1(net1501),
    .B2(\core.registers[6][4] ),
    .C1(net1552),
    .X(_04713_));
 sky130_fd_sc_hd__a211o_1 _09726_ (.A1(net1535),
    .A2(_04712_),
    .B1(_04713_),
    .C1(net1577),
    .X(_04714_));
 sky130_fd_sc_hd__a211o_1 _09727_ (.A1(net1533),
    .A2(_04708_),
    .B1(_04707_),
    .C1(net1576),
    .X(_04715_));
 sky130_fd_sc_hd__o211a_1 _09728_ (.A1(net1587),
    .A2(_04706_),
    .B1(_04715_),
    .C1(net1600),
    .X(_04716_));
 sky130_fd_sc_hd__o211a_1 _09729_ (.A1(net1588),
    .A2(_04711_),
    .B1(_04714_),
    .C1(net1596),
    .X(_04717_));
 sky130_fd_sc_hd__o31a_2 _09730_ (.A1(net1569),
    .A2(_04716_),
    .A3(_04717_),
    .B1(_04703_),
    .X(_04718_));
 sky130_fd_sc_hd__a22o_4 _09731_ (.A1(net1095),
    .A2(_04650_),
    .B1(_04718_),
    .B2(net1046),
    .X(_04719_));
 sky130_fd_sc_hd__mux2_8 _09732_ (.A0(net1748),
    .A1(_04719_),
    .S(net1260),
    .X(_04720_));
 sky130_fd_sc_hd__nand2_4 _09733_ (.A(_04686_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__inv_2 _09734_ (.A(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__or2_4 _09735_ (.A(_04686_),
    .B(_04720_),
    .X(_04723_));
 sky130_fd_sc_hd__nand2_4 _09736_ (.A(_04721_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__a32o_1 _09737_ (.A1(_03982_),
    .A2(net1458),
    .A3(_04024_),
    .B1(_04471_),
    .B2(_03977_),
    .X(_04725_));
 sky130_fd_sc_hd__mux2_8 _09738_ (.A0(net140),
    .A1(net135),
    .S(net1734),
    .X(_04726_));
 sky130_fd_sc_hd__o32a_1 _09739_ (.A1(net1638),
    .A2(net1620),
    .A3(_04726_),
    .B1(net1625),
    .B2(\coreWBInterface.readDataBuffered[3] ),
    .X(_04727_));
 sky130_fd_sc_hd__o21a_1 _09740_ (.A1(net1616),
    .A2(_04727_),
    .B1(_04029_),
    .X(_04728_));
 sky130_fd_sc_hd__o31a_1 _09741_ (.A1(net1617),
    .A2(_04035_),
    .A3(_04725_),
    .B1(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__a221o_4 _09742_ (.A1(\core.pipe1_csrData[3] ),
    .A2(net1247),
    .B1(_03935_),
    .B2(\core.pipe1_resultRegister[3] ),
    .C1(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__nor2_1 _09743_ (.A(net1143),
    .B(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__mux2_1 _09744_ (.A0(\core.registers[24][3] ),
    .A1(\core.registers[25][3] ),
    .S(net1377),
    .X(_04732_));
 sky130_fd_sc_hd__a221o_1 _09745_ (.A1(net1680),
    .A2(\core.registers[26][3] ),
    .B1(\core.registers[27][3] ),
    .B2(net1377),
    .C1(net1700),
    .X(_04733_));
 sky130_fd_sc_hd__o21a_1 _09746_ (.A1(net1770),
    .A2(_04732_),
    .B1(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__mux2_1 _09747_ (.A0(\core.registers[10][3] ),
    .A1(\core.registers[11][3] ),
    .S(net1377),
    .X(_04735_));
 sky130_fd_sc_hd__mux2_1 _09748_ (.A0(\core.registers[8][3] ),
    .A1(\core.registers[9][3] ),
    .S(net1377),
    .X(_04736_));
 sky130_fd_sc_hd__mux2_1 _09749_ (.A0(_04735_),
    .A1(_04736_),
    .S(net1330),
    .X(_04737_));
 sky130_fd_sc_hd__mux2_1 _09750_ (.A0(_04734_),
    .A1(_04737_),
    .S(net1709),
    .X(_04738_));
 sky130_fd_sc_hd__or2_1 _09751_ (.A(\core.registers[28][3] ),
    .B(net1377),
    .X(_04739_));
 sky130_fd_sc_hd__o211a_1 _09752_ (.A1(\core.registers[29][3] ),
    .A2(net1359),
    .B1(_04739_),
    .C1(net1700),
    .X(_04740_));
 sky130_fd_sc_hd__a31o_1 _09753_ (.A1(net1770),
    .A2(net1680),
    .A3(\core.registers[30][3] ),
    .B1(net1709),
    .X(_04741_));
 sky130_fd_sc_hd__a31o_1 _09754_ (.A1(net1770),
    .A2(\core.registers[31][3] ),
    .A3(net1377),
    .B1(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__mux4_1 _09755_ (.A0(\core.registers[16][3] ),
    .A1(\core.registers[17][3] ),
    .A2(\core.registers[20][3] ),
    .A3(\core.registers[21][3] ),
    .S0(net1381),
    .S1(net1448),
    .X(_04743_));
 sky130_fd_sc_hd__o22a_1 _09756_ (.A1(net1680),
    .A2(\core.registers[23][3] ),
    .B1(net1377),
    .B2(\core.registers[22][3] ),
    .X(_04744_));
 sky130_fd_sc_hd__o22a_1 _09757_ (.A1(net1680),
    .A2(\core.registers[19][3] ),
    .B1(net1381),
    .B2(\core.registers[18][3] ),
    .X(_04745_));
 sky130_fd_sc_hd__mux2_1 _09758_ (.A0(_04744_),
    .A1(_04745_),
    .S(net1435),
    .X(_04746_));
 sky130_fd_sc_hd__o21a_1 _09759_ (.A1(net1330),
    .A2(_04746_),
    .B1(net1324),
    .X(_04747_));
 sky130_fd_sc_hd__o21ai_1 _09760_ (.A1(net1344),
    .A2(_04743_),
    .B1(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__o22a_1 _09761_ (.A1(net1680),
    .A2(\core.registers[7][3] ),
    .B1(net1377),
    .B2(\core.registers[6][3] ),
    .X(_04749_));
 sky130_fd_sc_hd__o22a_1 _09762_ (.A1(net1680),
    .A2(\core.registers[3][3] ),
    .B1(net1380),
    .B2(\core.registers[2][3] ),
    .X(_04750_));
 sky130_fd_sc_hd__mux2_1 _09763_ (.A0(_04749_),
    .A1(_04750_),
    .S(net1435),
    .X(_04751_));
 sky130_fd_sc_hd__or2_1 _09764_ (.A(net1330),
    .B(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__mux4_1 _09765_ (.A0(\core.registers[0][3] ),
    .A1(\core.registers[1][3] ),
    .A2(\core.registers[4][3] ),
    .A3(\core.registers[5][3] ),
    .S0(net1384),
    .S1(net1450),
    .X(_04753_));
 sky130_fd_sc_hd__o21a_1 _09766_ (.A1(net1344),
    .A2(_04753_),
    .B1(net1320),
    .X(_04754_));
 sky130_fd_sc_hd__a21oi_1 _09767_ (.A1(_04752_),
    .A2(_04754_),
    .B1(net1429),
    .Y(_04755_));
 sky130_fd_sc_hd__nand2_1 _09768_ (.A(_04748_),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__mux2_1 _09769_ (.A0(\core.registers[12][3] ),
    .A1(\core.registers[13][3] ),
    .S(net1377),
    .X(_04757_));
 sky130_fd_sc_hd__mux2_1 _09770_ (.A0(\core.registers[14][3] ),
    .A1(\core.registers[15][3] ),
    .S(net1377),
    .X(_04758_));
 sky130_fd_sc_hd__mux2_1 _09771_ (.A0(_04757_),
    .A1(_04758_),
    .S(net1344),
    .X(_04759_));
 sky130_fd_sc_hd__o221a_1 _09772_ (.A1(_04740_),
    .A2(_04742_),
    .B1(_04759_),
    .B2(net1755),
    .C1(net1763),
    .X(_04760_));
 sky130_fd_sc_hd__a211o_2 _09773_ (.A1(net1705),
    .A2(_04738_),
    .B1(_04760_),
    .C1(net1427),
    .X(_04761_));
 sky130_fd_sc_hd__a21oi_4 _09774_ (.A1(_04756_),
    .A2(_04761_),
    .B1(net1148),
    .Y(_04762_));
 sky130_fd_sc_hd__o31a_1 _09775_ (.A1(_04095_),
    .A2(_04731_),
    .A3(_04762_),
    .B1(net1154),
    .X(_04763_));
 sky130_fd_sc_hd__a211o_2 _09776_ (.A1(_03844_),
    .A2(_04057_),
    .B1(net1093),
    .C1(_04763_),
    .X(_04764_));
 sky130_fd_sc_hd__nand2_2 _09777_ (.A(net1762),
    .B(net1093),
    .Y(_04765_));
 sky130_fd_sc_hd__a21oi_4 _09778_ (.A1(_04764_),
    .A2(_04765_),
    .B1(net1265),
    .Y(_04766_));
 sky130_fd_sc_hd__a21o_1 _09779_ (.A1(_04764_),
    .A2(_04765_),
    .B1(net1265),
    .X(_04767_));
 sky130_fd_sc_hd__or2_1 _09780_ (.A(net475),
    .B(net1260),
    .X(_04768_));
 sky130_fd_sc_hd__a221o_1 _09781_ (.A1(net1647),
    .A2(\core.registers[30][3] ),
    .B1(\core.registers[31][3] ),
    .B2(net1476),
    .C1(net1667),
    .X(_04769_));
 sky130_fd_sc_hd__mux2_1 _09782_ (.A0(\core.registers[28][3] ),
    .A1(\core.registers[29][3] ),
    .S(net1476),
    .X(_04770_));
 sky130_fd_sc_hd__o21a_1 _09783_ (.A1(net1788),
    .A2(_04770_),
    .B1(_04769_),
    .X(_04771_));
 sky130_fd_sc_hd__mux2_1 _09784_ (.A0(\core.registers[8][3] ),
    .A1(\core.registers[9][3] ),
    .S(net1476),
    .X(_04772_));
 sky130_fd_sc_hd__mux2_1 _09785_ (.A0(\core.registers[10][3] ),
    .A1(\core.registers[11][3] ),
    .S(net1476),
    .X(_04773_));
 sky130_fd_sc_hd__mux2_1 _09786_ (.A0(\core.registers[24][3] ),
    .A1(\core.registers[25][3] ),
    .S(net1476),
    .X(_04774_));
 sky130_fd_sc_hd__a221o_1 _09787_ (.A1(net1647),
    .A2(\core.registers[26][3] ),
    .B1(\core.registers[27][3] ),
    .B2(net1476),
    .C1(net1663),
    .X(_04775_));
 sky130_fd_sc_hd__mux2_1 _09788_ (.A0(_04772_),
    .A1(_04773_),
    .S(net1546),
    .X(_04776_));
 sky130_fd_sc_hd__nor2_1 _09789_ (.A(net1779),
    .B(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__o21ai_1 _09790_ (.A1(net1788),
    .A2(_04774_),
    .B1(_04775_),
    .Y(_04778_));
 sky130_fd_sc_hd__a211o_1 _09791_ (.A1(net1779),
    .A2(_04778_),
    .B1(_04777_),
    .C1(net1784),
    .X(_04779_));
 sky130_fd_sc_hd__mux2_1 _09792_ (.A0(\core.registers[12][3] ),
    .A1(\core.registers[13][3] ),
    .S(net1476),
    .X(_04780_));
 sky130_fd_sc_hd__mux2_1 _09793_ (.A0(\core.registers[14][3] ),
    .A1(\core.registers[15][3] ),
    .S(net1476),
    .X(_04781_));
 sky130_fd_sc_hd__mux2_1 _09794_ (.A0(_04780_),
    .A1(_04781_),
    .S(net1546),
    .X(_04782_));
 sky130_fd_sc_hd__mux2_1 _09795_ (.A0(_04771_),
    .A1(_04782_),
    .S(net1674),
    .X(_04783_));
 sky130_fd_sc_hd__a21oi_1 _09796_ (.A1(net1784),
    .A2(_04783_),
    .B1(net1562),
    .Y(_04784_));
 sky130_fd_sc_hd__mux2_1 _09797_ (.A0(\core.registers[18][3] ),
    .A1(\core.registers[19][3] ),
    .S(net1476),
    .X(_04785_));
 sky130_fd_sc_hd__mux2_1 _09798_ (.A0(\core.registers[16][3] ),
    .A1(\core.registers[17][3] ),
    .S(net1480),
    .X(_04786_));
 sky130_fd_sc_hd__mux2_1 _09799_ (.A0(_04785_),
    .A1(_04786_),
    .S(net1530),
    .X(_04787_));
 sky130_fd_sc_hd__o221a_1 _09800_ (.A1(net1647),
    .A2(\core.registers[23][3] ),
    .B1(net1476),
    .B2(\core.registers[22][3] ),
    .C1(net1546),
    .X(_04788_));
 sky130_fd_sc_hd__mux2_1 _09801_ (.A0(\core.registers[20][3] ),
    .A1(\core.registers[21][3] ),
    .S(net1480),
    .X(_04789_));
 sky130_fd_sc_hd__or2_1 _09802_ (.A(\core.registers[0][3] ),
    .B(net1483),
    .X(_04790_));
 sky130_fd_sc_hd__o211a_1 _09803_ (.A1(\core.registers[1][3] ),
    .A2(net1459),
    .B1(_04790_),
    .C1(net1530),
    .X(_04791_));
 sky130_fd_sc_hd__mux2_1 _09804_ (.A0(\core.registers[2][3] ),
    .A1(\core.registers[3][3] ),
    .S(net1479),
    .X(_04792_));
 sky130_fd_sc_hd__a211o_1 _09805_ (.A1(net1548),
    .A2(_04792_),
    .B1(_04791_),
    .C1(net1585),
    .X(_04793_));
 sky130_fd_sc_hd__mux2_1 _09806_ (.A0(\core.registers[4][3] ),
    .A1(\core.registers[5][3] ),
    .S(net1483),
    .X(_04794_));
 sky130_fd_sc_hd__o221a_1 _09807_ (.A1(net1647),
    .A2(\core.registers[7][3] ),
    .B1(net1481),
    .B2(\core.registers[6][3] ),
    .C1(net1546),
    .X(_04795_));
 sky130_fd_sc_hd__a211o_1 _09808_ (.A1(net1530),
    .A2(_04794_),
    .B1(_04795_),
    .C1(net1574),
    .X(_04796_));
 sky130_fd_sc_hd__a211o_1 _09809_ (.A1(net1530),
    .A2(_04789_),
    .B1(_04788_),
    .C1(net1574),
    .X(_04797_));
 sky130_fd_sc_hd__o211a_1 _09810_ (.A1(net1585),
    .A2(_04787_),
    .B1(_04797_),
    .C1(net1597),
    .X(_04798_));
 sky130_fd_sc_hd__a31o_1 _09811_ (.A1(net1594),
    .A2(_04793_),
    .A3(_04796_),
    .B1(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__a2bb2o_4 _09812_ (.A1_N(net1567),
    .A2_N(_04799_),
    .B1(_04784_),
    .B2(_04779_),
    .X(_04800_));
 sky130_fd_sc_hd__o2bb2a_2 _09813_ (.A1_N(net1096),
    .A2_N(_04730_),
    .B1(_04800_),
    .B2(net1044),
    .X(_04801_));
 sky130_fd_sc_hd__a21boi_4 _09814_ (.A1(net1260),
    .A2(_04801_),
    .B1_N(_04768_),
    .Y(_04802_));
 sky130_fd_sc_hd__clkinv_2 _09815_ (.A(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__nor2_4 _09816_ (.A(_04766_),
    .B(_04802_),
    .Y(_04804_));
 sky130_fd_sc_hd__nand2_2 _09817_ (.A(net748),
    .B(_04803_),
    .Y(_04805_));
 sky130_fd_sc_hd__nor2_4 _09818_ (.A(net748),
    .B(_04803_),
    .Y(_04806_));
 sky130_fd_sc_hd__and3_1 _09819_ (.A(_03982_),
    .B(_04016_),
    .C(_04135_),
    .X(_04807_));
 sky130_fd_sc_hd__a31o_1 _09820_ (.A1(_03982_),
    .A2(net1458),
    .A3(_04138_),
    .B1(net1617),
    .X(_04808_));
 sky130_fd_sc_hd__or3b_2 _09821_ (.A(_04808_),
    .B(_04807_),
    .C_N(_04144_),
    .X(_04809_));
 sky130_fd_sc_hd__mux2_8 _09822_ (.A0(net129),
    .A1(net134),
    .S(net1734),
    .X(_04810_));
 sky130_fd_sc_hd__o32a_1 _09823_ (.A1(net1638),
    .A2(net1619),
    .A3(_04810_),
    .B1(net1625),
    .B2(\coreWBInterface.readDataBuffered[2] ),
    .X(_04811_));
 sky130_fd_sc_hd__o211a_1 _09824_ (.A1(net1616),
    .A2(_04811_),
    .B1(_04809_),
    .C1(_04029_),
    .X(_04812_));
 sky130_fd_sc_hd__a221o_4 _09825_ (.A1(\core.pipe1_csrData[2] ),
    .A2(net1247),
    .B1(_03935_),
    .B2(\core.pipe1_resultRegister[2] ),
    .C1(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__or2_1 _09826_ (.A(\core.registers[13][2] ),
    .B(net1359),
    .X(_04814_));
 sky130_fd_sc_hd__o211a_1 _09827_ (.A1(\core.registers[12][2] ),
    .A2(net1387),
    .B1(net1340),
    .C1(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__a22o_1 _09828_ (.A1(net1681),
    .A2(\core.registers[14][2] ),
    .B1(\core.registers[15][2] ),
    .B2(net1387),
    .X(_04816_));
 sky130_fd_sc_hd__and2_1 _09829_ (.A(net1346),
    .B(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__or2_1 _09830_ (.A(\core.registers[9][2] ),
    .B(net1359),
    .X(_04818_));
 sky130_fd_sc_hd__o211a_1 _09831_ (.A1(\core.registers[8][2] ),
    .A2(net1387),
    .B1(net1331),
    .C1(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__a22o_1 _09832_ (.A1(net1683),
    .A2(\core.registers[10][2] ),
    .B1(\core.registers[11][2] ),
    .B2(net1387),
    .X(_04820_));
 sky130_fd_sc_hd__a21o_1 _09833_ (.A1(net1346),
    .A2(_04820_),
    .B1(net1764),
    .X(_04821_));
 sky130_fd_sc_hd__o32a_1 _09834_ (.A1(net1705),
    .A2(_04815_),
    .A3(_04817_),
    .B1(_04819_),
    .B2(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__mux2_1 _09835_ (.A0(\core.registers[28][2] ),
    .A1(\core.registers[29][2] ),
    .S(net1388),
    .X(_04823_));
 sky130_fd_sc_hd__a22o_1 _09836_ (.A1(net1683),
    .A2(\core.registers[30][2] ),
    .B1(\core.registers[31][2] ),
    .B2(net1388),
    .X(_04824_));
 sky130_fd_sc_hd__mux2_1 _09837_ (.A0(\core.registers[24][2] ),
    .A1(\core.registers[25][2] ),
    .S(net1388),
    .X(_04825_));
 sky130_fd_sc_hd__a22o_1 _09838_ (.A1(net1683),
    .A2(\core.registers[26][2] ),
    .B1(\core.registers[27][2] ),
    .B2(net1388),
    .X(_04826_));
 sky130_fd_sc_hd__mux4_1 _09839_ (.A0(_04823_),
    .A1(_04824_),
    .A2(_04825_),
    .A3(_04826_),
    .S0(net1772),
    .S1(net1705),
    .X(_04827_));
 sky130_fd_sc_hd__o21a_1 _09840_ (.A1(net1709),
    .A2(_04827_),
    .B1(net1431),
    .X(_04828_));
 sky130_fd_sc_hd__o21ai_2 _09841_ (.A1(net1755),
    .A2(_04822_),
    .B1(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__mux2_1 _09842_ (.A0(\core.registers[0][2] ),
    .A1(\core.registers[1][2] ),
    .S(net1401),
    .X(_04830_));
 sky130_fd_sc_hd__mux2_1 _09843_ (.A0(\core.registers[4][2] ),
    .A1(\core.registers[5][2] ),
    .S(net1390),
    .X(_04831_));
 sky130_fd_sc_hd__mux2_1 _09844_ (.A0(\core.registers[2][2] ),
    .A1(\core.registers[3][2] ),
    .S(net1388),
    .X(_04832_));
 sky130_fd_sc_hd__mux2_1 _09845_ (.A0(_04830_),
    .A1(_04832_),
    .S(net1349),
    .X(_04833_));
 sky130_fd_sc_hd__or3_1 _09846_ (.A(net1684),
    .B(\core.registers[7][2] ),
    .C(net1633),
    .X(_04834_));
 sky130_fd_sc_hd__o211a_1 _09847_ (.A1(\core.registers[6][2] ),
    .A2(net1387),
    .B1(net1346),
    .C1(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__a211o_1 _09848_ (.A1(net1331),
    .A2(_04831_),
    .B1(_04835_),
    .C1(net1440),
    .X(_04836_));
 sky130_fd_sc_hd__o211a_1 _09849_ (.A1(net1452),
    .A2(_04833_),
    .B1(_04836_),
    .C1(net1321),
    .X(_04837_));
 sky130_fd_sc_hd__mux2_1 _09850_ (.A0(\core.registers[16][2] ),
    .A1(\core.registers[17][2] ),
    .S(net1387),
    .X(_04838_));
 sky130_fd_sc_hd__mux2_1 _09851_ (.A0(\core.registers[20][2] ),
    .A1(\core.registers[21][2] ),
    .S(net1387),
    .X(_04839_));
 sky130_fd_sc_hd__mux2_1 _09852_ (.A0(\core.registers[18][2] ),
    .A1(\core.registers[19][2] ),
    .S(net1388),
    .X(_04840_));
 sky130_fd_sc_hd__mux2_1 _09853_ (.A0(_04838_),
    .A1(_04840_),
    .S(net1346),
    .X(_04841_));
 sky130_fd_sc_hd__or3_1 _09854_ (.A(net1684),
    .B(\core.registers[23][2] ),
    .C(net1634),
    .X(_04842_));
 sky130_fd_sc_hd__o211a_1 _09855_ (.A1(\core.registers[22][2] ),
    .A2(net1387),
    .B1(net1346),
    .C1(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__a211o_1 _09856_ (.A1(net1331),
    .A2(_04839_),
    .B1(_04843_),
    .C1(net1440),
    .X(_04844_));
 sky130_fd_sc_hd__o211a_1 _09857_ (.A1(net1452),
    .A2(_04841_),
    .B1(_04844_),
    .C1(net1325),
    .X(_04845_));
 sky130_fd_sc_hd__o21ai_2 _09858_ (.A1(_04837_),
    .A2(_04845_),
    .B1(net1428),
    .Y(_04846_));
 sky130_fd_sc_hd__nand3_4 _09859_ (.A(net1143),
    .B(_04829_),
    .C(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__o211ai_4 _09860_ (.A1(net1143),
    .A2(net1087),
    .B1(_04847_),
    .C1(net1239),
    .Y(_04848_));
 sky130_fd_sc_hd__nor2_1 _09861_ (.A(\core.pipe0_currentInstruction[9] ),
    .B(net1154),
    .Y(_04849_));
 sky130_fd_sc_hd__a211o_4 _09862_ (.A1(net1154),
    .A2(_04848_),
    .B1(_04849_),
    .C1(net1093),
    .X(_04850_));
 sky130_fd_sc_hd__nand2_2 _09863_ (.A(net1764),
    .B(net1093),
    .Y(_04851_));
 sky130_fd_sc_hd__a21oi_4 _09864_ (.A1(_04850_),
    .A2(_04851_),
    .B1(net1263),
    .Y(_04852_));
 sky130_fd_sc_hd__a21o_4 _09865_ (.A1(_04850_),
    .A2(_04851_),
    .B1(net1263),
    .X(_04853_));
 sky130_fd_sc_hd__nand2_1 _09866_ (.A(_03827_),
    .B(net1267),
    .Y(_04854_));
 sky130_fd_sc_hd__mux4_1 _09867_ (.A0(\core.registers[24][2] ),
    .A1(\core.registers[25][2] ),
    .A2(\core.registers[28][2] ),
    .A3(\core.registers[29][2] ),
    .S0(net1488),
    .S1(\core.pipe0_currentInstruction[17] ),
    .X(_04855_));
 sky130_fd_sc_hd__a221o_1 _09868_ (.A1(net1650),
    .A2(\core.registers[30][2] ),
    .B1(\core.registers[31][2] ),
    .B2(net1488),
    .C1(net1670),
    .X(_04856_));
 sky130_fd_sc_hd__a221o_1 _09869_ (.A1(net1650),
    .A2(\core.registers[26][2] ),
    .B1(\core.registers[27][2] ),
    .B2(net1488),
    .C1(net1785),
    .X(_04857_));
 sky130_fd_sc_hd__a31o_1 _09870_ (.A1(net1791),
    .A2(_04856_),
    .A3(_04857_),
    .B1(net1674),
    .X(_04858_));
 sky130_fd_sc_hd__a21oi_1 _09871_ (.A1(net1666),
    .A2(_04855_),
    .B1(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__mux4_1 _09872_ (.A0(\core.registers[8][2] ),
    .A1(\core.registers[9][2] ),
    .A2(\core.registers[12][2] ),
    .A3(\core.registers[13][2] ),
    .S0(net1487),
    .S1(net1784),
    .X(_04860_));
 sky130_fd_sc_hd__a221o_1 _09873_ (.A1(net1662),
    .A2(\core.registers[14][2] ),
    .B1(\core.registers[15][2] ),
    .B2(net1487),
    .C1(net1669),
    .X(_04861_));
 sky130_fd_sc_hd__a221o_1 _09874_ (.A1(net1650),
    .A2(\core.registers[10][2] ),
    .B1(\core.registers[11][2] ),
    .B2(net1487),
    .C1(net1784),
    .X(_04862_));
 sky130_fd_sc_hd__a31o_1 _09875_ (.A1(net1788),
    .A2(_04861_),
    .A3(_04862_),
    .B1(net1779),
    .X(_04863_));
 sky130_fd_sc_hd__a21oi_1 _09876_ (.A1(net1667),
    .A2(_04860_),
    .B1(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__nor2_1 _09877_ (.A(_04859_),
    .B(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__mux2_1 _09878_ (.A0(\core.registers[18][2] ),
    .A1(\core.registers[19][2] ),
    .S(net1488),
    .X(_04866_));
 sky130_fd_sc_hd__mux2_1 _09879_ (.A0(\core.registers[16][2] ),
    .A1(\core.registers[17][2] ),
    .S(net1487),
    .X(_04867_));
 sky130_fd_sc_hd__mux2_1 _09880_ (.A0(_04866_),
    .A1(_04867_),
    .S(net1532),
    .X(_04868_));
 sky130_fd_sc_hd__o221a_1 _09881_ (.A1(net1650),
    .A2(\core.registers[23][2] ),
    .B1(net1487),
    .B2(\core.registers[22][2] ),
    .C1(net1549),
    .X(_04869_));
 sky130_fd_sc_hd__mux2_1 _09882_ (.A0(\core.registers[20][2] ),
    .A1(\core.registers[21][2] ),
    .S(net1487),
    .X(_04870_));
 sky130_fd_sc_hd__or2_1 _09883_ (.A(\core.registers[0][2] ),
    .B(net1500),
    .X(_04871_));
 sky130_fd_sc_hd__o211a_1 _09884_ (.A1(\core.registers[1][2] ),
    .A2(net1459),
    .B1(_04871_),
    .C1(net1532),
    .X(_04872_));
 sky130_fd_sc_hd__mux2_1 _09885_ (.A0(\core.registers[2][2] ),
    .A1(\core.registers[3][2] ),
    .S(net1488),
    .X(_04873_));
 sky130_fd_sc_hd__a211o_1 _09886_ (.A1(net1549),
    .A2(_04873_),
    .B1(_04872_),
    .C1(net1586),
    .X(_04874_));
 sky130_fd_sc_hd__mux2_1 _09887_ (.A0(\core.registers[4][2] ),
    .A1(\core.registers[5][2] ),
    .S(net1489),
    .X(_04875_));
 sky130_fd_sc_hd__o221a_1 _09888_ (.A1(net1650),
    .A2(\core.registers[7][2] ),
    .B1(net1487),
    .B2(\core.registers[6][2] ),
    .C1(net1549),
    .X(_04876_));
 sky130_fd_sc_hd__a211o_1 _09889_ (.A1(net1532),
    .A2(_04875_),
    .B1(_04876_),
    .C1(net1575),
    .X(_04877_));
 sky130_fd_sc_hd__a211o_1 _09890_ (.A1(net1532),
    .A2(_04870_),
    .B1(_04869_),
    .C1(net1575),
    .X(_04878_));
 sky130_fd_sc_hd__o211a_1 _09891_ (.A1(net1586),
    .A2(_04868_),
    .B1(_04878_),
    .C1(net1598),
    .X(_04879_));
 sky130_fd_sc_hd__a311o_1 _09892_ (.A1(net1593),
    .A2(_04874_),
    .A3(_04877_),
    .B1(_04879_),
    .C1(net1567),
    .X(_04880_));
 sky130_fd_sc_hd__o21ai_2 _09893_ (.A1(net1562),
    .A2(_04865_),
    .B1(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__o2bb2a_2 _09894_ (.A1_N(net1096),
    .A2_N(net1087),
    .B1(_04881_),
    .B2(net1044),
    .X(_04882_));
 sky130_fd_sc_hd__a21bo_4 _09895_ (.A1(net1261),
    .A2(_04882_),
    .B1_N(_04854_),
    .X(_04883_));
 sky130_fd_sc_hd__inv_2 _09896_ (.A(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__nor2_1 _09897_ (.A(_04853_),
    .B(_04883_),
    .Y(_04885_));
 sky130_fd_sc_hd__nand2_2 _09898_ (.A(_04853_),
    .B(_04883_),
    .Y(_04886_));
 sky130_fd_sc_hd__a32o_4 _09899_ (.A1(_03898_),
    .A2(_03924_),
    .A3(_03926_),
    .B1(_04027_),
    .B2(_04028_),
    .X(_04887_));
 sky130_fd_sc_hd__a21oi_2 _09900_ (.A1(\core.pipe1_csrData[1] ),
    .A2(net1250),
    .B1(net1237),
    .Y(_04888_));
 sky130_fd_sc_hd__or3b_1 _09901_ (.A(_04225_),
    .B(_03981_),
    .C_N(_03988_),
    .X(_04889_));
 sky130_fd_sc_hd__or3_1 _09902_ (.A(_03981_),
    .B(_04017_),
    .C(_04221_),
    .X(_04890_));
 sky130_fd_sc_hd__and4_1 _09903_ (.A(_04029_),
    .B(_04233_),
    .C(_04889_),
    .D(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__a21oi_1 _09904_ (.A1(net1749),
    .A2(_04891_),
    .B1(_04888_),
    .Y(_04892_));
 sky130_fd_sc_hd__a31o_1 _09905_ (.A1(_04233_),
    .A2(_04889_),
    .A3(_04890_),
    .B1(_03830_),
    .X(_04893_));
 sky130_fd_sc_hd__mux2_8 _09906_ (.A0(net118),
    .A1(net133),
    .S(net1734),
    .X(_04894_));
 sky130_fd_sc_hd__nor2_1 _09907_ (.A(net1620),
    .B(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__o32a_1 _09908_ (.A1(net1639),
    .A2(net1620),
    .A3(_04894_),
    .B1(net1627),
    .B2(\coreWBInterface.readDataBuffered[1] ),
    .X(_04896_));
 sky130_fd_sc_hd__a21oi_1 _09909_ (.A1(_03830_),
    .A2(_04896_),
    .B1(_04030_),
    .Y(_04897_));
 sky130_fd_sc_hd__a21oi_1 _09910_ (.A1(_04893_),
    .A2(_04897_),
    .B1(_03935_),
    .Y(_04898_));
 sky130_fd_sc_hd__o22a_1 _09911_ (.A1(net1244),
    .A2(_04892_),
    .B1(_04898_),
    .B2(\core.pipe1_resultRegister[1] ),
    .X(_04899_));
 sky130_fd_sc_hd__mux2_1 _09912_ (.A0(\core.registers[16][1] ),
    .A1(\core.registers[17][1] ),
    .S(net1417),
    .X(_04900_));
 sky130_fd_sc_hd__o221a_1 _09913_ (.A1(net1777),
    .A2(\core.registers[20][1] ),
    .B1(\core.registers[21][1] ),
    .B2(net1362),
    .C1(net1457),
    .X(_04901_));
 sky130_fd_sc_hd__a211o_1 _09914_ (.A1(net1442),
    .A2(_04900_),
    .B1(_04901_),
    .C1(net1354),
    .X(_04902_));
 sky130_fd_sc_hd__o221a_1 _09915_ (.A1(net1695),
    .A2(\core.registers[19][1] ),
    .B1(net1417),
    .B2(\core.registers[18][1] ),
    .C1(net1442),
    .X(_04903_));
 sky130_fd_sc_hd__o221a_1 _09916_ (.A1(net1689),
    .A2(\core.registers[23][1] ),
    .B1(net1404),
    .B2(\core.registers[22][1] ),
    .C1(net1457),
    .X(_04904_));
 sky130_fd_sc_hd__mux2_1 _09917_ (.A0(\core.registers[0][1] ),
    .A1(\core.registers[1][1] ),
    .S(net1404),
    .X(_04905_));
 sky130_fd_sc_hd__o221a_1 _09918_ (.A1(net1777),
    .A2(\core.registers[4][1] ),
    .B1(\core.registers[5][1] ),
    .B2(net1362),
    .C1(net1457),
    .X(_04906_));
 sky130_fd_sc_hd__a211o_1 _09919_ (.A1(net1442),
    .A2(_04905_),
    .B1(_04906_),
    .C1(net1355),
    .X(_04907_));
 sky130_fd_sc_hd__o221a_1 _09920_ (.A1(net1689),
    .A2(\core.registers[3][1] ),
    .B1(net1405),
    .B2(\core.registers[2][1] ),
    .C1(net1442),
    .X(_04908_));
 sky130_fd_sc_hd__o221a_1 _09921_ (.A1(net1689),
    .A2(\core.registers[7][1] ),
    .B1(net1404),
    .B2(\core.registers[6][1] ),
    .C1(net1453),
    .X(_04909_));
 sky130_fd_sc_hd__o311a_1 _09922_ (.A1(net1333),
    .A2(_04908_),
    .A3(_04909_),
    .B1(net1323),
    .C1(_04907_),
    .X(_04910_));
 sky130_fd_sc_hd__o311a_1 _09923_ (.A1(net1333),
    .A2(_04903_),
    .A3(_04904_),
    .B1(net1327),
    .C1(_04902_),
    .X(_04911_));
 sky130_fd_sc_hd__o21a_1 _09924_ (.A1(_04910_),
    .A2(_04911_),
    .B1(_04077_),
    .X(_04912_));
 sky130_fd_sc_hd__mux2_1 _09925_ (.A0(\core.registers[8][1] ),
    .A1(\core.registers[9][1] ),
    .S(net1404),
    .X(_04913_));
 sky130_fd_sc_hd__a221o_1 _09926_ (.A1(net1689),
    .A2(\core.registers[10][1] ),
    .B1(\core.registers[11][1] ),
    .B2(net1399),
    .C1(net1332),
    .X(_04914_));
 sky130_fd_sc_hd__o21a_1 _09927_ (.A1(net1349),
    .A2(_04913_),
    .B1(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__a31o_1 _09928_ (.A1(net1777),
    .A2(\core.registers[25][1] ),
    .A3(net1631),
    .B1(net1774),
    .X(_04916_));
 sky130_fd_sc_hd__a21o_1 _09929_ (.A1(\core.registers[24][1] ),
    .A2(net1362),
    .B1(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__a221o_1 _09930_ (.A1(net1689),
    .A2(\core.registers[26][1] ),
    .B1(\core.registers[27][1] ),
    .B2(net1405),
    .C1(net1701),
    .X(_04918_));
 sky130_fd_sc_hd__a21o_1 _09931_ (.A1(_04917_),
    .A2(_04918_),
    .B1(net1765),
    .X(_04919_));
 sky130_fd_sc_hd__mux2_1 _09932_ (.A0(\core.registers[30][1] ),
    .A1(\core.registers[31][1] ),
    .S(net1405),
    .X(_04920_));
 sky130_fd_sc_hd__mux2_1 _09933_ (.A0(\core.registers[28][1] ),
    .A1(\core.registers[29][1] ),
    .S(net1405),
    .X(_04921_));
 sky130_fd_sc_hd__mux2_1 _09934_ (.A0(_04920_),
    .A1(_04921_),
    .S(net1334),
    .X(_04922_));
 sky130_fd_sc_hd__or2_1 _09935_ (.A(net1442),
    .B(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__mux2_1 _09936_ (.A0(\core.registers[14][1] ),
    .A1(\core.registers[15][1] ),
    .S(net1400),
    .X(_04924_));
 sky130_fd_sc_hd__mux2_1 _09937_ (.A0(\core.registers[12][1] ),
    .A1(\core.registers[13][1] ),
    .S(net1400),
    .X(_04925_));
 sky130_fd_sc_hd__mux2_1 _09938_ (.A0(_04924_),
    .A1(_04925_),
    .S(net1334),
    .X(_04926_));
 sky130_fd_sc_hd__o221a_1 _09939_ (.A1(net1765),
    .A2(_04915_),
    .B1(_04926_),
    .B2(net1441),
    .C1(net1323),
    .X(_04927_));
 sky130_fd_sc_hd__a31o_1 _09940_ (.A1(net1327),
    .A2(_04919_),
    .A3(_04923_),
    .B1(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__a211o_2 _09941_ (.A1(net1432),
    .A2(_04928_),
    .B1(_04912_),
    .C1(net1149),
    .X(_04929_));
 sky130_fd_sc_hd__o211ai_4 _09942_ (.A1(net1147),
    .A2(net1084),
    .B1(_04929_),
    .C1(net1241),
    .Y(_04930_));
 sky130_fd_sc_hd__nor2_1 _09943_ (.A(\core.pipe0_currentInstruction[8] ),
    .B(net1154),
    .Y(_04931_));
 sky130_fd_sc_hd__a211o_1 _09944_ (.A1(net1154),
    .A2(_04930_),
    .B1(_04931_),
    .C1(_04069_),
    .X(_04932_));
 sky130_fd_sc_hd__nand2_1 _09945_ (.A(net1771),
    .B(net1093),
    .Y(_04933_));
 sky130_fd_sc_hd__a21o_1 _09946_ (.A1(_04932_),
    .A2(_04933_),
    .B1(net1265),
    .X(_04934_));
 sky130_fd_sc_hd__inv_2 _09947_ (.A(net886),
    .Y(_04935_));
 sky130_fd_sc_hd__or2_1 _09948_ (.A(net461),
    .B(net1260),
    .X(_04936_));
 sky130_fd_sc_hd__mux2_1 _09949_ (.A0(\core.registers[28][1] ),
    .A1(\core.registers[29][1] ),
    .S(net1504),
    .X(_04937_));
 sky130_fd_sc_hd__a221o_1 _09950_ (.A1(net1654),
    .A2(\core.registers[30][1] ),
    .B1(\core.registers[31][1] ),
    .B2(net1504),
    .C1(net1665),
    .X(_04938_));
 sky130_fd_sc_hd__mux2_1 _09951_ (.A0(\core.registers[8][1] ),
    .A1(\core.registers[9][1] ),
    .S(net1503),
    .X(_04939_));
 sky130_fd_sc_hd__mux2_1 _09952_ (.A0(\core.registers[10][1] ),
    .A1(\core.registers[11][1] ),
    .S(net1503),
    .X(_04940_));
 sky130_fd_sc_hd__mux2_1 _09953_ (.A0(_04939_),
    .A1(_04940_),
    .S(net1553),
    .X(_04941_));
 sky130_fd_sc_hd__or2_1 _09954_ (.A(\core.registers[25][1] ),
    .B(net1460),
    .X(_04942_));
 sky130_fd_sc_hd__o21a_1 _09955_ (.A1(\core.registers[24][1] ),
    .A2(net1503),
    .B1(net1665),
    .X(_04943_));
 sky130_fd_sc_hd__a22o_1 _09956_ (.A1(net1653),
    .A2(\core.registers[26][1] ),
    .B1(\core.registers[27][1] ),
    .B2(net1504),
    .X(_04944_));
 sky130_fd_sc_hd__a221o_1 _09957_ (.A1(_04942_),
    .A2(_04943_),
    .B1(_04944_),
    .B2(net1791),
    .C1(net1672),
    .X(_04945_));
 sky130_fd_sc_hd__o211a_1 _09958_ (.A1(net1781),
    .A2(_04941_),
    .B1(_04945_),
    .C1(net1671),
    .X(_04946_));
 sky130_fd_sc_hd__o21a_1 _09959_ (.A1(net1792),
    .A2(_04937_),
    .B1(_04938_),
    .X(_04947_));
 sky130_fd_sc_hd__mux2_1 _09960_ (.A0(\core.registers[12][1] ),
    .A1(\core.registers[13][1] ),
    .S(net1498),
    .X(_04948_));
 sky130_fd_sc_hd__mux2_1 _09961_ (.A0(\core.registers[14][1] ),
    .A1(\core.registers[15][1] ),
    .S(net1498),
    .X(_04949_));
 sky130_fd_sc_hd__mux2_1 _09962_ (.A0(_04948_),
    .A1(_04949_),
    .S(net1550),
    .X(_04950_));
 sky130_fd_sc_hd__mux2_1 _09963_ (.A0(_04947_),
    .A1(_04950_),
    .S(net1673),
    .X(_04951_));
 sky130_fd_sc_hd__a21o_1 _09964_ (.A1(net1785),
    .A2(_04951_),
    .B1(net1563),
    .X(_04952_));
 sky130_fd_sc_hd__mux2_1 _09965_ (.A0(\core.registers[18][1] ),
    .A1(\core.registers[19][1] ),
    .S(net1515),
    .X(_04953_));
 sky130_fd_sc_hd__mux2_1 _09966_ (.A0(\core.registers[16][1] ),
    .A1(\core.registers[17][1] ),
    .S(net1515),
    .X(_04954_));
 sky130_fd_sc_hd__mux2_1 _09967_ (.A0(_04953_),
    .A1(_04954_),
    .S(net1540),
    .X(_04955_));
 sky130_fd_sc_hd__o221a_1 _09968_ (.A1(net1653),
    .A2(\core.registers[23][1] ),
    .B1(net1504),
    .B2(\core.registers[22][1] ),
    .C1(net1553),
    .X(_04956_));
 sky130_fd_sc_hd__mux2_1 _09969_ (.A0(\core.registers[20][1] ),
    .A1(\core.registers[21][1] ),
    .S(net1504),
    .X(_04957_));
 sky130_fd_sc_hd__mux2_1 _09970_ (.A0(\core.registers[0][1] ),
    .A1(\core.registers[1][1] ),
    .S(net1504),
    .X(_04958_));
 sky130_fd_sc_hd__mux2_1 _09971_ (.A0(\core.registers[2][1] ),
    .A1(\core.registers[3][1] ),
    .S(net1504),
    .X(_04959_));
 sky130_fd_sc_hd__mux2_1 _09972_ (.A0(_04958_),
    .A1(_04959_),
    .S(net1553),
    .X(_04960_));
 sky130_fd_sc_hd__mux2_1 _09973_ (.A0(\core.registers[4][1] ),
    .A1(\core.registers[5][1] ),
    .S(net1504),
    .X(_04961_));
 sky130_fd_sc_hd__o221a_1 _09974_ (.A1(net1654),
    .A2(\core.registers[7][1] ),
    .B1(net1503),
    .B2(\core.registers[6][1] ),
    .C1(net1553),
    .X(_04962_));
 sky130_fd_sc_hd__a211o_1 _09975_ (.A1(net1534),
    .A2(_04961_),
    .B1(_04962_),
    .C1(net1577),
    .X(_04963_));
 sky130_fd_sc_hd__a211o_1 _09976_ (.A1(net1535),
    .A2(_04957_),
    .B1(_04956_),
    .C1(net1577),
    .X(_04964_));
 sky130_fd_sc_hd__o211a_1 _09977_ (.A1(net1588),
    .A2(_04955_),
    .B1(_04964_),
    .C1(net1600),
    .X(_04965_));
 sky130_fd_sc_hd__o211a_1 _09978_ (.A1(net1588),
    .A2(_04960_),
    .B1(_04963_),
    .C1(net1596),
    .X(_04966_));
 sky130_fd_sc_hd__o32a_4 _09979_ (.A1(net1569),
    .A2(_04965_),
    .A3(_04966_),
    .B1(_04946_),
    .B2(_04952_),
    .X(_04967_));
 sky130_fd_sc_hd__a22oi_4 _09980_ (.A1(net1095),
    .A2(net1084),
    .B1(_04967_),
    .B2(net1046),
    .Y(_04968_));
 sky130_fd_sc_hd__a21boi_4 _09981_ (.A1(net1260),
    .A2(_04968_),
    .B1_N(_04936_),
    .Y(_04969_));
 sky130_fd_sc_hd__and2b_2 _09982_ (.A_N(net889),
    .B(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__xnor2_4 _09983_ (.A(net889),
    .B(_04969_),
    .Y(_04971_));
 sky130_fd_sc_hd__xor2_4 _09984_ (.A(net889),
    .B(_04969_),
    .X(_04972_));
 sky130_fd_sc_hd__a21oi_2 _09985_ (.A1(\core.pipe1_csrData[0] ),
    .A2(net1249),
    .B1(net1238),
    .Y(_04973_));
 sky130_fd_sc_hd__and3_1 _09986_ (.A(_03982_),
    .B(_04016_),
    .C(_04309_),
    .X(_04974_));
 sky130_fd_sc_hd__nor2_1 _09987_ (.A(net1242),
    .B(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hd__a31oi_2 _09988_ (.A1(net1750),
    .A2(_04319_),
    .A3(_04975_),
    .B1(_04973_),
    .Y(_04976_));
 sky130_fd_sc_hd__o21a_1 _09989_ (.A1(_04313_),
    .A2(_04974_),
    .B1(net1749),
    .X(_04977_));
 sky130_fd_sc_hd__mux2_4 _09990_ (.A0(net107),
    .A1(net132),
    .S(net1734),
    .X(_04978_));
 sky130_fd_sc_hd__nor2_1 _09991_ (.A(net1619),
    .B(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__nand2_1 _09992_ (.A(net1745),
    .B(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__o211a_1 _09993_ (.A1(\coreWBInterface.readDataBuffered[0] ),
    .A2(net1625),
    .B1(_04980_),
    .C1(net1712),
    .X(_04981_));
 sky130_fd_sc_hd__o31a_1 _09994_ (.A1(net1242),
    .A2(_04977_),
    .A3(_04981_),
    .B1(net1188),
    .X(_04982_));
 sky130_fd_sc_hd__o22a_4 _09995_ (.A1(net1244),
    .A2(_04976_),
    .B1(_04982_),
    .B2(\core.pipe1_resultRegister[0] ),
    .X(_04983_));
 sky130_fd_sc_hd__or2_1 _09996_ (.A(net1776),
    .B(\core.registers[20][0] ),
    .X(_04984_));
 sky130_fd_sc_hd__o221a_1 _09997_ (.A1(net1683),
    .A2(\core.registers[19][0] ),
    .B1(net1384),
    .B2(\core.registers[18][0] ),
    .C1(net1438),
    .X(_04985_));
 sky130_fd_sc_hd__o221a_1 _09998_ (.A1(net1683),
    .A2(\core.registers[23][0] ),
    .B1(net1385),
    .B2(\core.registers[22][0] ),
    .C1(net1450),
    .X(_04986_));
 sky130_fd_sc_hd__o221a_1 _09999_ (.A1(net1681),
    .A2(\core.registers[7][0] ),
    .B1(net1384),
    .B2(\core.registers[6][0] ),
    .C1(net1450),
    .X(_04987_));
 sky130_fd_sc_hd__o221a_1 _10000_ (.A1(net1683),
    .A2(\core.registers[3][0] ),
    .B1(net1387),
    .B2(\core.registers[2][0] ),
    .C1(net1438),
    .X(_04988_));
 sky130_fd_sc_hd__mux2_1 _10001_ (.A0(\core.registers[0][0] ),
    .A1(\core.registers[1][0] ),
    .S(net1387),
    .X(_04989_));
 sky130_fd_sc_hd__o221a_1 _10002_ (.A1(net1776),
    .A2(\core.registers[4][0] ),
    .B1(\core.registers[5][0] ),
    .B2(net1359),
    .C1(net1450),
    .X(_04990_));
 sky130_fd_sc_hd__a211o_1 _10003_ (.A1(net1438),
    .A2(_04989_),
    .B1(_04990_),
    .C1(net1346),
    .X(_04991_));
 sky130_fd_sc_hd__o311a_1 _10004_ (.A1(net1340),
    .A2(_04987_),
    .A3(_04988_),
    .B1(_04991_),
    .C1(net1320),
    .X(_04992_));
 sky130_fd_sc_hd__o211a_1 _10005_ (.A1(\core.registers[21][0] ),
    .A2(net1359),
    .B1(_04984_),
    .C1(net1450),
    .X(_04993_));
 sky130_fd_sc_hd__mux2_1 _10006_ (.A0(\core.registers[16][0] ),
    .A1(\core.registers[17][0] ),
    .S(net1388),
    .X(_04994_));
 sky130_fd_sc_hd__a211o_1 _10007_ (.A1(net1438),
    .A2(_04994_),
    .B1(_04993_),
    .C1(net1344),
    .X(_04995_));
 sky130_fd_sc_hd__o311a_1 _10008_ (.A1(net1331),
    .A2(_04985_),
    .A3(_04986_),
    .B1(_04995_),
    .C1(net1325),
    .X(_04996_));
 sky130_fd_sc_hd__or3_2 _10009_ (.A(_04076_),
    .B(_04992_),
    .C(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__mux2_1 _10010_ (.A0(\core.registers[10][0] ),
    .A1(\core.registers[11][0] ),
    .S(net1389),
    .X(_04998_));
 sky130_fd_sc_hd__mux2_1 _10011_ (.A0(\core.registers[8][0] ),
    .A1(\core.registers[9][0] ),
    .S(net1389),
    .X(_04999_));
 sky130_fd_sc_hd__mux2_1 _10012_ (.A0(_04998_),
    .A1(_04999_),
    .S(net1331),
    .X(_05000_));
 sky130_fd_sc_hd__mux2_1 _10013_ (.A0(\core.registers[14][0] ),
    .A1(\core.registers[15][0] ),
    .S(net1379),
    .X(_05001_));
 sky130_fd_sc_hd__mux2_1 _10014_ (.A0(\core.registers[12][0] ),
    .A1(\core.registers[13][0] ),
    .S(net1380),
    .X(_05002_));
 sky130_fd_sc_hd__mux2_1 _10015_ (.A0(_05001_),
    .A1(_05002_),
    .S(net1330),
    .X(_05003_));
 sky130_fd_sc_hd__o221a_1 _10016_ (.A1(net1763),
    .A2(_05000_),
    .B1(_05003_),
    .B2(net1436),
    .C1(net1320),
    .X(_05004_));
 sky130_fd_sc_hd__mux4_1 _10017_ (.A0(\core.registers[24][0] ),
    .A1(\core.registers[25][0] ),
    .A2(\core.registers[28][0] ),
    .A3(\core.registers[29][0] ),
    .S0(net1380),
    .S1(net1764),
    .X(_05005_));
 sky130_fd_sc_hd__a221o_1 _10018_ (.A1(net1681),
    .A2(\core.registers[30][0] ),
    .B1(\core.registers[31][0] ),
    .B2(net1384),
    .C1(net1705),
    .X(_05006_));
 sky130_fd_sc_hd__a221o_1 _10019_ (.A1(net1681),
    .A2(\core.registers[26][0] ),
    .B1(\core.registers[27][0] ),
    .B2(net1379),
    .C1(net1764),
    .X(_05007_));
 sky130_fd_sc_hd__and3_1 _10020_ (.A(net1770),
    .B(_05006_),
    .C(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__a21o_1 _10021_ (.A1(net1700),
    .A2(_05005_),
    .B1(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__a211o_1 _10022_ (.A1(net1755),
    .A2(_05009_),
    .B1(_05004_),
    .C1(net1427),
    .X(_05010_));
 sky130_fd_sc_hd__a21o_2 _10023_ (.A1(_04997_),
    .A2(_05010_),
    .B1(net1148),
    .X(_05011_));
 sky130_fd_sc_hd__o211ai_4 _10024_ (.A1(net1142),
    .A2(net1079),
    .B1(_05011_),
    .C1(net1240),
    .Y(_05012_));
 sky130_fd_sc_hd__nor2_1 _10025_ (.A(\core.pipe0_currentInstruction[7] ),
    .B(net1154),
    .Y(_05013_));
 sky130_fd_sc_hd__a211o_1 _10026_ (.A1(net1154),
    .A2(_05012_),
    .B1(_05013_),
    .C1(net1093),
    .X(_05014_));
 sky130_fd_sc_hd__nand2_1 _10027_ (.A(net1776),
    .B(net1093),
    .Y(_05015_));
 sky130_fd_sc_hd__a21o_1 _10028_ (.A1(_05014_),
    .A2(_05015_),
    .B1(net1263),
    .X(_05016_));
 sky130_fd_sc_hd__mux2_1 _10029_ (.A0(\core.registers[28][0] ),
    .A1(\core.registers[29][0] ),
    .S(net1479),
    .X(_05017_));
 sky130_fd_sc_hd__a221o_1 _10030_ (.A1(net1647),
    .A2(\core.registers[30][0] ),
    .B1(\core.registers[31][0] ),
    .B2(net1483),
    .C1(net1667),
    .X(_05018_));
 sky130_fd_sc_hd__mux2_1 _10031_ (.A0(\core.registers[8][0] ),
    .A1(\core.registers[9][0] ),
    .S(net1486),
    .X(_05019_));
 sky130_fd_sc_hd__mux2_1 _10032_ (.A0(\core.registers[10][0] ),
    .A1(\core.registers[11][0] ),
    .S(net1486),
    .X(_05020_));
 sky130_fd_sc_hd__mux2_1 _10033_ (.A0(_05019_),
    .A1(_05020_),
    .S(net1549),
    .X(_05021_));
 sky130_fd_sc_hd__mux2_1 _10034_ (.A0(\core.registers[24][0] ),
    .A1(\core.registers[25][0] ),
    .S(net1489),
    .X(_05022_));
 sky130_fd_sc_hd__a22o_1 _10035_ (.A1(net1649),
    .A2(\core.registers[26][0] ),
    .B1(\core.registers[27][0] ),
    .B2(net1479),
    .X(_05023_));
 sky130_fd_sc_hd__mux2_1 _10036_ (.A0(_05022_),
    .A1(_05023_),
    .S(net1788),
    .X(_05024_));
 sky130_fd_sc_hd__mux2_1 _10037_ (.A0(_05021_),
    .A1(_05024_),
    .S(net1779),
    .X(_05025_));
 sky130_fd_sc_hd__mux2_1 _10038_ (.A0(\core.registers[12][0] ),
    .A1(\core.registers[13][0] ),
    .S(net1478),
    .X(_05026_));
 sky130_fd_sc_hd__mux2_1 _10039_ (.A0(\core.registers[14][0] ),
    .A1(\core.registers[15][0] ),
    .S(net1478),
    .X(_05027_));
 sky130_fd_sc_hd__mux2_1 _10040_ (.A0(_05026_),
    .A1(_05027_),
    .S(net1546),
    .X(_05028_));
 sky130_fd_sc_hd__nor2_1 _10041_ (.A(net1779),
    .B(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__o21ai_1 _10042_ (.A1(net1788),
    .A2(_05017_),
    .B1(_05018_),
    .Y(_05030_));
 sky130_fd_sc_hd__a211o_1 _10043_ (.A1(net1779),
    .A2(_05030_),
    .B1(_05029_),
    .C1(net1669),
    .X(_05031_));
 sky130_fd_sc_hd__a21oi_1 _10044_ (.A1(net1669),
    .A2(_05025_),
    .B1(net1562),
    .Y(_05032_));
 sky130_fd_sc_hd__mux2_1 _10045_ (.A0(\core.registers[18][0] ),
    .A1(\core.registers[19][0] ),
    .S(net1483),
    .X(_05033_));
 sky130_fd_sc_hd__mux2_1 _10046_ (.A0(\core.registers[16][0] ),
    .A1(\core.registers[17][0] ),
    .S(net1484),
    .X(_05034_));
 sky130_fd_sc_hd__mux2_1 _10047_ (.A0(_05033_),
    .A1(_05034_),
    .S(net1531),
    .X(_05035_));
 sky130_fd_sc_hd__o221a_1 _10048_ (.A1(net1649),
    .A2(\core.registers[23][0] ),
    .B1(net1484),
    .B2(\core.registers[22][0] ),
    .C1(net1547),
    .X(_05036_));
 sky130_fd_sc_hd__mux2_1 _10049_ (.A0(\core.registers[20][0] ),
    .A1(\core.registers[21][0] ),
    .S(net1484),
    .X(_05037_));
 sky130_fd_sc_hd__or2_1 _10050_ (.A(\core.registers[0][0] ),
    .B(net1487),
    .X(_05038_));
 sky130_fd_sc_hd__o211a_1 _10051_ (.A1(\core.registers[1][0] ),
    .A2(net1459),
    .B1(_05038_),
    .C1(net1532),
    .X(_05039_));
 sky130_fd_sc_hd__mux2_1 _10052_ (.A0(\core.registers[2][0] ),
    .A1(\core.registers[3][0] ),
    .S(net1487),
    .X(_05040_));
 sky130_fd_sc_hd__a211o_1 _10053_ (.A1(net1549),
    .A2(_05040_),
    .B1(_05039_),
    .C1(net1586),
    .X(_05041_));
 sky130_fd_sc_hd__mux2_1 _10054_ (.A0(\core.registers[4][0] ),
    .A1(\core.registers[5][0] ),
    .S(net1487),
    .X(_05042_));
 sky130_fd_sc_hd__o221a_1 _10055_ (.A1(net1649),
    .A2(\core.registers[7][0] ),
    .B1(net1483),
    .B2(\core.registers[6][0] ),
    .C1(net1547),
    .X(_05043_));
 sky130_fd_sc_hd__a211o_1 _10056_ (.A1(net1530),
    .A2(_05042_),
    .B1(_05043_),
    .C1(net1574),
    .X(_05044_));
 sky130_fd_sc_hd__a211o_1 _10057_ (.A1(net1531),
    .A2(_05037_),
    .B1(_05036_),
    .C1(net1575),
    .X(_05045_));
 sky130_fd_sc_hd__o211a_1 _10058_ (.A1(net1586),
    .A2(_05035_),
    .B1(_05045_),
    .C1(net1598),
    .X(_05046_));
 sky130_fd_sc_hd__a31o_1 _10059_ (.A1(net1594),
    .A2(_05041_),
    .A3(_05044_),
    .B1(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__o2bb2a_1 _10060_ (.A1_N(_05031_),
    .A2_N(_05032_),
    .B1(_05047_),
    .B2(net1567),
    .X(_05048_));
 sky130_fd_sc_hd__a22o_2 _10061_ (.A1(net1094),
    .A2(net1079),
    .B1(_05048_),
    .B2(net1046),
    .X(_05049_));
 sky130_fd_sc_hd__mux2_8 _10062_ (.A0(net450),
    .A1(_05049_),
    .S(net1258),
    .X(_05050_));
 sky130_fd_sc_hd__and2b_1 _10063_ (.A_N(net885),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__nand2b_1 _10064_ (.A_N(net885),
    .B(_05050_),
    .Y(_05052_));
 sky130_fd_sc_hd__nor2_2 _10065_ (.A(_04972_),
    .B(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__nor2_4 _10066_ (.A(_04970_),
    .B(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__a211o_1 _10067_ (.A1(_04971_),
    .A2(_05051_),
    .B1(_04885_),
    .C1(_04970_),
    .X(_05055_));
 sky130_fd_sc_hd__nand2_2 _10068_ (.A(_04886_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__a21o_1 _10069_ (.A1(_04886_),
    .A2(_05055_),
    .B1(_04806_),
    .X(_05057_));
 sky130_fd_sc_hd__nand2_2 _10070_ (.A(_04805_),
    .B(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__a31o_4 _10071_ (.A1(_04723_),
    .A2(_04805_),
    .A3(_05057_),
    .B1(_04722_),
    .X(_05059_));
 sky130_fd_sc_hd__a21oi_4 _10072_ (.A1(_04635_),
    .A2(_05059_),
    .B1(_04633_),
    .Y(_05060_));
 sky130_fd_sc_hd__a211o_1 _10073_ (.A1(_04635_),
    .A2(_05059_),
    .B1(_04548_),
    .C1(_04633_),
    .X(_05061_));
 sky130_fd_sc_hd__nand2_2 _10074_ (.A(_04549_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__a21oi_1 _10075_ (.A1(_04549_),
    .A2(_05061_),
    .B1(_04462_),
    .Y(_05063_));
 sky130_fd_sc_hd__or2_4 _10076_ (.A(_04463_),
    .B(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__o21ai_4 _10077_ (.A1(_04392_),
    .A2(_05064_),
    .B1(_04389_),
    .Y(_05065_));
 sky130_fd_sc_hd__a21boi_4 _10078_ (.A1(_04307_),
    .A2(_05065_),
    .B1_N(_04304_),
    .Y(_05066_));
 sky130_fd_sc_hd__o21ba_4 _10079_ (.A1(_04218_),
    .A2(_05066_),
    .B1_N(_04216_),
    .X(_05067_));
 sky130_fd_sc_hd__xnor2_4 _10080_ (.A(_04133_),
    .B(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__a21o_1 _10081_ (.A1(net1751),
    .A2(net1039),
    .B1(net1263),
    .X(_05069_));
 sky130_fd_sc_hd__a21o_1 _10082_ (.A1(\core.pipe1_csrData[30] ),
    .A2(net1250),
    .B1(net1237),
    .X(_05070_));
 sky130_fd_sc_hd__a31o_1 _10083_ (.A1(net1616),
    .A2(_04006_),
    .A3(_04012_),
    .B1(net1242),
    .X(_05071_));
 sky130_fd_sc_hd__nor2_1 _10084_ (.A(_03986_),
    .B(_04473_),
    .Y(_05072_));
 sky130_fd_sc_hd__nand2_2 _10085_ (.A(net1617),
    .B(_04014_),
    .Y(_05073_));
 sky130_fd_sc_hd__nor2_1 _10086_ (.A(_05072_),
    .B(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__o21a_1 _10087_ (.A1(net1186),
    .A2(_05074_),
    .B1(_05070_),
    .X(_05075_));
 sky130_fd_sc_hd__o22a_4 _10088_ (.A1(\core.pipe1_resultRegister[30] ),
    .A2(_03934_),
    .B1(_05075_),
    .B2(net1245),
    .X(_05076_));
 sky130_fd_sc_hd__nor2_1 _10089_ (.A(net1144),
    .B(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__mux2_1 _10090_ (.A0(\core.registers[12][30] ),
    .A1(\core.registers[13][30] ),
    .S(net1414),
    .X(_05078_));
 sky130_fd_sc_hd__mux2_1 _10091_ (.A0(\core.registers[14][30] ),
    .A1(\core.registers[15][30] ),
    .S(net1409),
    .X(_05079_));
 sky130_fd_sc_hd__mux2_1 _10092_ (.A0(_05078_),
    .A1(_05079_),
    .S(net1350),
    .X(_05080_));
 sky130_fd_sc_hd__nor2_1 _10093_ (.A(net1759),
    .B(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__a221o_1 _10094_ (.A1(net1691),
    .A2(\core.registers[30][30] ),
    .B1(\core.registers[31][30] ),
    .B2(net1409),
    .C1(net1701),
    .X(_05082_));
 sky130_fd_sc_hd__mux2_1 _10095_ (.A0(\core.registers[28][30] ),
    .A1(\core.registers[29][30] ),
    .S(net1409),
    .X(_05083_));
 sky130_fd_sc_hd__o21ai_1 _10096_ (.A1(net1773),
    .A2(_05083_),
    .B1(_05082_),
    .Y(_05084_));
 sky130_fd_sc_hd__a211o_1 _10097_ (.A1(net1759),
    .A2(_05084_),
    .B1(_05081_),
    .C1(net1706),
    .X(_05085_));
 sky130_fd_sc_hd__mux2_1 _10098_ (.A0(\core.registers[8][30] ),
    .A1(\core.registers[9][30] ),
    .S(net1410),
    .X(_05086_));
 sky130_fd_sc_hd__mux2_1 _10099_ (.A0(\core.registers[10][30] ),
    .A1(\core.registers[11][30] ),
    .S(net1410),
    .X(_05087_));
 sky130_fd_sc_hd__mux2_2 _10100_ (.A0(_05086_),
    .A1(_05087_),
    .S(net1350),
    .X(_05088_));
 sky130_fd_sc_hd__or2_1 _10101_ (.A(\core.registers[25][30] ),
    .B(net1361),
    .X(_05089_));
 sky130_fd_sc_hd__o211a_1 _10102_ (.A1(\core.registers[24][30] ),
    .A2(net1408),
    .B1(_05089_),
    .C1(net1701),
    .X(_05090_));
 sky130_fd_sc_hd__and3_1 _10103_ (.A(net1773),
    .B(\core.registers[27][30] ),
    .C(net1408),
    .X(_05091_));
 sky130_fd_sc_hd__a211o_1 _10104_ (.A1(\core.registers[26][30] ),
    .A2(net1319),
    .B1(_05091_),
    .C1(net1710),
    .X(_05092_));
 sky130_fd_sc_hd__o221ai_4 _10105_ (.A1(net1759),
    .A2(_05088_),
    .B1(_05090_),
    .B2(_05092_),
    .C1(net1706),
    .Y(_05093_));
 sky130_fd_sc_hd__mux4_1 _10106_ (.A0(\core.registers[16][30] ),
    .A1(\core.registers[17][30] ),
    .A2(\core.registers[20][30] ),
    .A3(\core.registers[21][30] ),
    .S0(net1414),
    .S1(net1454),
    .X(_05094_));
 sky130_fd_sc_hd__o22a_1 _10107_ (.A1(net1694),
    .A2(\core.registers[23][30] ),
    .B1(net1414),
    .B2(\core.registers[22][30] ),
    .X(_05095_));
 sky130_fd_sc_hd__o22a_1 _10108_ (.A1(net1694),
    .A2(\core.registers[19][30] ),
    .B1(net1414),
    .B2(\core.registers[18][30] ),
    .X(_05096_));
 sky130_fd_sc_hd__mux2_1 _10109_ (.A0(_05095_),
    .A1(_05096_),
    .S(net1443),
    .X(_05097_));
 sky130_fd_sc_hd__o21a_1 _10110_ (.A1(net1336),
    .A2(_05097_),
    .B1(net1326),
    .X(_05098_));
 sky130_fd_sc_hd__o21ai_2 _10111_ (.A1(net1350),
    .A2(_05094_),
    .B1(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__o22a_1 _10112_ (.A1(net1691),
    .A2(\core.registers[7][30] ),
    .B1(net1408),
    .B2(\core.registers[6][30] ),
    .X(_05100_));
 sky130_fd_sc_hd__o22a_1 _10113_ (.A1(net1691),
    .A2(\core.registers[3][30] ),
    .B1(net1408),
    .B2(\core.registers[2][30] ),
    .X(_05101_));
 sky130_fd_sc_hd__mux2_1 _10114_ (.A0(_05100_),
    .A1(_05101_),
    .S(net1443),
    .X(_05102_));
 sky130_fd_sc_hd__or2_1 _10115_ (.A(net1335),
    .B(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__mux4_1 _10116_ (.A0(\core.registers[0][30] ),
    .A1(\core.registers[1][30] ),
    .A2(\core.registers[4][30] ),
    .A3(\core.registers[5][30] ),
    .S0(net1411),
    .S1(net1454),
    .X(_05104_));
 sky130_fd_sc_hd__o21a_1 _10117_ (.A1(net1350),
    .A2(_05104_),
    .B1(net1322),
    .X(_05105_));
 sky130_fd_sc_hd__a21oi_1 _10118_ (.A1(_05103_),
    .A2(_05105_),
    .B1(net1433),
    .Y(_05106_));
 sky130_fd_sc_hd__a32o_4 _10119_ (.A1(net1433),
    .A2(_05085_),
    .A3(_05093_),
    .B1(_05099_),
    .B2(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__a211o_4 _10120_ (.A1(net1144),
    .A2(_05107_),
    .B1(_05077_),
    .C1(_04095_),
    .X(_05108_));
 sky130_fd_sc_hd__nor2_1 _10121_ (.A(net1040),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__o22a_2 _10122_ (.A1(net1752),
    .A2(net1257),
    .B1(net1006),
    .B2(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__mux2_1 _10123_ (.A0(\core.registers[18][30] ),
    .A1(\core.registers[19][30] ),
    .S(net1510),
    .X(_05111_));
 sky130_fd_sc_hd__mux2_1 _10124_ (.A0(\core.registers[16][30] ),
    .A1(\core.registers[17][30] ),
    .S(net1510),
    .X(_05112_));
 sky130_fd_sc_hd__mux2_1 _10125_ (.A0(_05111_),
    .A1(_05112_),
    .S(net1536),
    .X(_05113_));
 sky130_fd_sc_hd__o221a_1 _10126_ (.A1(net1656),
    .A2(\core.registers[23][30] ),
    .B1(net1510),
    .B2(\core.registers[22][30] ),
    .C1(net1556),
    .X(_05114_));
 sky130_fd_sc_hd__mux2_1 _10127_ (.A0(\core.registers[20][30] ),
    .A1(\core.registers[21][30] ),
    .S(net1510),
    .X(_05115_));
 sky130_fd_sc_hd__or2_1 _10128_ (.A(\core.registers[0][30] ),
    .B(net1509),
    .X(_05116_));
 sky130_fd_sc_hd__o211a_1 _10129_ (.A1(\core.registers[1][30] ),
    .A2(net1460),
    .B1(_05116_),
    .C1(net1537),
    .X(_05117_));
 sky130_fd_sc_hd__mux2_1 _10130_ (.A0(\core.registers[2][30] ),
    .A1(\core.registers[3][30] ),
    .S(net1506),
    .X(_05118_));
 sky130_fd_sc_hd__a211o_1 _10131_ (.A1(net1555),
    .A2(_05118_),
    .B1(_05117_),
    .C1(net1589),
    .X(_05119_));
 sky130_fd_sc_hd__mux2_1 _10132_ (.A0(\core.registers[4][30] ),
    .A1(\core.registers[5][30] ),
    .S(net1507),
    .X(_05120_));
 sky130_fd_sc_hd__o221a_1 _10133_ (.A1(net1656),
    .A2(\core.registers[7][30] ),
    .B1(net1507),
    .B2(\core.registers[6][30] ),
    .C1(net1555),
    .X(_05121_));
 sky130_fd_sc_hd__a211o_1 _10134_ (.A1(net1537),
    .A2(_05120_),
    .B1(_05121_),
    .C1(net1580),
    .X(_05122_));
 sky130_fd_sc_hd__a211o_1 _10135_ (.A1(net1536),
    .A2(_05115_),
    .B1(_05114_),
    .C1(net1580),
    .X(_05123_));
 sky130_fd_sc_hd__o211a_1 _10136_ (.A1(net1589),
    .A2(_05113_),
    .B1(_05123_),
    .C1(net1599),
    .X(_05124_));
 sky130_fd_sc_hd__a311o_2 _10137_ (.A1(net1595),
    .A2(_05119_),
    .A3(_05122_),
    .B1(_05124_),
    .C1(net1568),
    .X(_05125_));
 sky130_fd_sc_hd__mux2_1 _10138_ (.A0(\core.registers[28][30] ),
    .A1(\core.registers[29][30] ),
    .S(net1507),
    .X(_05126_));
 sky130_fd_sc_hd__a221o_1 _10139_ (.A1(net1656),
    .A2(\core.registers[30][30] ),
    .B1(\core.registers[31][30] ),
    .B2(net1506),
    .C1(net1664),
    .X(_05127_));
 sky130_fd_sc_hd__mux2_1 _10140_ (.A0(\core.registers[8][30] ),
    .A1(\core.registers[9][30] ),
    .S(net1508),
    .X(_05128_));
 sky130_fd_sc_hd__mux2_1 _10141_ (.A0(\core.registers[10][30] ),
    .A1(\core.registers[11][30] ),
    .S(net1508),
    .X(_05129_));
 sky130_fd_sc_hd__mux2_1 _10142_ (.A0(_05128_),
    .A1(_05129_),
    .S(net1555),
    .X(_05130_));
 sky130_fd_sc_hd__or2_1 _10143_ (.A(\core.registers[25][30] ),
    .B(net1461),
    .X(_05131_));
 sky130_fd_sc_hd__o21a_1 _10144_ (.A1(\core.registers[24][30] ),
    .A2(net1506),
    .B1(net1665),
    .X(_05132_));
 sky130_fd_sc_hd__a22o_1 _10145_ (.A1(net1656),
    .A2(\core.registers[26][30] ),
    .B1(\core.registers[27][30] ),
    .B2(net1506),
    .X(_05133_));
 sky130_fd_sc_hd__a221o_1 _10146_ (.A1(_05131_),
    .A2(_05132_),
    .B1(_05133_),
    .B2(net1790),
    .C1(net1672),
    .X(_05134_));
 sky130_fd_sc_hd__o211a_1 _10147_ (.A1(net1781),
    .A2(_05130_),
    .B1(_05134_),
    .C1(net1670),
    .X(_05135_));
 sky130_fd_sc_hd__o21a_1 _10148_ (.A1(net1790),
    .A2(_05126_),
    .B1(_05127_),
    .X(_05136_));
 sky130_fd_sc_hd__mux2_1 _10149_ (.A0(\core.registers[12][30] ),
    .A1(\core.registers[13][30] ),
    .S(net1510),
    .X(_05137_));
 sky130_fd_sc_hd__mux2_1 _10150_ (.A0(\core.registers[14][30] ),
    .A1(\core.registers[15][30] ),
    .S(net1507),
    .X(_05138_));
 sky130_fd_sc_hd__mux2_1 _10151_ (.A0(_05137_),
    .A1(_05138_),
    .S(net1555),
    .X(_05139_));
 sky130_fd_sc_hd__mux2_1 _10152_ (.A0(_05136_),
    .A1(_05139_),
    .S(net1672),
    .X(_05140_));
 sky130_fd_sc_hd__a21o_1 _10153_ (.A1(net1785),
    .A2(_05140_),
    .B1(net1564),
    .X(_05141_));
 sky130_fd_sc_hd__o21ai_4 _10154_ (.A1(_05135_),
    .A2(_05141_),
    .B1(_05125_),
    .Y(_05142_));
 sky130_fd_sc_hd__o2bb2a_4 _10155_ (.A1_N(net1095),
    .A2_N(_05076_),
    .B1(_05142_),
    .B2(net1044),
    .X(_05143_));
 sky130_fd_sc_hd__inv_2 _10156_ (.A(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__mux2_4 _10157_ (.A0(net473),
    .A1(_05144_),
    .S(net1255),
    .X(_05145_));
 sky130_fd_sc_hd__and2_2 _10158_ (.A(_05110_),
    .B(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__nor2_1 _10159_ (.A(_05110_),
    .B(_05145_),
    .Y(_05147_));
 sky130_fd_sc_hd__or2_4 _10160_ (.A(_05146_),
    .B(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__inv_6 _10161_ (.A(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__nor2_1 _10162_ (.A(_03986_),
    .B(_04558_),
    .Y(_05150_));
 sky130_fd_sc_hd__nor2_1 _10163_ (.A(_05073_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__a21o_1 _10164_ (.A1(\core.pipe1_csrData[29] ),
    .A2(net1250),
    .B1(net1237),
    .X(_05152_));
 sky130_fd_sc_hd__o21a_1 _10165_ (.A1(net1187),
    .A2(_05151_),
    .B1(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__o22a_4 _10166_ (.A1(\core.pipe1_resultRegister[29] ),
    .A2(_03934_),
    .B1(_05153_),
    .B2(net1245),
    .X(_05154_));
 sky130_fd_sc_hd__mux2_1 _10167_ (.A0(\core.registers[14][29] ),
    .A1(\core.registers[15][29] ),
    .S(net1409),
    .X(_05155_));
 sky130_fd_sc_hd__mux2_1 _10168_ (.A0(\core.registers[12][29] ),
    .A1(\core.registers[13][29] ),
    .S(net1409),
    .X(_05156_));
 sky130_fd_sc_hd__mux2_1 _10169_ (.A0(_05155_),
    .A1(_05156_),
    .S(net1335),
    .X(_05157_));
 sky130_fd_sc_hd__mux2_1 _10170_ (.A0(\core.registers[28][29] ),
    .A1(\core.registers[29][29] ),
    .S(net1408),
    .X(_05158_));
 sky130_fd_sc_hd__a221o_1 _10171_ (.A1(net1691),
    .A2(\core.registers[30][29] ),
    .B1(\core.registers[31][29] ),
    .B2(net1408),
    .C1(net1701),
    .X(_05159_));
 sky130_fd_sc_hd__o21a_1 _10172_ (.A1(net1773),
    .A2(_05158_),
    .B1(_05159_),
    .X(_05160_));
 sky130_fd_sc_hd__mux2_1 _10173_ (.A0(\core.registers[8][29] ),
    .A1(\core.registers[9][29] ),
    .S(net1408),
    .X(_05161_));
 sky130_fd_sc_hd__mux2_1 _10174_ (.A0(\core.registers[10][29] ),
    .A1(\core.registers[11][29] ),
    .S(net1408),
    .X(_05162_));
 sky130_fd_sc_hd__mux2_1 _10175_ (.A0(_05161_),
    .A1(_05162_),
    .S(net1350),
    .X(_05163_));
 sky130_fd_sc_hd__mux2_1 _10176_ (.A0(\core.registers[24][29] ),
    .A1(\core.registers[25][29] ),
    .S(net1408),
    .X(_05164_));
 sky130_fd_sc_hd__a22o_1 _10177_ (.A1(net1691),
    .A2(\core.registers[26][29] ),
    .B1(\core.registers[27][29] ),
    .B2(net1408),
    .X(_05165_));
 sky130_fd_sc_hd__mux2_1 _10178_ (.A0(_05164_),
    .A1(_05165_),
    .S(net1773),
    .X(_05166_));
 sky130_fd_sc_hd__mux4_2 _10179_ (.A0(_05157_),
    .A1(_05160_),
    .A2(_05163_),
    .A3(_05166_),
    .S0(net1759),
    .S1(net1706),
    .X(_05167_));
 sky130_fd_sc_hd__nand2_1 _10180_ (.A(net1432),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__mux4_1 _10181_ (.A0(\core.registers[16][29] ),
    .A1(\core.registers[17][29] ),
    .A2(\core.registers[20][29] ),
    .A3(\core.registers[21][29] ),
    .S0(net1414),
    .S1(net1454),
    .X(_05169_));
 sky130_fd_sc_hd__o22a_1 _10182_ (.A1(net1694),
    .A2(\core.registers[23][29] ),
    .B1(net1414),
    .B2(\core.registers[22][29] ),
    .X(_05170_));
 sky130_fd_sc_hd__o22a_1 _10183_ (.A1(net1694),
    .A2(\core.registers[19][29] ),
    .B1(net1414),
    .B2(\core.registers[18][29] ),
    .X(_05171_));
 sky130_fd_sc_hd__mux2_1 _10184_ (.A0(_05170_),
    .A1(_05171_),
    .S(net1443),
    .X(_05172_));
 sky130_fd_sc_hd__o21a_1 _10185_ (.A1(net1336),
    .A2(_05172_),
    .B1(net1326),
    .X(_05173_));
 sky130_fd_sc_hd__o21a_1 _10186_ (.A1(net1350),
    .A2(_05169_),
    .B1(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__o22a_1 _10187_ (.A1(net1694),
    .A2(\core.registers[7][29] ),
    .B1(net1414),
    .B2(\core.registers[6][29] ),
    .X(_05175_));
 sky130_fd_sc_hd__o22a_1 _10188_ (.A1(net1694),
    .A2(\core.registers[3][29] ),
    .B1(net1414),
    .B2(\core.registers[2][29] ),
    .X(_05176_));
 sky130_fd_sc_hd__mux2_1 _10189_ (.A0(_05175_),
    .A1(_05176_),
    .S(net1443),
    .X(_05177_));
 sky130_fd_sc_hd__or2_2 _10190_ (.A(net1336),
    .B(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__mux4_1 _10191_ (.A0(\core.registers[0][29] ),
    .A1(\core.registers[1][29] ),
    .A2(\core.registers[4][29] ),
    .A3(\core.registers[5][29] ),
    .S0(net1414),
    .S1(net1454),
    .X(_05179_));
 sky130_fd_sc_hd__o21a_1 _10192_ (.A1(net1351),
    .A2(_05179_),
    .B1(net1322),
    .X(_05180_));
 sky130_fd_sc_hd__a21oi_4 _10193_ (.A1(_05178_),
    .A2(_05180_),
    .B1(_05174_),
    .Y(_05181_));
 sky130_fd_sc_hd__o211ai_4 _10194_ (.A1(net1432),
    .A2(_05181_),
    .B1(_05168_),
    .C1(net1147),
    .Y(_05182_));
 sky130_fd_sc_hd__o211ai_4 _10195_ (.A1(net1144),
    .A2(_05154_),
    .B1(_05182_),
    .C1(net1241),
    .Y(_05183_));
 sky130_fd_sc_hd__nor2_1 _10196_ (.A(net1041),
    .B(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__o22a_4 _10197_ (.A1(\core.pipe0_currentInstruction[29] ),
    .A2(net1257),
    .B1(net1006),
    .B2(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__mux2_1 _10198_ (.A0(\core.registers[18][29] ),
    .A1(\core.registers[19][29] ),
    .S(net1510),
    .X(_05186_));
 sky130_fd_sc_hd__mux2_1 _10199_ (.A0(\core.registers[16][29] ),
    .A1(\core.registers[17][29] ),
    .S(net1513),
    .X(_05187_));
 sky130_fd_sc_hd__mux2_1 _10200_ (.A0(_05186_),
    .A1(_05187_),
    .S(net1536),
    .X(_05188_));
 sky130_fd_sc_hd__o221a_1 _10201_ (.A1(net1657),
    .A2(\core.registers[23][29] ),
    .B1(net1513),
    .B2(\core.registers[22][29] ),
    .C1(net1556),
    .X(_05189_));
 sky130_fd_sc_hd__mux2_1 _10202_ (.A0(\core.registers[20][29] ),
    .A1(\core.registers[21][29] ),
    .S(net1510),
    .X(_05190_));
 sky130_fd_sc_hd__mux2_1 _10203_ (.A0(\core.registers[0][29] ),
    .A1(\core.registers[1][29] ),
    .S(net1512),
    .X(_05191_));
 sky130_fd_sc_hd__mux2_1 _10204_ (.A0(\core.registers[2][29] ),
    .A1(\core.registers[3][29] ),
    .S(net1510),
    .X(_05192_));
 sky130_fd_sc_hd__mux2_1 _10205_ (.A0(_05191_),
    .A1(_05192_),
    .S(net1556),
    .X(_05193_));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(\core.registers[4][29] ),
    .A1(\core.registers[5][29] ),
    .S(net1510),
    .X(_05194_));
 sky130_fd_sc_hd__o221a_1 _10207_ (.A1(net1657),
    .A2(\core.registers[7][29] ),
    .B1(net1510),
    .B2(\core.registers[6][29] ),
    .C1(net1556),
    .X(_05195_));
 sky130_fd_sc_hd__a211o_1 _10208_ (.A1(net1536),
    .A2(_05194_),
    .B1(_05195_),
    .C1(net1580),
    .X(_05196_));
 sky130_fd_sc_hd__a211o_1 _10209_ (.A1(net1536),
    .A2(_05190_),
    .B1(_05189_),
    .C1(net1580),
    .X(_05197_));
 sky130_fd_sc_hd__o211a_2 _10210_ (.A1(net1589),
    .A2(_05188_),
    .B1(_05197_),
    .C1(net1599),
    .X(_05198_));
 sky130_fd_sc_hd__o211a_2 _10211_ (.A1(net1592),
    .A2(_05193_),
    .B1(_05196_),
    .C1(net1595),
    .X(_05199_));
 sky130_fd_sc_hd__mux2_1 _10212_ (.A0(\core.registers[28][29] ),
    .A1(\core.registers[29][29] ),
    .S(net1506),
    .X(_05200_));
 sky130_fd_sc_hd__a221o_1 _10213_ (.A1(net1656),
    .A2(\core.registers[30][29] ),
    .B1(\core.registers[31][29] ),
    .B2(net1506),
    .C1(net1664),
    .X(_05201_));
 sky130_fd_sc_hd__mux2_1 _10214_ (.A0(\core.registers[8][29] ),
    .A1(\core.registers[9][29] ),
    .S(net1506),
    .X(_05202_));
 sky130_fd_sc_hd__mux2_1 _10215_ (.A0(\core.registers[10][29] ),
    .A1(\core.registers[11][29] ),
    .S(net1506),
    .X(_05203_));
 sky130_fd_sc_hd__mux2_1 _10216_ (.A0(_05202_),
    .A1(_05203_),
    .S(net1555),
    .X(_05204_));
 sky130_fd_sc_hd__or2_1 _10217_ (.A(\core.registers[25][29] ),
    .B(net1461),
    .X(_05205_));
 sky130_fd_sc_hd__o21a_1 _10218_ (.A1(\core.registers[24][29] ),
    .A2(net1506),
    .B1(net1664),
    .X(_05206_));
 sky130_fd_sc_hd__a22o_1 _10219_ (.A1(net1656),
    .A2(\core.registers[26][29] ),
    .B1(\core.registers[27][29] ),
    .B2(net1506),
    .X(_05207_));
 sky130_fd_sc_hd__a221o_1 _10220_ (.A1(_05205_),
    .A2(_05206_),
    .B1(_05207_),
    .B2(net1790),
    .C1(net1672),
    .X(_05208_));
 sky130_fd_sc_hd__o211a_1 _10221_ (.A1(net1781),
    .A2(_05204_),
    .B1(_05208_),
    .C1(net1670),
    .X(_05209_));
 sky130_fd_sc_hd__o21a_1 _10222_ (.A1(net1790),
    .A2(_05200_),
    .B1(_05201_),
    .X(_05210_));
 sky130_fd_sc_hd__mux2_1 _10223_ (.A0(\core.registers[12][29] ),
    .A1(\core.registers[13][29] ),
    .S(net1507),
    .X(_05211_));
 sky130_fd_sc_hd__mux2_1 _10224_ (.A0(\core.registers[14][29] ),
    .A1(\core.registers[15][29] ),
    .S(net1507),
    .X(_05212_));
 sky130_fd_sc_hd__mux2_1 _10225_ (.A0(_05211_),
    .A1(_05212_),
    .S(net1555),
    .X(_05213_));
 sky130_fd_sc_hd__mux2_1 _10226_ (.A0(_05210_),
    .A1(_05213_),
    .S(net1672),
    .X(_05214_));
 sky130_fd_sc_hd__a21o_1 _10227_ (.A1(net1786),
    .A2(_05214_),
    .B1(net1564),
    .X(_05215_));
 sky130_fd_sc_hd__o32a_4 _10228_ (.A1(net1568),
    .A2(_05198_),
    .A3(_05199_),
    .B1(_05209_),
    .B2(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__a22o_4 _10229_ (.A1(net1096),
    .A2(_05154_),
    .B1(_05216_),
    .B2(net1046),
    .X(_05217_));
 sky130_fd_sc_hd__mux2_4 _10230_ (.A0(net471),
    .A1(_05217_),
    .S(net1254),
    .X(_05218_));
 sky130_fd_sc_hd__nor2_2 _10231_ (.A(_05185_),
    .B(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__inv_2 _10232_ (.A(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hd__and2_2 _10233_ (.A(_05185_),
    .B(_05218_),
    .X(_05221_));
 sky130_fd_sc_hd__nor2_1 _10234_ (.A(_03986_),
    .B(_04644_),
    .Y(_05222_));
 sky130_fd_sc_hd__nor2_1 _10235_ (.A(_05073_),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__a21o_1 _10236_ (.A1(\core.pipe1_csrData[28] ),
    .A2(net1250),
    .B1(net1237),
    .X(_05224_));
 sky130_fd_sc_hd__o21a_1 _10237_ (.A1(net1187),
    .A2(_05223_),
    .B1(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__o22a_2 _10238_ (.A1(\core.pipe1_resultRegister[28] ),
    .A2(net1188),
    .B1(_05225_),
    .B2(net1245),
    .X(_05226_));
 sky130_fd_sc_hd__nor2_1 _10239_ (.A(net1145),
    .B(net872),
    .Y(_05227_));
 sky130_fd_sc_hd__mux2_1 _10240_ (.A0(\core.registers[12][28] ),
    .A1(\core.registers[13][28] ),
    .S(net1397),
    .X(_05228_));
 sky130_fd_sc_hd__mux2_1 _10241_ (.A0(\core.registers[14][28] ),
    .A1(\core.registers[15][28] ),
    .S(net1397),
    .X(_05229_));
 sky130_fd_sc_hd__mux2_1 _10242_ (.A0(_05228_),
    .A1(_05229_),
    .S(net1350),
    .X(_05230_));
 sky130_fd_sc_hd__nor2_1 _10243_ (.A(net1759),
    .B(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__a221o_1 _10244_ (.A1(net1688),
    .A2(\core.registers[30][28] ),
    .B1(\core.registers[31][28] ),
    .B2(net1397),
    .C1(net1701),
    .X(_05232_));
 sky130_fd_sc_hd__mux2_1 _10245_ (.A0(\core.registers[28][28] ),
    .A1(\core.registers[29][28] ),
    .S(net1397),
    .X(_05233_));
 sky130_fd_sc_hd__o21ai_1 _10246_ (.A1(net1773),
    .A2(_05233_),
    .B1(_05232_),
    .Y(_05234_));
 sky130_fd_sc_hd__a211o_1 _10247_ (.A1(net1759),
    .A2(_05234_),
    .B1(_05231_),
    .C1(net1706),
    .X(_05235_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(\core.registers[8][28] ),
    .A1(\core.registers[9][28] ),
    .S(net1397),
    .X(_05236_));
 sky130_fd_sc_hd__mux2_1 _10249_ (.A0(\core.registers[10][28] ),
    .A1(\core.registers[11][28] ),
    .S(net1398),
    .X(_05237_));
 sky130_fd_sc_hd__mux2_2 _10250_ (.A0(_05236_),
    .A1(_05237_),
    .S(net1350),
    .X(_05238_));
 sky130_fd_sc_hd__or2_1 _10251_ (.A(\core.registers[24][28] ),
    .B(net1397),
    .X(_05239_));
 sky130_fd_sc_hd__o211a_1 _10252_ (.A1(\core.registers[25][28] ),
    .A2(net1362),
    .B1(_05239_),
    .C1(net1701),
    .X(_05240_));
 sky130_fd_sc_hd__and3_1 _10253_ (.A(net1773),
    .B(\core.registers[27][28] ),
    .C(net1397),
    .X(_05241_));
 sky130_fd_sc_hd__a211o_1 _10254_ (.A1(\core.registers[26][28] ),
    .A2(net1319),
    .B1(_05241_),
    .C1(net1710),
    .X(_05242_));
 sky130_fd_sc_hd__o221ai_4 _10255_ (.A1(net1759),
    .A2(_05238_),
    .B1(_05240_),
    .B2(_05242_),
    .C1(net1706),
    .Y(_05243_));
 sky130_fd_sc_hd__mux4_1 _10256_ (.A0(\core.registers[16][28] ),
    .A1(\core.registers[17][28] ),
    .A2(\core.registers[20][28] ),
    .A3(\core.registers[21][28] ),
    .S0(net1397),
    .S1(net1453),
    .X(_05244_));
 sky130_fd_sc_hd__o22a_1 _10257_ (.A1(net1688),
    .A2(\core.registers[23][28] ),
    .B1(net1397),
    .B2(\core.registers[22][28] ),
    .X(_05245_));
 sky130_fd_sc_hd__o22a_1 _10258_ (.A1(net1688),
    .A2(\core.registers[19][28] ),
    .B1(net1397),
    .B2(\core.registers[18][28] ),
    .X(_05246_));
 sky130_fd_sc_hd__mux2_1 _10259_ (.A0(_05245_),
    .A1(_05246_),
    .S(net1441),
    .X(_05247_));
 sky130_fd_sc_hd__o21a_1 _10260_ (.A1(net1332),
    .A2(_05247_),
    .B1(net1327),
    .X(_05248_));
 sky130_fd_sc_hd__o21ai_1 _10261_ (.A1(net1348),
    .A2(_05244_),
    .B1(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__o22a_1 _10262_ (.A1(net1689),
    .A2(\core.registers[7][28] ),
    .B1(net1400),
    .B2(\core.registers[6][28] ),
    .X(_05250_));
 sky130_fd_sc_hd__o22a_1 _10263_ (.A1(net1688),
    .A2(\core.registers[3][28] ),
    .B1(net1400),
    .B2(\core.registers[2][28] ),
    .X(_05251_));
 sky130_fd_sc_hd__mux2_1 _10264_ (.A0(_05250_),
    .A1(_05251_),
    .S(net1441),
    .X(_05252_));
 sky130_fd_sc_hd__or2_1 _10265_ (.A(net1334),
    .B(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__mux4_1 _10266_ (.A0(\core.registers[0][28] ),
    .A1(\core.registers[1][28] ),
    .A2(\core.registers[4][28] ),
    .A3(\core.registers[5][28] ),
    .S0(net1400),
    .S1(net1453),
    .X(_05254_));
 sky130_fd_sc_hd__o21a_1 _10267_ (.A1(net1348),
    .A2(_05254_),
    .B1(net1323),
    .X(_05255_));
 sky130_fd_sc_hd__a21oi_1 _10268_ (.A1(_05253_),
    .A2(_05255_),
    .B1(net1432),
    .Y(_05256_));
 sky130_fd_sc_hd__a32o_2 _10269_ (.A1(net1432),
    .A2(_05235_),
    .A3(_05243_),
    .B1(_05249_),
    .B2(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__a211o_4 _10270_ (.A1(net1145),
    .A2(_05257_),
    .B1(_05227_),
    .C1(_04095_),
    .X(_05258_));
 sky130_fd_sc_hd__nor2_1 _10271_ (.A(net1040),
    .B(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__o22a_2 _10272_ (.A1(\core.pipe0_currentInstruction[28] ),
    .A2(net1253),
    .B1(net1006),
    .B2(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__mux2_1 _10273_ (.A0(\core.registers[18][28] ),
    .A1(\core.registers[19][28] ),
    .S(net1495),
    .X(_05261_));
 sky130_fd_sc_hd__mux2_1 _10274_ (.A0(\core.registers[16][28] ),
    .A1(\core.registers[17][28] ),
    .S(net1495),
    .X(_05262_));
 sky130_fd_sc_hd__mux2_1 _10275_ (.A0(_05261_),
    .A1(_05262_),
    .S(net1534),
    .X(_05263_));
 sky130_fd_sc_hd__o221a_1 _10276_ (.A1(net1651),
    .A2(\core.registers[23][28] ),
    .B1(net1495),
    .B2(\core.registers[22][28] ),
    .C1(net1550),
    .X(_05264_));
 sky130_fd_sc_hd__mux2_1 _10277_ (.A0(\core.registers[20][28] ),
    .A1(\core.registers[21][28] ),
    .S(net1495),
    .X(_05265_));
 sky130_fd_sc_hd__mux2_1 _10278_ (.A0(\core.registers[0][28] ),
    .A1(\core.registers[1][28] ),
    .S(net1498),
    .X(_05266_));
 sky130_fd_sc_hd__mux2_1 _10279_ (.A0(\core.registers[2][28] ),
    .A1(\core.registers[3][28] ),
    .S(net1498),
    .X(_05267_));
 sky130_fd_sc_hd__mux2_1 _10280_ (.A0(_05266_),
    .A1(_05267_),
    .S(net1554),
    .X(_05268_));
 sky130_fd_sc_hd__mux2_1 _10281_ (.A0(\core.registers[4][28] ),
    .A1(\core.registers[5][28] ),
    .S(net1498),
    .X(_05269_));
 sky130_fd_sc_hd__o221a_1 _10282_ (.A1(net1655),
    .A2(\core.registers[7][28] ),
    .B1(net1498),
    .B2(\core.registers[6][28] ),
    .C1(net1550),
    .X(_05270_));
 sky130_fd_sc_hd__a211o_1 _10283_ (.A1(net1534),
    .A2(_05269_),
    .B1(_05270_),
    .C1(net1576),
    .X(_05271_));
 sky130_fd_sc_hd__a211o_1 _10284_ (.A1(net1534),
    .A2(_05265_),
    .B1(_05264_),
    .C1(net1576),
    .X(_05272_));
 sky130_fd_sc_hd__o211a_1 _10285_ (.A1(net1587),
    .A2(_05263_),
    .B1(_05272_),
    .C1(net1600),
    .X(_05273_));
 sky130_fd_sc_hd__o211a_1 _10286_ (.A1(net1587),
    .A2(_05268_),
    .B1(_05271_),
    .C1(net1596),
    .X(_05274_));
 sky130_fd_sc_hd__mux2_1 _10287_ (.A0(\core.registers[28][28] ),
    .A1(\core.registers[29][28] ),
    .S(net1495),
    .X(_05275_));
 sky130_fd_sc_hd__a221o_1 _10288_ (.A1(net1651),
    .A2(\core.registers[30][28] ),
    .B1(\core.registers[31][28] ),
    .B2(net1495),
    .C1(net1664),
    .X(_05276_));
 sky130_fd_sc_hd__mux2_1 _10289_ (.A0(\core.registers[8][28] ),
    .A1(\core.registers[9][28] ),
    .S(net1495),
    .X(_05277_));
 sky130_fd_sc_hd__mux2_1 _10290_ (.A0(\core.registers[10][28] ),
    .A1(\core.registers[11][28] ),
    .S(net1499),
    .X(_05278_));
 sky130_fd_sc_hd__mux2_1 _10291_ (.A0(_05277_),
    .A1(_05278_),
    .S(net1550),
    .X(_05279_));
 sky130_fd_sc_hd__or2_1 _10292_ (.A(\core.registers[25][28] ),
    .B(net1460),
    .X(_05280_));
 sky130_fd_sc_hd__o21a_1 _10293_ (.A1(\core.registers[24][28] ),
    .A2(net1499),
    .B1(net1664),
    .X(_05281_));
 sky130_fd_sc_hd__a22o_1 _10294_ (.A1(net1651),
    .A2(\core.registers[26][28] ),
    .B1(\core.registers[27][28] ),
    .B2(net1495),
    .X(_05282_));
 sky130_fd_sc_hd__a221o_1 _10295_ (.A1(_05280_),
    .A2(_05281_),
    .B1(_05282_),
    .B2(net1790),
    .C1(net1672),
    .X(_05283_));
 sky130_fd_sc_hd__o211a_1 _10296_ (.A1(net1781),
    .A2(_05279_),
    .B1(_05283_),
    .C1(net1670),
    .X(_05284_));
 sky130_fd_sc_hd__o21a_1 _10297_ (.A1(net1790),
    .A2(_05275_),
    .B1(_05276_),
    .X(_05285_));
 sky130_fd_sc_hd__mux2_1 _10298_ (.A0(\core.registers[12][28] ),
    .A1(\core.registers[13][28] ),
    .S(net1495),
    .X(_05286_));
 sky130_fd_sc_hd__mux2_1 _10299_ (.A0(\core.registers[14][28] ),
    .A1(\core.registers[15][28] ),
    .S(net1495),
    .X(_05287_));
 sky130_fd_sc_hd__mux2_1 _10300_ (.A0(_05286_),
    .A1(_05287_),
    .S(net1550),
    .X(_05288_));
 sky130_fd_sc_hd__mux2_1 _10301_ (.A0(_05285_),
    .A1(_05288_),
    .S(net1672),
    .X(_05289_));
 sky130_fd_sc_hd__a21o_1 _10302_ (.A1(net1785),
    .A2(_05289_),
    .B1(net1564),
    .X(_05290_));
 sky130_fd_sc_hd__o32a_4 _10303_ (.A1(net1569),
    .A2(_05273_),
    .A3(_05274_),
    .B1(_05284_),
    .B2(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__a22o_4 _10304_ (.A1(net1097),
    .A2(net872),
    .B1(_05291_),
    .B2(_03945_),
    .X(_05292_));
 sky130_fd_sc_hd__mux2_4 _10305_ (.A0(net470),
    .A1(_05292_),
    .S(net1254),
    .X(_05293_));
 sky130_fd_sc_hd__or2_4 _10306_ (.A(_05260_),
    .B(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__and2_2 _10307_ (.A(_05260_),
    .B(_05293_),
    .X(_05295_));
 sky130_fd_sc_hd__clkinv_2 _10308_ (.A(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__nor2_1 _10309_ (.A(_03987_),
    .B(_05073_),
    .Y(_05297_));
 sky130_fd_sc_hd__a21o_1 _10310_ (.A1(\core.pipe1_csrData[27] ),
    .A2(net1250),
    .B1(net1237),
    .X(_05298_));
 sky130_fd_sc_hd__o21a_1 _10311_ (.A1(net1187),
    .A2(_05297_),
    .B1(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__o22a_4 _10312_ (.A1(\core.pipe1_resultRegister[27] ),
    .A2(_03934_),
    .B1(_05299_),
    .B2(net1245),
    .X(_05300_));
 sky130_fd_sc_hd__mux2_1 _10313_ (.A0(\core.registers[14][27] ),
    .A1(\core.registers[15][27] ),
    .S(net1392),
    .X(_05301_));
 sky130_fd_sc_hd__mux2_1 _10314_ (.A0(\core.registers[12][27] ),
    .A1(\core.registers[13][27] ),
    .S(net1391),
    .X(_05302_));
 sky130_fd_sc_hd__mux2_1 _10315_ (.A0(_05301_),
    .A1(_05302_),
    .S(net1332),
    .X(_05303_));
 sky130_fd_sc_hd__mux2_1 _10316_ (.A0(\core.registers[28][27] ),
    .A1(\core.registers[29][27] ),
    .S(net1391),
    .X(_05304_));
 sky130_fd_sc_hd__a221o_1 _10317_ (.A1(net1687),
    .A2(\core.registers[30][27] ),
    .B1(\core.registers[31][27] ),
    .B2(net1391),
    .C1(net1702),
    .X(_05305_));
 sky130_fd_sc_hd__o21a_1 _10318_ (.A1(net1772),
    .A2(_05304_),
    .B1(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__mux2_1 _10319_ (.A0(\core.registers[8][27] ),
    .A1(\core.registers[9][27] ),
    .S(net1391),
    .X(_05307_));
 sky130_fd_sc_hd__mux2_1 _10320_ (.A0(\core.registers[10][27] ),
    .A1(\core.registers[11][27] ),
    .S(net1395),
    .X(_05308_));
 sky130_fd_sc_hd__mux2_1 _10321_ (.A0(_05307_),
    .A1(_05308_),
    .S(net1347),
    .X(_05309_));
 sky130_fd_sc_hd__mux2_1 _10322_ (.A0(\core.registers[24][27] ),
    .A1(\core.registers[25][27] ),
    .S(net1391),
    .X(_05310_));
 sky130_fd_sc_hd__a22o_1 _10323_ (.A1(net1687),
    .A2(\core.registers[26][27] ),
    .B1(\core.registers[27][27] ),
    .B2(net1391),
    .X(_05311_));
 sky130_fd_sc_hd__mux2_1 _10324_ (.A0(_05310_),
    .A1(_05311_),
    .S(net1772),
    .X(_05312_));
 sky130_fd_sc_hd__mux4_2 _10325_ (.A0(_05303_),
    .A1(_05306_),
    .A2(_05309_),
    .A3(_05312_),
    .S0(net1757),
    .S1(net1707),
    .X(_05313_));
 sky130_fd_sc_hd__nand2_1 _10326_ (.A(net1431),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__mux4_1 _10327_ (.A0(\core.registers[16][27] ),
    .A1(\core.registers[17][27] ),
    .A2(\core.registers[20][27] ),
    .A3(\core.registers[21][27] ),
    .S0(net1413),
    .S1(net1454),
    .X(_05315_));
 sky130_fd_sc_hd__o22a_1 _10328_ (.A1(net1694),
    .A2(\core.registers[23][27] ),
    .B1(net1412),
    .B2(\core.registers[22][27] ),
    .X(_05316_));
 sky130_fd_sc_hd__o22a_1 _10329_ (.A1(net1694),
    .A2(\core.registers[19][27] ),
    .B1(net1413),
    .B2(\core.registers[18][27] ),
    .X(_05317_));
 sky130_fd_sc_hd__mux2_1 _10330_ (.A0(_05316_),
    .A1(_05317_),
    .S(net1443),
    .X(_05318_));
 sky130_fd_sc_hd__o21a_1 _10331_ (.A1(net1336),
    .A2(_05318_),
    .B1(net1326),
    .X(_05319_));
 sky130_fd_sc_hd__o21a_2 _10332_ (.A1(net1351),
    .A2(_05315_),
    .B1(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__o22a_1 _10333_ (.A1(net1694),
    .A2(\core.registers[7][27] ),
    .B1(net1412),
    .B2(\core.registers[6][27] ),
    .X(_05321_));
 sky130_fd_sc_hd__o22a_1 _10334_ (.A1(net1694),
    .A2(\core.registers[3][27] ),
    .B1(net1412),
    .B2(\core.registers[2][27] ),
    .X(_05322_));
 sky130_fd_sc_hd__mux2_1 _10335_ (.A0(_05321_),
    .A1(_05322_),
    .S(net1443),
    .X(_05323_));
 sky130_fd_sc_hd__or2_2 _10336_ (.A(net1336),
    .B(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__mux4_1 _10337_ (.A0(\core.registers[0][27] ),
    .A1(\core.registers[1][27] ),
    .A2(\core.registers[4][27] ),
    .A3(\core.registers[5][27] ),
    .S0(net1412),
    .S1(net1457),
    .X(_05325_));
 sky130_fd_sc_hd__o21a_1 _10338_ (.A1(net1351),
    .A2(_05325_),
    .B1(net1322),
    .X(_05326_));
 sky130_fd_sc_hd__a21oi_4 _10339_ (.A1(_05324_),
    .A2(_05326_),
    .B1(_05320_),
    .Y(_05327_));
 sky130_fd_sc_hd__o211ai_4 _10340_ (.A1(net1431),
    .A2(_05327_),
    .B1(_05314_),
    .C1(net1146),
    .Y(_05328_));
 sky130_fd_sc_hd__o211ai_4 _10341_ (.A1(net1146),
    .A2(net868),
    .B1(_05328_),
    .C1(net1240),
    .Y(_05329_));
 sky130_fd_sc_hd__nor2_1 _10342_ (.A(net1041),
    .B(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__o22a_4 _10343_ (.A1(\core.pipe0_currentInstruction[27] ),
    .A2(net1258),
    .B1(net1006),
    .B2(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__mux2_1 _10344_ (.A0(\core.registers[18][27] ),
    .A1(\core.registers[19][27] ),
    .S(net1512),
    .X(_05332_));
 sky130_fd_sc_hd__mux2_1 _10345_ (.A0(\core.registers[16][27] ),
    .A1(\core.registers[17][27] ),
    .S(net1512),
    .X(_05333_));
 sky130_fd_sc_hd__mux2_1 _10346_ (.A0(_05332_),
    .A1(_05333_),
    .S(net1537),
    .X(_05334_));
 sky130_fd_sc_hd__o221a_1 _10347_ (.A1(net1657),
    .A2(\core.registers[23][27] ),
    .B1(net1512),
    .B2(\core.registers[22][27] ),
    .C1(net1556),
    .X(_05335_));
 sky130_fd_sc_hd__mux2_1 _10348_ (.A0(\core.registers[20][27] ),
    .A1(\core.registers[21][27] ),
    .S(net1512),
    .X(_05336_));
 sky130_fd_sc_hd__or2_1 _10349_ (.A(\core.registers[0][27] ),
    .B(net1511),
    .X(_05337_));
 sky130_fd_sc_hd__o211a_1 _10350_ (.A1(\core.registers[1][27] ),
    .A2(net1460),
    .B1(_05337_),
    .C1(net1537),
    .X(_05338_));
 sky130_fd_sc_hd__mux2_1 _10351_ (.A0(\core.registers[2][27] ),
    .A1(\core.registers[3][27] ),
    .S(net1511),
    .X(_05339_));
 sky130_fd_sc_hd__a211o_1 _10352_ (.A1(net1556),
    .A2(_05339_),
    .B1(_05338_),
    .C1(net1589),
    .X(_05340_));
 sky130_fd_sc_hd__mux2_1 _10353_ (.A0(\core.registers[4][27] ),
    .A1(\core.registers[5][27] ),
    .S(net1511),
    .X(_05341_));
 sky130_fd_sc_hd__o221a_1 _10354_ (.A1(net1657),
    .A2(\core.registers[7][27] ),
    .B1(net1511),
    .B2(\core.registers[6][27] ),
    .C1(net1556),
    .X(_05342_));
 sky130_fd_sc_hd__a211o_1 _10355_ (.A1(net1536),
    .A2(_05341_),
    .B1(_05342_),
    .C1(net1580),
    .X(_05343_));
 sky130_fd_sc_hd__a211o_1 _10356_ (.A1(net1536),
    .A2(_05336_),
    .B1(_05335_),
    .C1(net1580),
    .X(_05344_));
 sky130_fd_sc_hd__o211a_1 _10357_ (.A1(net1589),
    .A2(_05334_),
    .B1(_05344_),
    .C1(net1599),
    .X(_05345_));
 sky130_fd_sc_hd__a311o_4 _10358_ (.A1(net1595),
    .A2(_05340_),
    .A3(_05343_),
    .B1(_05345_),
    .C1(net1568),
    .X(_05346_));
 sky130_fd_sc_hd__mux2_1 _10359_ (.A0(\core.registers[28][27] ),
    .A1(\core.registers[29][27] ),
    .S(net1490),
    .X(_05347_));
 sky130_fd_sc_hd__a221o_1 _10360_ (.A1(net1652),
    .A2(\core.registers[30][27] ),
    .B1(\core.registers[31][27] ),
    .B2(net1490),
    .C1(net1666),
    .X(_05348_));
 sky130_fd_sc_hd__mux2_1 _10361_ (.A0(\core.registers[8][27] ),
    .A1(\core.registers[9][27] ),
    .S(net1490),
    .X(_05349_));
 sky130_fd_sc_hd__mux2_1 _10362_ (.A0(\core.registers[10][27] ),
    .A1(\core.registers[11][27] ),
    .S(net1491),
    .X(_05350_));
 sky130_fd_sc_hd__mux2_1 _10363_ (.A0(_05349_),
    .A1(_05350_),
    .S(net1551),
    .X(_05351_));
 sky130_fd_sc_hd__or2_1 _10364_ (.A(\core.registers[25][27] ),
    .B(net1460),
    .X(_05352_));
 sky130_fd_sc_hd__o21a_1 _10365_ (.A1(\core.registers[24][27] ),
    .A2(net1490),
    .B1(net1666),
    .X(_05353_));
 sky130_fd_sc_hd__a22o_1 _10366_ (.A1(net1652),
    .A2(\core.registers[26][27] ),
    .B1(\core.registers[27][27] ),
    .B2(net1490),
    .X(_05354_));
 sky130_fd_sc_hd__a221o_1 _10367_ (.A1(_05352_),
    .A2(_05353_),
    .B1(_05354_),
    .B2(net1791),
    .C1(net1673),
    .X(_05355_));
 sky130_fd_sc_hd__o211a_1 _10368_ (.A1(net1782),
    .A2(_05351_),
    .B1(_05355_),
    .C1(net1670),
    .X(_05356_));
 sky130_fd_sc_hd__mux2_1 _10369_ (.A0(\core.registers[12][27] ),
    .A1(\core.registers[13][27] ),
    .S(net1490),
    .X(_05357_));
 sky130_fd_sc_hd__mux2_1 _10370_ (.A0(\core.registers[14][27] ),
    .A1(\core.registers[15][27] ),
    .S(net1490),
    .X(_05358_));
 sky130_fd_sc_hd__mux2_1 _10371_ (.A0(_05357_),
    .A1(_05358_),
    .S(net1551),
    .X(_05359_));
 sky130_fd_sc_hd__o21a_1 _10372_ (.A1(net1791),
    .A2(_05347_),
    .B1(_05348_),
    .X(_05360_));
 sky130_fd_sc_hd__mux2_1 _10373_ (.A0(_05359_),
    .A1(_05360_),
    .S(net1782),
    .X(_05361_));
 sky130_fd_sc_hd__a21o_1 _10374_ (.A1(net1785),
    .A2(_05361_),
    .B1(net1563),
    .X(_05362_));
 sky130_fd_sc_hd__o21ai_4 _10375_ (.A1(_05356_),
    .A2(_05362_),
    .B1(_05346_),
    .Y(_05363_));
 sky130_fd_sc_hd__o2bb2a_4 _10376_ (.A1_N(net1096),
    .A2_N(net868),
    .B1(_05363_),
    .B2(net1044),
    .X(_05364_));
 sky130_fd_sc_hd__inv_2 _10377_ (.A(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__mux2_8 _10378_ (.A0(net469),
    .A1(_05365_),
    .S(net1251),
    .X(_05366_));
 sky130_fd_sc_hd__nor2_4 _10379_ (.A(_05331_),
    .B(_05366_),
    .Y(_05367_));
 sky130_fd_sc_hd__inv_2 _10380_ (.A(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__and2_4 _10381_ (.A(_05331_),
    .B(_05366_),
    .X(_05369_));
 sky130_fd_sc_hd__a31o_1 _10382_ (.A1(net1618),
    .A2(_04014_),
    .A3(_04136_),
    .B1(net1186),
    .X(_05370_));
 sky130_fd_sc_hd__a21o_1 _10383_ (.A1(\core.pipe1_csrData[26] ),
    .A2(net1250),
    .B1(net1237),
    .X(_05371_));
 sky130_fd_sc_hd__a21o_1 _10384_ (.A1(_05370_),
    .A2(_05371_),
    .B1(net1244),
    .X(_05372_));
 sky130_fd_sc_hd__o21a_4 _10385_ (.A1(\core.pipe1_resultRegister[26] ),
    .A2(net1188),
    .B1(_05372_),
    .X(_05373_));
 sky130_fd_sc_hd__mux2_1 _10386_ (.A0(\core.registers[14][26] ),
    .A1(\core.registers[15][26] ),
    .S(net1363),
    .X(_05374_));
 sky130_fd_sc_hd__mux2_1 _10387_ (.A0(\core.registers[12][26] ),
    .A1(\core.registers[13][26] ),
    .S(net1363),
    .X(_05375_));
 sky130_fd_sc_hd__mux2_1 _10388_ (.A0(_05374_),
    .A1(_05375_),
    .S(net1328),
    .X(_05376_));
 sky130_fd_sc_hd__mux2_1 _10389_ (.A0(\core.registers[28][26] ),
    .A1(\core.registers[29][26] ),
    .S(net1374),
    .X(_05377_));
 sky130_fd_sc_hd__a221o_1 _10390_ (.A1(net1676),
    .A2(\core.registers[30][26] ),
    .B1(\core.registers[31][26] ),
    .B2(net1364),
    .C1(net1699),
    .X(_05378_));
 sky130_fd_sc_hd__o21a_1 _10391_ (.A1(net1769),
    .A2(_05377_),
    .B1(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_1 _10392_ (.A0(\core.registers[8][26] ),
    .A1(\core.registers[9][26] ),
    .S(net1364),
    .X(_05380_));
 sky130_fd_sc_hd__mux2_1 _10393_ (.A0(\core.registers[10][26] ),
    .A1(\core.registers[11][26] ),
    .S(net1363),
    .X(_05381_));
 sky130_fd_sc_hd__mux2_1 _10394_ (.A0(_05380_),
    .A1(_05381_),
    .S(net1341),
    .X(_05382_));
 sky130_fd_sc_hd__mux2_1 _10395_ (.A0(\core.registers[24][26] ),
    .A1(\core.registers[25][26] ),
    .S(net1364),
    .X(_05383_));
 sky130_fd_sc_hd__a22o_1 _10396_ (.A1(net1676),
    .A2(\core.registers[26][26] ),
    .B1(\core.registers[27][26] ),
    .B2(net1364),
    .X(_05384_));
 sky130_fd_sc_hd__mux2_1 _10397_ (.A0(_05383_),
    .A1(_05384_),
    .S(net1769),
    .X(_05385_));
 sky130_fd_sc_hd__mux4_2 _10398_ (.A0(_05376_),
    .A1(_05379_),
    .A2(_05382_),
    .A3(_05385_),
    .S0(net1753),
    .S1(net1704),
    .X(_05386_));
 sky130_fd_sc_hd__nand2_2 _10399_ (.A(net1429),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__mux4_1 _10400_ (.A0(\core.registers[16][26] ),
    .A1(\core.registers[17][26] ),
    .A2(\core.registers[20][26] ),
    .A3(\core.registers[21][26] ),
    .S0(net1423),
    .S1(net1456),
    .X(_05388_));
 sky130_fd_sc_hd__o22a_1 _10401_ (.A1(net1696),
    .A2(\core.registers[23][26] ),
    .B1(net1423),
    .B2(\core.registers[22][26] ),
    .X(_05389_));
 sky130_fd_sc_hd__o22a_1 _10402_ (.A1(net1697),
    .A2(\core.registers[19][26] ),
    .B1(net1423),
    .B2(\core.registers[18][26] ),
    .X(_05390_));
 sky130_fd_sc_hd__mux2_1 _10403_ (.A0(_05389_),
    .A1(_05390_),
    .S(net1444),
    .X(_05391_));
 sky130_fd_sc_hd__o21a_1 _10404_ (.A1(net1337),
    .A2(_05391_),
    .B1(net1326),
    .X(_05392_));
 sky130_fd_sc_hd__o21a_1 _10405_ (.A1(net1353),
    .A2(_05388_),
    .B1(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__o22a_1 _10406_ (.A1(net1697),
    .A2(\core.registers[7][26] ),
    .B1(net1425),
    .B2(\core.registers[6][26] ),
    .X(_05394_));
 sky130_fd_sc_hd__o22a_1 _10407_ (.A1(net1697),
    .A2(\core.registers[3][26] ),
    .B1(net1425),
    .B2(\core.registers[2][26] ),
    .X(_05395_));
 sky130_fd_sc_hd__mux2_1 _10408_ (.A0(_05394_),
    .A1(_05395_),
    .S(net1445),
    .X(_05396_));
 sky130_fd_sc_hd__or2_2 _10409_ (.A(net1338),
    .B(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__mux4_1 _10410_ (.A0(\core.registers[0][26] ),
    .A1(\core.registers[1][26] ),
    .A2(\core.registers[4][26] ),
    .A3(\core.registers[5][26] ),
    .S0(net1425),
    .S1(net1456),
    .X(_05398_));
 sky130_fd_sc_hd__o21a_1 _10411_ (.A1(net1353),
    .A2(_05398_),
    .B1(net1322),
    .X(_05399_));
 sky130_fd_sc_hd__a21oi_4 _10412_ (.A1(_05397_),
    .A2(_05399_),
    .B1(_05393_),
    .Y(_05400_));
 sky130_fd_sc_hd__o211ai_4 _10413_ (.A1(net1429),
    .A2(_05400_),
    .B1(_05387_),
    .C1(net1142),
    .Y(_05401_));
 sky130_fd_sc_hd__o211ai_4 _10414_ (.A1(net1142),
    .A2(net1004),
    .B1(_05401_),
    .C1(net1240),
    .Y(_05402_));
 sky130_fd_sc_hd__nor2_1 _10415_ (.A(net1041),
    .B(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__o22a_4 _10416_ (.A1(\core.pipe0_currentInstruction[26] ),
    .A2(net1257),
    .B1(net1006),
    .B2(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__mux2_1 _10417_ (.A0(\core.registers[18][26] ),
    .A1(\core.registers[19][26] ),
    .S(net1523),
    .X(_05405_));
 sky130_fd_sc_hd__mux2_1 _10418_ (.A0(\core.registers[16][26] ),
    .A1(\core.registers[17][26] ),
    .S(net1523),
    .X(_05406_));
 sky130_fd_sc_hd__mux2_1 _10419_ (.A0(_05405_),
    .A1(_05406_),
    .S(net1539),
    .X(_05407_));
 sky130_fd_sc_hd__o221a_1 _10420_ (.A1(net1659),
    .A2(\core.registers[23][26] ),
    .B1(net1521),
    .B2(\core.registers[22][26] ),
    .C1(net1558),
    .X(_05408_));
 sky130_fd_sc_hd__mux2_1 _10421_ (.A0(\core.registers[20][26] ),
    .A1(\core.registers[21][26] ),
    .S(net1521),
    .X(_05409_));
 sky130_fd_sc_hd__or2_1 _10422_ (.A(\core.registers[0][26] ),
    .B(net1521),
    .X(_05410_));
 sky130_fd_sc_hd__o211a_1 _10423_ (.A1(\core.registers[1][26] ),
    .A2(net1460),
    .B1(_05410_),
    .C1(net1539),
    .X(_05411_));
 sky130_fd_sc_hd__mux2_1 _10424_ (.A0(\core.registers[2][26] ),
    .A1(\core.registers[3][26] ),
    .S(net1521),
    .X(_05412_));
 sky130_fd_sc_hd__a211o_1 _10425_ (.A1(net1558),
    .A2(_05412_),
    .B1(_05411_),
    .C1(net1591),
    .X(_05413_));
 sky130_fd_sc_hd__mux2_1 _10426_ (.A0(\core.registers[4][26] ),
    .A1(\core.registers[5][26] ),
    .S(net1523),
    .X(_05414_));
 sky130_fd_sc_hd__o221a_1 _10427_ (.A1(net1660),
    .A2(\core.registers[7][26] ),
    .B1(net1521),
    .B2(\core.registers[6][26] ),
    .C1(net1558),
    .X(_05415_));
 sky130_fd_sc_hd__a211o_1 _10428_ (.A1(net1538),
    .A2(_05414_),
    .B1(_05415_),
    .C1(net1579),
    .X(_05416_));
 sky130_fd_sc_hd__a211o_1 _10429_ (.A1(net1539),
    .A2(_05409_),
    .B1(_05408_),
    .C1(net1579),
    .X(_05417_));
 sky130_fd_sc_hd__o211a_1 _10430_ (.A1(net1590),
    .A2(_05407_),
    .B1(_05417_),
    .C1(net1599),
    .X(_05418_));
 sky130_fd_sc_hd__a31o_4 _10431_ (.A1(net1596),
    .A2(_05413_),
    .A3(_05416_),
    .B1(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__mux2_1 _10432_ (.A0(\core.registers[28][26] ),
    .A1(\core.registers[29][26] ),
    .S(net1472),
    .X(_05420_));
 sky130_fd_sc_hd__a221o_1 _10433_ (.A1(net1642),
    .A2(\core.registers[30][26] ),
    .B1(\core.registers[31][26] ),
    .B2(net1463),
    .C1(net1663),
    .X(_05421_));
 sky130_fd_sc_hd__mux2_1 _10434_ (.A0(\core.registers[8][26] ),
    .A1(\core.registers[9][26] ),
    .S(net1462),
    .X(_05422_));
 sky130_fd_sc_hd__mux2_1 _10435_ (.A0(\core.registers[10][26] ),
    .A1(\core.registers[11][26] ),
    .S(net1462),
    .X(_05423_));
 sky130_fd_sc_hd__mux2_1 _10436_ (.A0(_05422_),
    .A1(_05423_),
    .S(net1543),
    .X(_05424_));
 sky130_fd_sc_hd__mux2_1 _10437_ (.A0(\core.registers[24][26] ),
    .A1(\core.registers[25][26] ),
    .S(net1462),
    .X(_05425_));
 sky130_fd_sc_hd__a22o_1 _10438_ (.A1(net1642),
    .A2(\core.registers[26][26] ),
    .B1(\core.registers[27][26] ),
    .B2(net1463),
    .X(_05426_));
 sky130_fd_sc_hd__mux2_1 _10439_ (.A0(_05425_),
    .A1(_05426_),
    .S(net1787),
    .X(_05427_));
 sky130_fd_sc_hd__mux2_1 _10440_ (.A0(_05424_),
    .A1(_05427_),
    .S(net1778),
    .X(_05428_));
 sky130_fd_sc_hd__mux2_1 _10441_ (.A0(\core.registers[12][26] ),
    .A1(\core.registers[13][26] ),
    .S(net1470),
    .X(_05429_));
 sky130_fd_sc_hd__mux2_1 _10442_ (.A0(\core.registers[14][26] ),
    .A1(\core.registers[15][26] ),
    .S(net1470),
    .X(_05430_));
 sky130_fd_sc_hd__mux2_1 _10443_ (.A0(_05429_),
    .A1(_05430_),
    .S(net1544),
    .X(_05431_));
 sky130_fd_sc_hd__nor2_1 _10444_ (.A(net1778),
    .B(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__o21ai_1 _10445_ (.A1(net1787),
    .A2(_05420_),
    .B1(_05421_),
    .Y(_05433_));
 sky130_fd_sc_hd__a211o_1 _10446_ (.A1(net1778),
    .A2(_05433_),
    .B1(_05432_),
    .C1(net1668),
    .X(_05434_));
 sky130_fd_sc_hd__a21oi_2 _10447_ (.A1(net1668),
    .A2(_05428_),
    .B1(net1562),
    .Y(_05435_));
 sky130_fd_sc_hd__a2bb2o_1 _10448_ (.A1_N(net1567),
    .A2_N(_05419_),
    .B1(_05434_),
    .B2(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__o2bb2a_2 _10449_ (.A1_N(net1094),
    .A2_N(net1004),
    .B1(_05436_),
    .B2(net1045),
    .X(_05437_));
 sky130_fd_sc_hd__inv_2 _10450_ (.A(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hd__mux2_4 _10451_ (.A0(net468),
    .A1(_05438_),
    .S(net1251),
    .X(_05439_));
 sky130_fd_sc_hd__and2_2 _10452_ (.A(_05404_),
    .B(_05439_),
    .X(_05440_));
 sky130_fd_sc_hd__nor2_1 _10453_ (.A(_05404_),
    .B(_05439_),
    .Y(_05441_));
 sky130_fd_sc_hd__or2_4 _10454_ (.A(_05440_),
    .B(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__clkinv_4 _10455_ (.A(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__a31o_1 _10456_ (.A1(net1617),
    .A2(_04014_),
    .A3(_04222_),
    .B1(net1187),
    .X(_05444_));
 sky130_fd_sc_hd__a21o_1 _10457_ (.A1(\core.pipe1_csrData[25] ),
    .A2(net1249),
    .B1(net1237),
    .X(_05445_));
 sky130_fd_sc_hd__a21o_1 _10458_ (.A1(_05444_),
    .A2(_05445_),
    .B1(net1244),
    .X(_05446_));
 sky130_fd_sc_hd__o21a_4 _10459_ (.A1(\core.pipe1_resultRegister[25] ),
    .A2(net1188),
    .B1(_05446_),
    .X(_05447_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(\core.registers[14][25] ),
    .A1(\core.registers[15][25] ),
    .S(net1373),
    .X(_05448_));
 sky130_fd_sc_hd__mux2_1 _10461_ (.A0(\core.registers[12][25] ),
    .A1(\core.registers[13][25] ),
    .S(net1373),
    .X(_05449_));
 sky130_fd_sc_hd__mux2_1 _10462_ (.A0(_05448_),
    .A1(_05449_),
    .S(net1329),
    .X(_05450_));
 sky130_fd_sc_hd__mux2_1 _10463_ (.A0(\core.registers[28][25] ),
    .A1(\core.registers[29][25] ),
    .S(net1374),
    .X(_05451_));
 sky130_fd_sc_hd__a221o_1 _10464_ (.A1(net1685),
    .A2(\core.registers[30][25] ),
    .B1(\core.registers[31][25] ),
    .B2(net1373),
    .C1(net1700),
    .X(_05452_));
 sky130_fd_sc_hd__o21a_1 _10465_ (.A1(net1771),
    .A2(_05451_),
    .B1(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__mux2_1 _10466_ (.A0(\core.registers[8][25] ),
    .A1(\core.registers[9][25] ),
    .S(net1374),
    .X(_05454_));
 sky130_fd_sc_hd__mux2_1 _10467_ (.A0(\core.registers[10][25] ),
    .A1(\core.registers[11][25] ),
    .S(net1374),
    .X(_05455_));
 sky130_fd_sc_hd__mux2_1 _10468_ (.A0(_05454_),
    .A1(_05455_),
    .S(net1343),
    .X(_05456_));
 sky130_fd_sc_hd__mux2_1 _10469_ (.A0(\core.registers[24][25] ),
    .A1(\core.registers[25][25] ),
    .S(net1373),
    .X(_05457_));
 sky130_fd_sc_hd__a22o_1 _10470_ (.A1(net1685),
    .A2(\core.registers[26][25] ),
    .B1(\core.registers[27][25] ),
    .B2(net1372),
    .X(_05458_));
 sky130_fd_sc_hd__mux2_1 _10471_ (.A0(_05457_),
    .A1(_05458_),
    .S(net1771),
    .X(_05459_));
 sky130_fd_sc_hd__mux4_2 _10472_ (.A0(_05450_),
    .A1(_05453_),
    .A2(_05456_),
    .A3(_05459_),
    .S0(net1754),
    .S1(net1704),
    .X(_05460_));
 sky130_fd_sc_hd__nand2_1 _10473_ (.A(net1430),
    .B(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__mux4_1 _10474_ (.A0(\core.registers[16][25] ),
    .A1(\core.registers[17][25] ),
    .A2(\core.registers[20][25] ),
    .A3(\core.registers[21][25] ),
    .S0(net1389),
    .S1(net1449),
    .X(_05462_));
 sky130_fd_sc_hd__o22a_1 _10475_ (.A1(net1677),
    .A2(\core.registers[23][25] ),
    .B1(net1389),
    .B2(\core.registers[22][25] ),
    .X(_05463_));
 sky130_fd_sc_hd__o22a_1 _10476_ (.A1(net1677),
    .A2(\core.registers[19][25] ),
    .B1(net1389),
    .B2(\core.registers[18][25] ),
    .X(_05464_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(_05463_),
    .A1(_05464_),
    .S(net1437),
    .X(_05465_));
 sky130_fd_sc_hd__o21a_1 _10478_ (.A1(net1331),
    .A2(_05465_),
    .B1(net1324),
    .X(_05466_));
 sky130_fd_sc_hd__o21a_1 _10479_ (.A1(net1346),
    .A2(_05462_),
    .B1(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__o22a_1 _10480_ (.A1(net1681),
    .A2(\core.registers[7][25] ),
    .B1(net1389),
    .B2(\core.registers[6][25] ),
    .X(_05468_));
 sky130_fd_sc_hd__o22a_1 _10481_ (.A1(net1681),
    .A2(\core.registers[3][25] ),
    .B1(net1389),
    .B2(\core.registers[2][25] ),
    .X(_05469_));
 sky130_fd_sc_hd__mux2_1 _10482_ (.A0(_05468_),
    .A1(_05469_),
    .S(net1437),
    .X(_05470_));
 sky130_fd_sc_hd__or2_2 _10483_ (.A(net1331),
    .B(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__mux4_1 _10484_ (.A0(\core.registers[0][25] ),
    .A1(\core.registers[1][25] ),
    .A2(\core.registers[4][25] ),
    .A3(\core.registers[5][25] ),
    .S0(net1389),
    .S1(net1449),
    .X(_05472_));
 sky130_fd_sc_hd__o21a_1 _10485_ (.A1(net1356),
    .A2(_05472_),
    .B1(net1321),
    .X(_05473_));
 sky130_fd_sc_hd__a21oi_4 _10486_ (.A1(_05471_),
    .A2(_05473_),
    .B1(_05467_),
    .Y(_05474_));
 sky130_fd_sc_hd__o211ai_4 _10487_ (.A1(net1430),
    .A2(_05474_),
    .B1(_05461_),
    .C1(net1141),
    .Y(_05475_));
 sky130_fd_sc_hd__o211ai_4 _10488_ (.A1(net1141),
    .A2(net999),
    .B1(_05475_),
    .C1(net1239),
    .Y(_05476_));
 sky130_fd_sc_hd__nor2_1 _10489_ (.A(net1039),
    .B(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__o22a_4 _10490_ (.A1(\core.pipe0_currentInstruction[25] ),
    .A2(net1252),
    .B1(net1005),
    .B2(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__mux2_1 _10491_ (.A0(\core.registers[18][25] ),
    .A1(\core.registers[19][25] ),
    .S(net1486),
    .X(_05479_));
 sky130_fd_sc_hd__mux2_1 _10492_ (.A0(\core.registers[16][25] ),
    .A1(\core.registers[17][25] ),
    .S(net1486),
    .X(_05480_));
 sky130_fd_sc_hd__mux2_1 _10493_ (.A0(_05479_),
    .A1(_05480_),
    .S(net1529),
    .X(_05481_));
 sky130_fd_sc_hd__o221a_1 _10494_ (.A1(net1646),
    .A2(\core.registers[23][25] ),
    .B1(net1486),
    .B2(\core.registers[22][25] ),
    .C1(net1549),
    .X(_05482_));
 sky130_fd_sc_hd__mux2_1 _10495_ (.A0(\core.registers[20][25] ),
    .A1(\core.registers[21][25] ),
    .S(net1486),
    .X(_05483_));
 sky130_fd_sc_hd__or2_1 _10496_ (.A(\core.registers[0][25] ),
    .B(net1489),
    .X(_05484_));
 sky130_fd_sc_hd__o211a_1 _10497_ (.A1(\core.registers[1][25] ),
    .A2(net1459),
    .B1(_05484_),
    .C1(net1532),
    .X(_05485_));
 sky130_fd_sc_hd__mux2_1 _10498_ (.A0(\core.registers[2][25] ),
    .A1(\core.registers[3][25] ),
    .S(net1486),
    .X(_05486_));
 sky130_fd_sc_hd__a211o_1 _10499_ (.A1(net1549),
    .A2(_05486_),
    .B1(_05485_),
    .C1(net1586),
    .X(_05487_));
 sky130_fd_sc_hd__mux2_1 _10500_ (.A0(\core.registers[4][25] ),
    .A1(\core.registers[5][25] ),
    .S(net1486),
    .X(_05488_));
 sky130_fd_sc_hd__o221a_1 _10501_ (.A1(net1650),
    .A2(\core.registers[7][25] ),
    .B1(net1486),
    .B2(\core.registers[6][25] ),
    .C1(net1549),
    .X(_05489_));
 sky130_fd_sc_hd__a211o_1 _10502_ (.A1(net1529),
    .A2(_05488_),
    .B1(_05489_),
    .C1(net1573),
    .X(_05490_));
 sky130_fd_sc_hd__a211o_1 _10503_ (.A1(net1529),
    .A2(_05483_),
    .B1(_05482_),
    .C1(net1573),
    .X(_05491_));
 sky130_fd_sc_hd__o211a_1 _10504_ (.A1(net1584),
    .A2(_05481_),
    .B1(_05491_),
    .C1(net1597),
    .X(_05492_));
 sky130_fd_sc_hd__a31o_2 _10505_ (.A1(net1593),
    .A2(_05487_),
    .A3(_05490_),
    .B1(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__mux2_1 _10506_ (.A0(\core.registers[8][25] ),
    .A1(\core.registers[9][25] ),
    .S(net1475),
    .X(_05494_));
 sky130_fd_sc_hd__mux2_1 _10507_ (.A0(\core.registers[10][25] ),
    .A1(\core.registers[11][25] ),
    .S(net1475),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _10508_ (.A0(\core.registers[28][25] ),
    .A1(\core.registers[29][25] ),
    .S(net1472),
    .X(_05496_));
 sky130_fd_sc_hd__a221o_1 _10509_ (.A1(net1645),
    .A2(\core.registers[30][25] ),
    .B1(\core.registers[31][25] ),
    .B2(net1472),
    .C1(net1663),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _10510_ (.A0(_05494_),
    .A1(_05495_),
    .S(net1544),
    .X(_05498_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(\core.registers[24][25] ),
    .A1(\core.registers[25][25] ),
    .S(net1475),
    .X(_05499_));
 sky130_fd_sc_hd__a22o_1 _10512_ (.A1(net1645),
    .A2(\core.registers[26][25] ),
    .B1(\core.registers[27][25] ),
    .B2(net1471),
    .X(_05500_));
 sky130_fd_sc_hd__mux2_1 _10513_ (.A0(_05499_),
    .A1(_05500_),
    .S(net1789),
    .X(_05501_));
 sky130_fd_sc_hd__mux2_1 _10514_ (.A0(_05498_),
    .A1(_05501_),
    .S(net1780),
    .X(_05502_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(\core.registers[12][25] ),
    .A1(\core.registers[13][25] ),
    .S(net1471),
    .X(_05503_));
 sky130_fd_sc_hd__mux2_1 _10516_ (.A0(\core.registers[14][25] ),
    .A1(\core.registers[15][25] ),
    .S(net1471),
    .X(_05504_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(_05503_),
    .A1(_05504_),
    .S(net1544),
    .X(_05505_));
 sky130_fd_sc_hd__nor2_1 _10518_ (.A(net1780),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__o21ai_1 _10519_ (.A1(net1789),
    .A2(_05496_),
    .B1(_05497_),
    .Y(_05507_));
 sky130_fd_sc_hd__a211o_1 _10520_ (.A1(net1780),
    .A2(_05507_),
    .B1(_05506_),
    .C1(net1668),
    .X(_05508_));
 sky130_fd_sc_hd__a21oi_1 _10521_ (.A1(net1668),
    .A2(_05502_),
    .B1(net1562),
    .Y(_05509_));
 sky130_fd_sc_hd__a2bb2o_1 _10522_ (.A1_N(net1567),
    .A2_N(_05493_),
    .B1(_05508_),
    .B2(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__o2bb2a_2 _10523_ (.A1_N(net1094),
    .A2_N(net997),
    .B1(_05510_),
    .B2(net1045),
    .X(_05511_));
 sky130_fd_sc_hd__inv_2 _10524_ (.A(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__mux2_4 _10525_ (.A0(net467),
    .A1(_05512_),
    .S(net1251),
    .X(_05513_));
 sky130_fd_sc_hd__nor2_2 _10526_ (.A(_05478_),
    .B(_05513_),
    .Y(_05514_));
 sky130_fd_sc_hd__and2_2 _10527_ (.A(_05478_),
    .B(_05513_),
    .X(_05515_));
 sky130_fd_sc_hd__a31o_1 _10528_ (.A1(net1617),
    .A2(_04014_),
    .A3(_04310_),
    .B1(net1186),
    .X(_05516_));
 sky130_fd_sc_hd__a21o_1 _10529_ (.A1(\core.pipe1_csrData[24] ),
    .A2(net1249),
    .B1(net1238),
    .X(_05517_));
 sky130_fd_sc_hd__a21o_1 _10530_ (.A1(_05516_),
    .A2(_05517_),
    .B1(net1244),
    .X(_05518_));
 sky130_fd_sc_hd__o21a_4 _10531_ (.A1(\core.pipe1_resultRegister[24] ),
    .A2(net1188),
    .B1(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__nor2_1 _10532_ (.A(net1141),
    .B(net995),
    .Y(_05520_));
 sky130_fd_sc_hd__mux2_1 _10533_ (.A0(\core.registers[12][24] ),
    .A1(\core.registers[13][24] ),
    .S(net1373),
    .X(_05521_));
 sky130_fd_sc_hd__mux2_1 _10534_ (.A0(\core.registers[14][24] ),
    .A1(\core.registers[15][24] ),
    .S(net1372),
    .X(_05522_));
 sky130_fd_sc_hd__mux2_1 _10535_ (.A0(_05521_),
    .A1(_05522_),
    .S(net1343),
    .X(_05523_));
 sky130_fd_sc_hd__nor2_1 _10536_ (.A(net1755),
    .B(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__a221o_1 _10537_ (.A1(net1676),
    .A2(\core.registers[30][24] ),
    .B1(\core.registers[31][24] ),
    .B2(net1375),
    .C1(net1699),
    .X(_05525_));
 sky130_fd_sc_hd__mux2_1 _10538_ (.A0(\core.registers[28][24] ),
    .A1(\core.registers[29][24] ),
    .S(net1373),
    .X(_05526_));
 sky130_fd_sc_hd__o21ai_1 _10539_ (.A1(net1769),
    .A2(_05526_),
    .B1(_05525_),
    .Y(_05527_));
 sky130_fd_sc_hd__a211o_1 _10540_ (.A1(net1754),
    .A2(_05527_),
    .B1(_05524_),
    .C1(net1705),
    .X(_05528_));
 sky130_fd_sc_hd__mux2_1 _10541_ (.A0(\core.registers[8][24] ),
    .A1(\core.registers[9][24] ),
    .S(net1372),
    .X(_05529_));
 sky130_fd_sc_hd__mux2_1 _10542_ (.A0(\core.registers[10][24] ),
    .A1(\core.registers[11][24] ),
    .S(net1372),
    .X(_05530_));
 sky130_fd_sc_hd__mux2_4 _10543_ (.A0(_05529_),
    .A1(_05530_),
    .S(net1343),
    .X(_05531_));
 sky130_fd_sc_hd__or2_1 _10544_ (.A(\core.registers[24][24] ),
    .B(net1373),
    .X(_05532_));
 sky130_fd_sc_hd__o211a_1 _10545_ (.A1(\core.registers[25][24] ),
    .A2(net1358),
    .B1(_05532_),
    .C1(net1700),
    .X(_05533_));
 sky130_fd_sc_hd__and3_1 _10546_ (.A(net1769),
    .B(\core.registers[27][24] ),
    .C(net1373),
    .X(_05534_));
 sky130_fd_sc_hd__a211o_1 _10547_ (.A1(\core.registers[26][24] ),
    .A2(net1319),
    .B1(_05534_),
    .C1(net1708),
    .X(_05535_));
 sky130_fd_sc_hd__o221ai_4 _10548_ (.A1(net1754),
    .A2(_05531_),
    .B1(_05533_),
    .B2(_05535_),
    .C1(net1704),
    .Y(_05536_));
 sky130_fd_sc_hd__mux4_1 _10549_ (.A0(\core.registers[16][24] ),
    .A1(\core.registers[17][24] ),
    .A2(\core.registers[20][24] ),
    .A3(\core.registers[21][24] ),
    .S0(net1375),
    .S1(net1448),
    .X(_05537_));
 sky130_fd_sc_hd__o22a_1 _10550_ (.A1(net1676),
    .A2(\core.registers[23][24] ),
    .B1(net1375),
    .B2(\core.registers[22][24] ),
    .X(_05538_));
 sky130_fd_sc_hd__o22a_1 _10551_ (.A1(net1676),
    .A2(\core.registers[19][24] ),
    .B1(net1375),
    .B2(\core.registers[18][24] ),
    .X(_05539_));
 sky130_fd_sc_hd__mux2_1 _10552_ (.A0(_05538_),
    .A1(_05539_),
    .S(net1434),
    .X(_05540_));
 sky130_fd_sc_hd__o21a_1 _10553_ (.A1(net1329),
    .A2(_05540_),
    .B1(net1324),
    .X(_05541_));
 sky130_fd_sc_hd__o21ai_1 _10554_ (.A1(net1343),
    .A2(_05537_),
    .B1(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__o22a_1 _10555_ (.A1(net1677),
    .A2(\core.registers[7][24] ),
    .B1(net1376),
    .B2(\core.registers[6][24] ),
    .X(_05543_));
 sky130_fd_sc_hd__o22a_1 _10556_ (.A1(net1677),
    .A2(\core.registers[3][24] ),
    .B1(net1375),
    .B2(\core.registers[2][24] ),
    .X(_05544_));
 sky130_fd_sc_hd__mux2_1 _10557_ (.A0(_05543_),
    .A1(_05544_),
    .S(net1436),
    .X(_05545_));
 sky130_fd_sc_hd__or2_1 _10558_ (.A(net1329),
    .B(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__mux4_1 _10559_ (.A0(\core.registers[0][24] ),
    .A1(\core.registers[1][24] ),
    .A2(\core.registers[4][24] ),
    .A3(\core.registers[5][24] ),
    .S0(net1375),
    .S1(net1448),
    .X(_05547_));
 sky130_fd_sc_hd__o21a_1 _10560_ (.A1(net1343),
    .A2(_05547_),
    .B1(net1320),
    .X(_05548_));
 sky130_fd_sc_hd__a21oi_1 _10561_ (.A1(_05546_),
    .A2(_05548_),
    .B1(net1429),
    .Y(_05549_));
 sky130_fd_sc_hd__a32o_1 _10562_ (.A1(net1430),
    .A2(_05528_),
    .A3(_05536_),
    .B1(_05542_),
    .B2(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__a211o_1 _10563_ (.A1(net1141),
    .A2(_05550_),
    .B1(_05520_),
    .C1(_04095_),
    .X(_05551_));
 sky130_fd_sc_hd__nor2_1 _10564_ (.A(net1039),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__o22a_4 _10565_ (.A1(net1754),
    .A2(net1252),
    .B1(net1005),
    .B2(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__mux2_1 _10566_ (.A0(\core.registers[18][24] ),
    .A1(\core.registers[19][24] ),
    .S(net1473),
    .X(_05554_));
 sky130_fd_sc_hd__mux2_1 _10567_ (.A0(\core.registers[16][24] ),
    .A1(\core.registers[17][24] ),
    .S(net1473),
    .X(_05555_));
 sky130_fd_sc_hd__mux2_1 _10568_ (.A0(_05554_),
    .A1(_05555_),
    .S(net1529),
    .X(_05556_));
 sky130_fd_sc_hd__o221a_1 _10569_ (.A1(net1645),
    .A2(\core.registers[23][24] ),
    .B1(net1473),
    .B2(\core.registers[22][24] ),
    .C1(net1544),
    .X(_05557_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(\core.registers[20][24] ),
    .A1(\core.registers[21][24] ),
    .S(net1473),
    .X(_05558_));
 sky130_fd_sc_hd__or2_1 _10571_ (.A(\core.registers[0][24] ),
    .B(net1473),
    .X(_05559_));
 sky130_fd_sc_hd__o211a_1 _10572_ (.A1(\core.registers[1][24] ),
    .A2(net1459),
    .B1(_05559_),
    .C1(net1529),
    .X(_05560_));
 sky130_fd_sc_hd__mux2_1 _10573_ (.A0(\core.registers[2][24] ),
    .A1(\core.registers[3][24] ),
    .S(net1474),
    .X(_05561_));
 sky130_fd_sc_hd__a211o_1 _10574_ (.A1(net1545),
    .A2(_05561_),
    .B1(_05560_),
    .C1(net1584),
    .X(_05562_));
 sky130_fd_sc_hd__mux2_1 _10575_ (.A0(\core.registers[4][24] ),
    .A1(\core.registers[5][24] ),
    .S(net1474),
    .X(_05563_));
 sky130_fd_sc_hd__o221a_1 _10576_ (.A1(net1645),
    .A2(\core.registers[7][24] ),
    .B1(net1474),
    .B2(\core.registers[6][24] ),
    .C1(net1545),
    .X(_05564_));
 sky130_fd_sc_hd__a211o_1 _10577_ (.A1(net1527),
    .A2(_05563_),
    .B1(_05564_),
    .C1(net1573),
    .X(_05565_));
 sky130_fd_sc_hd__a211o_1 _10578_ (.A1(net1527),
    .A2(_05558_),
    .B1(_05557_),
    .C1(net1573),
    .X(_05566_));
 sky130_fd_sc_hd__o211a_1 _10579_ (.A1(net1584),
    .A2(_05556_),
    .B1(_05566_),
    .C1(net1597),
    .X(_05567_));
 sky130_fd_sc_hd__a31o_1 _10580_ (.A1(net1593),
    .A2(_05562_),
    .A3(_05565_),
    .B1(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__mux2_1 _10581_ (.A0(\core.registers[8][24] ),
    .A1(\core.registers[9][24] ),
    .S(net1471),
    .X(_05569_));
 sky130_fd_sc_hd__mux2_1 _10582_ (.A0(\core.registers[10][24] ),
    .A1(\core.registers[11][24] ),
    .S(net1471),
    .X(_05570_));
 sky130_fd_sc_hd__mux2_1 _10583_ (.A0(\core.registers[28][24] ),
    .A1(\core.registers[29][24] ),
    .S(net1472),
    .X(_05571_));
 sky130_fd_sc_hd__a221o_1 _10584_ (.A1(net1645),
    .A2(\core.registers[30][24] ),
    .B1(\core.registers[31][24] ),
    .B2(net1473),
    .C1(net1663),
    .X(_05572_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(_05569_),
    .A1(_05570_),
    .S(net1544),
    .X(_05573_));
 sky130_fd_sc_hd__mux2_1 _10586_ (.A0(\core.registers[24][24] ),
    .A1(\core.registers[25][24] ),
    .S(net1472),
    .X(_05574_));
 sky130_fd_sc_hd__a22o_1 _10587_ (.A1(net1645),
    .A2(\core.registers[26][24] ),
    .B1(\core.registers[27][24] ),
    .B2(net1472),
    .X(_05575_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(_05574_),
    .A1(_05575_),
    .S(net1787),
    .X(_05576_));
 sky130_fd_sc_hd__mux2_1 _10589_ (.A0(_05573_),
    .A1(_05576_),
    .S(net1779),
    .X(_05577_));
 sky130_fd_sc_hd__o21ai_1 _10590_ (.A1(net1787),
    .A2(_05571_),
    .B1(_05572_),
    .Y(_05578_));
 sky130_fd_sc_hd__mux2_1 _10591_ (.A0(\core.registers[12][24] ),
    .A1(\core.registers[13][24] ),
    .S(net1470),
    .X(_05579_));
 sky130_fd_sc_hd__mux2_1 _10592_ (.A0(\core.registers[14][24] ),
    .A1(\core.registers[15][24] ),
    .S(net1470),
    .X(_05580_));
 sky130_fd_sc_hd__mux2_1 _10593_ (.A0(_05579_),
    .A1(_05580_),
    .S(net1544),
    .X(_05581_));
 sky130_fd_sc_hd__nor2_1 _10594_ (.A(net1778),
    .B(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__a211o_1 _10595_ (.A1(net1779),
    .A2(_05578_),
    .B1(_05582_),
    .C1(net1668),
    .X(_05583_));
 sky130_fd_sc_hd__a21oi_1 _10596_ (.A1(net1668),
    .A2(_05577_),
    .B1(net1561),
    .Y(_05584_));
 sky130_fd_sc_hd__a2bb2o_1 _10597_ (.A1_N(net1567),
    .A2_N(_05568_),
    .B1(_05583_),
    .B2(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__o2bb2a_2 _10598_ (.A1_N(net1094),
    .A2_N(net993),
    .B1(_05585_),
    .B2(net1045),
    .X(_05586_));
 sky130_fd_sc_hd__inv_2 _10599_ (.A(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__mux2_4 _10600_ (.A0(net466),
    .A1(_05587_),
    .S(net1251),
    .X(_05588_));
 sky130_fd_sc_hd__and2_4 _10601_ (.A(_05553_),
    .B(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__nor2_4 _10602_ (.A(_05553_),
    .B(_05588_),
    .Y(_05590_));
 sky130_fd_sc_hd__nor2_8 _10603_ (.A(_05589_),
    .B(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__inv_2 _10604_ (.A(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__a21o_1 _10605_ (.A1(_03997_),
    .A2(net1243),
    .B1(_04022_),
    .X(_05593_));
 sky130_fd_sc_hd__a21o_1 _10606_ (.A1(net1617),
    .A2(_05593_),
    .B1(net1186),
    .X(_05594_));
 sky130_fd_sc_hd__a21o_1 _10607_ (.A1(\core.pipe1_csrData[23] ),
    .A2(net1248),
    .B1(net1238),
    .X(_05595_));
 sky130_fd_sc_hd__a21o_1 _10608_ (.A1(_05594_),
    .A2(_05595_),
    .B1(net1246),
    .X(_05596_));
 sky130_fd_sc_hd__o21a_4 _10609_ (.A1(\core.pipe1_resultRegister[23] ),
    .A2(net1189),
    .B1(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__mux2_1 _10610_ (.A0(\core.registers[14][23] ),
    .A1(\core.registers[15][23] ),
    .S(net1372),
    .X(_05598_));
 sky130_fd_sc_hd__mux2_1 _10611_ (.A0(\core.registers[12][23] ),
    .A1(\core.registers[13][23] ),
    .S(net1372),
    .X(_05599_));
 sky130_fd_sc_hd__mux2_1 _10612_ (.A0(_05598_),
    .A1(_05599_),
    .S(net1329),
    .X(_05600_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(\core.registers[28][23] ),
    .A1(\core.registers[29][23] ),
    .S(net1373),
    .X(_05601_));
 sky130_fd_sc_hd__a221o_1 _10614_ (.A1(net1679),
    .A2(\core.registers[30][23] ),
    .B1(\core.registers[31][23] ),
    .B2(net1374),
    .C1(net1699),
    .X(_05602_));
 sky130_fd_sc_hd__o21a_1 _10615_ (.A1(net1769),
    .A2(_05601_),
    .B1(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__mux2_1 _10616_ (.A0(\core.registers[8][23] ),
    .A1(\core.registers[9][23] ),
    .S(net1372),
    .X(_05604_));
 sky130_fd_sc_hd__mux2_1 _10617_ (.A0(\core.registers[10][23] ),
    .A1(\core.registers[11][23] ),
    .S(net1372),
    .X(_05605_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(_05604_),
    .A1(_05605_),
    .S(net1343),
    .X(_05606_));
 sky130_fd_sc_hd__mux2_1 _10619_ (.A0(\core.registers[24][23] ),
    .A1(\core.registers[25][23] ),
    .S(net1372),
    .X(_05607_));
 sky130_fd_sc_hd__a22o_1 _10620_ (.A1(net1679),
    .A2(\core.registers[26][23] ),
    .B1(\core.registers[27][23] ),
    .B2(net1372),
    .X(_05608_));
 sky130_fd_sc_hd__mux2_1 _10621_ (.A0(_05607_),
    .A1(_05608_),
    .S(net1769),
    .X(_05609_));
 sky130_fd_sc_hd__mux4_2 _10622_ (.A0(_05600_),
    .A1(_05603_),
    .A2(_05606_),
    .A3(_05609_),
    .S0(net1753),
    .S1(net1704),
    .X(_05610_));
 sky130_fd_sc_hd__nand2_1 _10623_ (.A(net1430),
    .B(_05610_),
    .Y(_05611_));
 sky130_fd_sc_hd__mux4_1 _10624_ (.A0(\core.registers[16][23] ),
    .A1(\core.registers[17][23] ),
    .A2(\core.registers[20][23] ),
    .A3(\core.registers[21][23] ),
    .S0(net1375),
    .S1(net1449),
    .X(_05612_));
 sky130_fd_sc_hd__o22a_1 _10625_ (.A1(net1685),
    .A2(\core.registers[23][23] ),
    .B1(net1375),
    .B2(\core.registers[22][23] ),
    .X(_05613_));
 sky130_fd_sc_hd__o22a_1 _10626_ (.A1(net1676),
    .A2(\core.registers[19][23] ),
    .B1(net1375),
    .B2(\core.registers[18][23] ),
    .X(_05614_));
 sky130_fd_sc_hd__mux2_1 _10627_ (.A0(_05613_),
    .A1(_05614_),
    .S(net1437),
    .X(_05615_));
 sky130_fd_sc_hd__o21a_1 _10628_ (.A1(net1329),
    .A2(_05615_),
    .B1(net1324),
    .X(_05616_));
 sky130_fd_sc_hd__o21a_1 _10629_ (.A1(net1343),
    .A2(_05612_),
    .B1(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__o22a_1 _10630_ (.A1(net1677),
    .A2(\core.registers[7][23] ),
    .B1(net1376),
    .B2(\core.registers[6][23] ),
    .X(_05618_));
 sky130_fd_sc_hd__o22a_1 _10631_ (.A1(net1677),
    .A2(\core.registers[3][23] ),
    .B1(net1376),
    .B2(\core.registers[2][23] ),
    .X(_05619_));
 sky130_fd_sc_hd__mux2_1 _10632_ (.A0(_05618_),
    .A1(_05619_),
    .S(net1437),
    .X(_05620_));
 sky130_fd_sc_hd__or2_1 _10633_ (.A(net1329),
    .B(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__mux4_1 _10634_ (.A0(\core.registers[0][23] ),
    .A1(\core.registers[1][23] ),
    .A2(\core.registers[4][23] ),
    .A3(\core.registers[5][23] ),
    .S0(net1376),
    .S1(net1449),
    .X(_05622_));
 sky130_fd_sc_hd__o21a_1 _10635_ (.A1(net1343),
    .A2(_05622_),
    .B1(net1321),
    .X(_05623_));
 sky130_fd_sc_hd__a21oi_1 _10636_ (.A1(_05621_),
    .A2(_05623_),
    .B1(_05617_),
    .Y(_05624_));
 sky130_fd_sc_hd__o211ai_2 _10637_ (.A1(net1430),
    .A2(_05624_),
    .B1(_05611_),
    .C1(net1142),
    .Y(_05625_));
 sky130_fd_sc_hd__o211a_2 _10638_ (.A1(net1141),
    .A2(net862),
    .B1(_05625_),
    .C1(net1239),
    .X(_05626_));
 sky130_fd_sc_hd__a21o_1 _10639_ (.A1(_04072_),
    .A2(_05626_),
    .B1(net1005),
    .X(_05627_));
 sky130_fd_sc_hd__o21ai_4 _10640_ (.A1(net1762),
    .A2(net1257),
    .B1(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__mux2_1 _10641_ (.A0(\core.registers[18][23] ),
    .A1(\core.registers[19][23] ),
    .S(net1473),
    .X(_05629_));
 sky130_fd_sc_hd__mux2_1 _10642_ (.A0(\core.registers[16][23] ),
    .A1(\core.registers[17][23] ),
    .S(net1473),
    .X(_05630_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(_05629_),
    .A1(_05630_),
    .S(net1529),
    .X(_05631_));
 sky130_fd_sc_hd__o221a_1 _10644_ (.A1(net1645),
    .A2(\core.registers[23][23] ),
    .B1(net1473),
    .B2(\core.registers[22][23] ),
    .C1(net1544),
    .X(_05632_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(\core.registers[20][23] ),
    .A1(\core.registers[21][23] ),
    .S(net1473),
    .X(_05633_));
 sky130_fd_sc_hd__or2_1 _10646_ (.A(\core.registers[0][23] ),
    .B(net1474),
    .X(_05634_));
 sky130_fd_sc_hd__o211a_1 _10647_ (.A1(\core.registers[1][23] ),
    .A2(net1459),
    .B1(_05634_),
    .C1(net1529),
    .X(_05635_));
 sky130_fd_sc_hd__mux2_1 _10648_ (.A0(\core.registers[2][23] ),
    .A1(\core.registers[3][23] ),
    .S(net1474),
    .X(_05636_));
 sky130_fd_sc_hd__a211o_1 _10649_ (.A1(net1545),
    .A2(_05636_),
    .B1(_05635_),
    .C1(net1584),
    .X(_05637_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(\core.registers[4][23] ),
    .A1(\core.registers[5][23] ),
    .S(net1474),
    .X(_05638_));
 sky130_fd_sc_hd__o221a_1 _10651_ (.A1(net1645),
    .A2(\core.registers[7][23] ),
    .B1(net1474),
    .B2(\core.registers[6][23] ),
    .C1(net1544),
    .X(_05639_));
 sky130_fd_sc_hd__a211o_1 _10652_ (.A1(net1529),
    .A2(_05638_),
    .B1(_05639_),
    .C1(net1573),
    .X(_05640_));
 sky130_fd_sc_hd__a211o_1 _10653_ (.A1(net1541),
    .A2(_05633_),
    .B1(_05632_),
    .C1(net1573),
    .X(_05641_));
 sky130_fd_sc_hd__o211a_1 _10654_ (.A1(net1584),
    .A2(_05631_),
    .B1(_05641_),
    .C1(net1597),
    .X(_05642_));
 sky130_fd_sc_hd__a31o_1 _10655_ (.A1(net1593),
    .A2(_05637_),
    .A3(_05640_),
    .B1(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__mux2_1 _10656_ (.A0(\core.registers[28][23] ),
    .A1(\core.registers[29][23] ),
    .S(net1472),
    .X(_05644_));
 sky130_fd_sc_hd__a221o_1 _10657_ (.A1(net1645),
    .A2(\core.registers[30][23] ),
    .B1(\core.registers[31][23] ),
    .B2(net1472),
    .C1(net1663),
    .X(_05645_));
 sky130_fd_sc_hd__mux2_1 _10658_ (.A0(\core.registers[8][23] ),
    .A1(\core.registers[9][23] ),
    .S(net1470),
    .X(_05646_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(\core.registers[10][23] ),
    .A1(\core.registers[11][23] ),
    .S(net1470),
    .X(_05647_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(_05646_),
    .A1(_05647_),
    .S(net1544),
    .X(_05648_));
 sky130_fd_sc_hd__mux2_1 _10661_ (.A0(\core.registers[24][23] ),
    .A1(\core.registers[25][23] ),
    .S(net1470),
    .X(_05649_));
 sky130_fd_sc_hd__a22o_1 _10662_ (.A1(net1645),
    .A2(\core.registers[26][23] ),
    .B1(\core.registers[27][23] ),
    .B2(net1470),
    .X(_05650_));
 sky130_fd_sc_hd__mux2_1 _10663_ (.A0(_05649_),
    .A1(_05650_),
    .S(net1787),
    .X(_05651_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(_05648_),
    .A1(_05651_),
    .S(net1778),
    .X(_05652_));
 sky130_fd_sc_hd__o21ai_1 _10665_ (.A1(net1787),
    .A2(_05644_),
    .B1(_05645_),
    .Y(_05653_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(\core.registers[12][23] ),
    .A1(\core.registers[13][23] ),
    .S(net1470),
    .X(_05654_));
 sky130_fd_sc_hd__mux2_1 _10667_ (.A0(\core.registers[14][23] ),
    .A1(\core.registers[15][23] ),
    .S(net1470),
    .X(_05655_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(_05654_),
    .A1(_05655_),
    .S(net1544),
    .X(_05656_));
 sky130_fd_sc_hd__nor2_1 _10669_ (.A(net1778),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__a211o_1 _10670_ (.A1(net1779),
    .A2(_05653_),
    .B1(_05657_),
    .C1(net1668),
    .X(_05658_));
 sky130_fd_sc_hd__a21oi_1 _10671_ (.A1(net1668),
    .A2(_05652_),
    .B1(net1562),
    .Y(_05659_));
 sky130_fd_sc_hd__a2bb2o_1 _10672_ (.A1_N(net1567),
    .A2_N(_05643_),
    .B1(_05658_),
    .B2(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__o2bb2a_4 _10673_ (.A1_N(net1094),
    .A2_N(net861),
    .B1(_05660_),
    .B2(net1045),
    .X(_05661_));
 sky130_fd_sc_hd__mux2_8 _10674_ (.A0(_03824_),
    .A1(_05661_),
    .S(net1251),
    .X(_05662_));
 sky130_fd_sc_hd__inv_2 _10675_ (.A(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__nor2_4 _10676_ (.A(_05628_),
    .B(_05662_),
    .Y(_05664_));
 sky130_fd_sc_hd__and2_4 _10677_ (.A(_05628_),
    .B(_05662_),
    .X(_05665_));
 sky130_fd_sc_hd__a21oi_2 _10678_ (.A1(net1243),
    .A2(_04475_),
    .B1(_04022_),
    .Y(_05666_));
 sky130_fd_sc_hd__nor2_2 _10679_ (.A(net1616),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__a21o_1 _10680_ (.A1(\core.pipe1_csrData[22] ),
    .A2(net1248),
    .B1(net1238),
    .X(_05668_));
 sky130_fd_sc_hd__o21a_1 _10681_ (.A1(net1186),
    .A2(_05667_),
    .B1(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__o22a_2 _10682_ (.A1(\core.pipe1_resultRegister[22] ),
    .A2(net1189),
    .B1(_05669_),
    .B2(net1246),
    .X(_05670_));
 sky130_fd_sc_hd__mux2_1 _10683_ (.A0(\core.registers[12][22] ),
    .A1(\core.registers[13][22] ),
    .S(net1383),
    .X(_05671_));
 sky130_fd_sc_hd__mux2_1 _10684_ (.A0(\core.registers[14][22] ),
    .A1(\core.registers[15][22] ),
    .S(net1383),
    .X(_05672_));
 sky130_fd_sc_hd__mux2_1 _10685_ (.A0(_05671_),
    .A1(_05672_),
    .S(net1345),
    .X(_05673_));
 sky130_fd_sc_hd__a221o_1 _10686_ (.A1(net1682),
    .A2(\core.registers[30][22] ),
    .B1(\core.registers[31][22] ),
    .B2(net1391),
    .C1(net1702),
    .X(_05674_));
 sky130_fd_sc_hd__mux2_1 _10687_ (.A0(\core.registers[28][22] ),
    .A1(\core.registers[29][22] ),
    .S(net1391),
    .X(_05675_));
 sky130_fd_sc_hd__o21a_1 _10688_ (.A1(net1772),
    .A2(_05675_),
    .B1(_05674_),
    .X(_05676_));
 sky130_fd_sc_hd__mux2_1 _10689_ (.A0(_05673_),
    .A1(_05676_),
    .S(net1757),
    .X(_05677_));
 sky130_fd_sc_hd__mux2_1 _10690_ (.A0(\core.registers[8][22] ),
    .A1(\core.registers[9][22] ),
    .S(net1383),
    .X(_05678_));
 sky130_fd_sc_hd__mux2_1 _10691_ (.A0(\core.registers[10][22] ),
    .A1(\core.registers[11][22] ),
    .S(net1383),
    .X(_05679_));
 sky130_fd_sc_hd__mux2_1 _10692_ (.A0(_05678_),
    .A1(_05679_),
    .S(net1345),
    .X(_05680_));
 sky130_fd_sc_hd__mux2_1 _10693_ (.A0(\core.registers[24][22] ),
    .A1(\core.registers[25][22] ),
    .S(net1383),
    .X(_05681_));
 sky130_fd_sc_hd__and3_1 _10694_ (.A(net1772),
    .B(\core.registers[27][22] ),
    .C(net1383),
    .X(_05682_));
 sky130_fd_sc_hd__a211o_1 _10695_ (.A1(\core.registers[26][22] ),
    .A2(_04445_),
    .B1(_05682_),
    .C1(net1710),
    .X(_05683_));
 sky130_fd_sc_hd__a21o_1 _10696_ (.A1(net1702),
    .A2(_05681_),
    .B1(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__o211a_1 _10697_ (.A1(net1757),
    .A2(_05680_),
    .B1(_05684_),
    .C1(net1707),
    .X(_05685_));
 sky130_fd_sc_hd__mux4_1 _10698_ (.A0(\core.registers[16][22] ),
    .A1(\core.registers[17][22] ),
    .A2(\core.registers[20][22] ),
    .A3(\core.registers[21][22] ),
    .S0(net1383),
    .S1(net1451),
    .X(_05686_));
 sky130_fd_sc_hd__o22a_1 _10699_ (.A1(net1682),
    .A2(\core.registers[23][22] ),
    .B1(net1391),
    .B2(\core.registers[22][22] ),
    .X(_05687_));
 sky130_fd_sc_hd__o22a_1 _10700_ (.A1(net1682),
    .A2(\core.registers[19][22] ),
    .B1(net1393),
    .B2(\core.registers[18][22] ),
    .X(_05688_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(_05687_),
    .A1(_05688_),
    .S(net1439),
    .X(_05689_));
 sky130_fd_sc_hd__o21a_1 _10702_ (.A1(net1332),
    .A2(_05689_),
    .B1(net1325),
    .X(_05690_));
 sky130_fd_sc_hd__o21ai_1 _10703_ (.A1(net1347),
    .A2(_05686_),
    .B1(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__o22a_1 _10704_ (.A1(net1682),
    .A2(\core.registers[7][22] ),
    .B1(net1385),
    .B2(\core.registers[6][22] ),
    .X(_05692_));
 sky130_fd_sc_hd__o22a_1 _10705_ (.A1(net1682),
    .A2(\core.registers[3][22] ),
    .B1(net1385),
    .B2(\core.registers[2][22] ),
    .X(_05693_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(_05692_),
    .A1(_05693_),
    .S(net1439),
    .X(_05694_));
 sky130_fd_sc_hd__or2_1 _10707_ (.A(net1331),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__mux4_1 _10708_ (.A0(\core.registers[0][22] ),
    .A1(\core.registers[1][22] ),
    .A2(\core.registers[4][22] ),
    .A3(\core.registers[5][22] ),
    .S0(net1393),
    .S1(net1451),
    .X(_05696_));
 sky130_fd_sc_hd__o21a_1 _10709_ (.A1(net1348),
    .A2(_05696_),
    .B1(net1321),
    .X(_05697_));
 sky130_fd_sc_hd__a21oi_1 _10710_ (.A1(_05695_),
    .A2(_05697_),
    .B1(net1431),
    .Y(_05698_));
 sky130_fd_sc_hd__a21o_1 _10711_ (.A1(net1764),
    .A2(_05677_),
    .B1(net1428),
    .X(_05699_));
 sky130_fd_sc_hd__o2bb2a_2 _10712_ (.A1_N(_05691_),
    .A2_N(_05698_),
    .B1(_05699_),
    .B2(_05685_),
    .X(_05700_));
 sky130_fd_sc_hd__o21a_1 _10713_ (.A1(net1146),
    .A2(net859),
    .B1(net1241),
    .X(_05701_));
 sky130_fd_sc_hd__o21ai_4 _10714_ (.A1(net1149),
    .A2(_05700_),
    .B1(_05701_),
    .Y(_05702_));
 sky130_fd_sc_hd__nor2_1 _10715_ (.A(net1039),
    .B(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__o22a_4 _10716_ (.A1(net1764),
    .A2(net1252),
    .B1(net1005),
    .B2(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__mux2_1 _10717_ (.A0(\core.registers[18][22] ),
    .A1(\core.registers[19][22] ),
    .S(net1492),
    .X(_05705_));
 sky130_fd_sc_hd__mux2_1 _10718_ (.A0(\core.registers[16][22] ),
    .A1(\core.registers[17][22] ),
    .S(net1482),
    .X(_05706_));
 sky130_fd_sc_hd__mux2_1 _10719_ (.A0(_05705_),
    .A1(_05706_),
    .S(net1531),
    .X(_05707_));
 sky130_fd_sc_hd__o221a_1 _10720_ (.A1(net1648),
    .A2(\core.registers[23][22] ),
    .B1(net1490),
    .B2(\core.registers[22][22] ),
    .C1(net1551),
    .X(_05708_));
 sky130_fd_sc_hd__mux2_1 _10721_ (.A0(\core.registers[20][22] ),
    .A1(\core.registers[21][22] ),
    .S(net1494),
    .X(_05709_));
 sky130_fd_sc_hd__or2_1 _10722_ (.A(\core.registers[0][22] ),
    .B(net1484),
    .X(_05710_));
 sky130_fd_sc_hd__o211a_1 _10723_ (.A1(\core.registers[1][22] ),
    .A2(net1459),
    .B1(_05710_),
    .C1(net1531),
    .X(_05711_));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(\core.registers[2][22] ),
    .A1(\core.registers[3][22] ),
    .S(net1484),
    .X(_05712_));
 sky130_fd_sc_hd__a211o_1 _10725_ (.A1(net1547),
    .A2(_05712_),
    .B1(_05711_),
    .C1(net1585),
    .X(_05713_));
 sky130_fd_sc_hd__mux2_1 _10726_ (.A0(\core.registers[4][22] ),
    .A1(\core.registers[5][22] ),
    .S(net1484),
    .X(_05714_));
 sky130_fd_sc_hd__o221a_1 _10727_ (.A1(net1649),
    .A2(\core.registers[7][22] ),
    .B1(net1484),
    .B2(\core.registers[6][22] ),
    .C1(net1547),
    .X(_05715_));
 sky130_fd_sc_hd__a211o_1 _10728_ (.A1(net1531),
    .A2(_05714_),
    .B1(_05715_),
    .C1(net1574),
    .X(_05716_));
 sky130_fd_sc_hd__a211o_1 _10729_ (.A1(net1531),
    .A2(_05709_),
    .B1(_05708_),
    .C1(net1575),
    .X(_05717_));
 sky130_fd_sc_hd__o211a_1 _10730_ (.A1(net1585),
    .A2(_05707_),
    .B1(_05717_),
    .C1(net1598),
    .X(_05718_));
 sky130_fd_sc_hd__a311o_2 _10731_ (.A1(net1594),
    .A2(_05713_),
    .A3(_05716_),
    .B1(_05718_),
    .C1(net1570),
    .X(_05719_));
 sky130_fd_sc_hd__mux2_1 _10732_ (.A0(\core.registers[8][22] ),
    .A1(\core.registers[9][22] ),
    .S(net1482),
    .X(_05720_));
 sky130_fd_sc_hd__mux2_1 _10733_ (.A0(\core.registers[10][22] ),
    .A1(\core.registers[11][22] ),
    .S(net1482),
    .X(_05721_));
 sky130_fd_sc_hd__mux2_1 _10734_ (.A0(\core.registers[28][22] ),
    .A1(\core.registers[29][22] ),
    .S(net1482),
    .X(_05722_));
 sky130_fd_sc_hd__a221o_1 _10735_ (.A1(net1648),
    .A2(\core.registers[30][22] ),
    .B1(\core.registers[31][22] ),
    .B2(net1490),
    .C1(net1666),
    .X(_05723_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(_05720_),
    .A1(_05721_),
    .S(net1547),
    .X(_05724_));
 sky130_fd_sc_hd__or2_1 _10737_ (.A(\core.registers[24][22] ),
    .B(net1482),
    .X(_05725_));
 sky130_fd_sc_hd__o21a_1 _10738_ (.A1(\core.registers[25][22] ),
    .A2(net1459),
    .B1(net1666),
    .X(_05726_));
 sky130_fd_sc_hd__a22o_1 _10739_ (.A1(net1648),
    .A2(\core.registers[26][22] ),
    .B1(\core.registers[27][22] ),
    .B2(net1482),
    .X(_05727_));
 sky130_fd_sc_hd__a221o_1 _10740_ (.A1(_05725_),
    .A2(_05726_),
    .B1(_05727_),
    .B2(net1791),
    .C1(net1673),
    .X(_05728_));
 sky130_fd_sc_hd__o211a_1 _10741_ (.A1(net1782),
    .A2(_05724_),
    .B1(_05728_),
    .C1(net1670),
    .X(_05729_));
 sky130_fd_sc_hd__o21a_1 _10742_ (.A1(net1791),
    .A2(_05722_),
    .B1(_05723_),
    .X(_05730_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\core.registers[12][22] ),
    .A1(\core.registers[13][22] ),
    .S(net1482),
    .X(_05731_));
 sky130_fd_sc_hd__mux2_1 _10744_ (.A0(\core.registers[14][22] ),
    .A1(\core.registers[15][22] ),
    .S(net1482),
    .X(_05732_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(_05731_),
    .A1(_05732_),
    .S(net1547),
    .X(_05733_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(_05730_),
    .A1(_05733_),
    .S(net1673),
    .X(_05734_));
 sky130_fd_sc_hd__a21o_1 _10747_ (.A1(net1785),
    .A2(_05734_),
    .B1(_03886_),
    .X(_05735_));
 sky130_fd_sc_hd__o21ai_4 _10748_ (.A1(_05729_),
    .A2(_05735_),
    .B1(_05719_),
    .Y(_05736_));
 sky130_fd_sc_hd__o2bb2a_4 _10749_ (.A1_N(net1096),
    .A2_N(net859),
    .B1(_05736_),
    .B2(net1044),
    .X(_05737_));
 sky130_fd_sc_hd__inv_2 _10750_ (.A(_05737_),
    .Y(_05738_));
 sky130_fd_sc_hd__mux2_4 _10751_ (.A0(net464),
    .A1(_05738_),
    .S(net1251),
    .X(_05739_));
 sky130_fd_sc_hd__and2_4 _10752_ (.A(_05704_),
    .B(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__nor2_4 _10753_ (.A(_05704_),
    .B(_05739_),
    .Y(_05741_));
 sky130_fd_sc_hd__nor2_8 _10754_ (.A(_05740_),
    .B(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__clkinv_2 _10755_ (.A(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__a21oi_1 _10756_ (.A1(net1243),
    .A2(_04560_),
    .B1(_04022_),
    .Y(_05744_));
 sky130_fd_sc_hd__nor2_1 _10757_ (.A(net1616),
    .B(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__a21o_1 _10758_ (.A1(\core.pipe1_csrData[21] ),
    .A2(net1248),
    .B1(net1238),
    .X(_05746_));
 sky130_fd_sc_hd__o21a_1 _10759_ (.A1(net1186),
    .A2(_05745_),
    .B1(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__o22a_4 _10760_ (.A1(\core.pipe1_resultRegister[21] ),
    .A2(net1189),
    .B1(_05747_),
    .B2(net1246),
    .X(_05748_));
 sky130_fd_sc_hd__mux2_1 _10761_ (.A0(\core.registers[12][21] ),
    .A1(\core.registers[13][21] ),
    .S(net1363),
    .X(_05749_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(\core.registers[14][21] ),
    .A1(\core.registers[15][21] ),
    .S(net1363),
    .X(_05750_));
 sky130_fd_sc_hd__mux2_1 _10763_ (.A0(_05749_),
    .A1(_05750_),
    .S(net1341),
    .X(_05751_));
 sky130_fd_sc_hd__a221o_1 _10764_ (.A1(net1675),
    .A2(\core.registers[30][21] ),
    .B1(\core.registers[31][21] ),
    .B2(net1365),
    .C1(net1699),
    .X(_05752_));
 sky130_fd_sc_hd__mux2_1 _10765_ (.A0(\core.registers[28][21] ),
    .A1(\core.registers[29][21] ),
    .S(net1364),
    .X(_05753_));
 sky130_fd_sc_hd__o21a_1 _10766_ (.A1(net1768),
    .A2(_05753_),
    .B1(_05752_),
    .X(_05754_));
 sky130_fd_sc_hd__mux2_1 _10767_ (.A0(_05751_),
    .A1(_05754_),
    .S(net1753),
    .X(_05755_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(\core.registers[8][21] ),
    .A1(\core.registers[9][21] ),
    .S(net1363),
    .X(_05756_));
 sky130_fd_sc_hd__mux2_1 _10769_ (.A0(\core.registers[10][21] ),
    .A1(\core.registers[11][21] ),
    .S(net1363),
    .X(_05757_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(_05756_),
    .A1(_05757_),
    .S(net1341),
    .X(_05758_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(\core.registers[24][21] ),
    .A1(\core.registers[25][21] ),
    .S(net1371),
    .X(_05759_));
 sky130_fd_sc_hd__and3_1 _10772_ (.A(net1768),
    .B(\core.registers[27][21] ),
    .C(net1371),
    .X(_05760_));
 sky130_fd_sc_hd__a211o_1 _10773_ (.A1(\core.registers[26][21] ),
    .A2(net1319),
    .B1(_05760_),
    .C1(net1708),
    .X(_05761_));
 sky130_fd_sc_hd__a21o_1 _10774_ (.A1(net1699),
    .A2(_05759_),
    .B1(_05761_),
    .X(_05762_));
 sky130_fd_sc_hd__o211a_1 _10775_ (.A1(net1753),
    .A2(_05758_),
    .B1(_05762_),
    .C1(net1704),
    .X(_05763_));
 sky130_fd_sc_hd__mux4_1 _10776_ (.A0(\core.registers[16][21] ),
    .A1(\core.registers[17][21] ),
    .A2(\core.registers[20][21] ),
    .A3(\core.registers[21][21] ),
    .S0(net1368),
    .S1(net1447),
    .X(_05764_));
 sky130_fd_sc_hd__o22a_1 _10777_ (.A1(net1675),
    .A2(\core.registers[23][21] ),
    .B1(net1368),
    .B2(\core.registers[22][21] ),
    .X(_05765_));
 sky130_fd_sc_hd__o22a_1 _10778_ (.A1(net1675),
    .A2(\core.registers[19][21] ),
    .B1(net1368),
    .B2(\core.registers[18][21] ),
    .X(_05766_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(_05765_),
    .A1(_05766_),
    .S(net1434),
    .X(_05767_));
 sky130_fd_sc_hd__o21a_1 _10780_ (.A1(net1328),
    .A2(_05767_),
    .B1(net1324),
    .X(_05768_));
 sky130_fd_sc_hd__o21ai_1 _10781_ (.A1(net1341),
    .A2(_05764_),
    .B1(_05768_),
    .Y(_05769_));
 sky130_fd_sc_hd__o22a_1 _10782_ (.A1(net1678),
    .A2(\core.registers[7][21] ),
    .B1(net1369),
    .B2(\core.registers[6][21] ),
    .X(_05770_));
 sky130_fd_sc_hd__o22a_1 _10783_ (.A1(net1677),
    .A2(\core.registers[3][21] ),
    .B1(net1369),
    .B2(\core.registers[2][21] ),
    .X(_05771_));
 sky130_fd_sc_hd__mux2_1 _10784_ (.A0(_05770_),
    .A1(_05771_),
    .S(net1434),
    .X(_05772_));
 sky130_fd_sc_hd__or2_1 _10785_ (.A(net1328),
    .B(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__mux4_1 _10786_ (.A0(\core.registers[0][21] ),
    .A1(\core.registers[1][21] ),
    .A2(\core.registers[4][21] ),
    .A3(\core.registers[5][21] ),
    .S0(net1369),
    .S1(net1448),
    .X(_05774_));
 sky130_fd_sc_hd__o21a_1 _10787_ (.A1(net1342),
    .A2(_05774_),
    .B1(net1320),
    .X(_05775_));
 sky130_fd_sc_hd__a21oi_1 _10788_ (.A1(_05773_),
    .A2(_05775_),
    .B1(net1429),
    .Y(_05776_));
 sky130_fd_sc_hd__a21o_1 _10789_ (.A1(net1763),
    .A2(_05755_),
    .B1(net1427),
    .X(_05777_));
 sky130_fd_sc_hd__o2bb2a_2 _10790_ (.A1_N(_05769_),
    .A2_N(_05776_),
    .B1(_05777_),
    .B2(_05763_),
    .X(_05778_));
 sky130_fd_sc_hd__o21a_1 _10791_ (.A1(net1148),
    .A2(_05778_),
    .B1(net1239),
    .X(_05779_));
 sky130_fd_sc_hd__o21ai_1 _10792_ (.A1(net1141),
    .A2(net854),
    .B1(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__nor2_1 _10793_ (.A(net1039),
    .B(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__o22a_2 _10794_ (.A1(net1771),
    .A2(net1252),
    .B1(net1005),
    .B2(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(\core.registers[18][21] ),
    .A1(\core.registers[19][21] ),
    .S(net1467),
    .X(_05783_));
 sky130_fd_sc_hd__mux2_1 _10796_ (.A0(\core.registers[16][21] ),
    .A1(\core.registers[17][21] ),
    .S(net1467),
    .X(_05784_));
 sky130_fd_sc_hd__mux2_1 _10797_ (.A0(_05783_),
    .A1(_05784_),
    .S(net1526),
    .X(_05785_));
 sky130_fd_sc_hd__o221a_1 _10798_ (.A1(net1642),
    .A2(\core.registers[23][21] ),
    .B1(net1467),
    .B2(\core.registers[22][21] ),
    .C1(net1542),
    .X(_05786_));
 sky130_fd_sc_hd__mux2_1 _10799_ (.A0(\core.registers[20][21] ),
    .A1(\core.registers[21][21] ),
    .S(net1467),
    .X(_05787_));
 sky130_fd_sc_hd__or2_1 _10800_ (.A(\core.registers[0][21] ),
    .B(net1468),
    .X(_05788_));
 sky130_fd_sc_hd__o211a_1 _10801_ (.A1(\core.registers[1][21] ),
    .A2(net1459),
    .B1(_05788_),
    .C1(net1528),
    .X(_05789_));
 sky130_fd_sc_hd__mux2_1 _10802_ (.A0(\core.registers[2][21] ),
    .A1(\core.registers[3][21] ),
    .S(net1468),
    .X(_05790_));
 sky130_fd_sc_hd__a211o_1 _10803_ (.A1(net1542),
    .A2(_05790_),
    .B1(_05789_),
    .C1(net1583),
    .X(_05791_));
 sky130_fd_sc_hd__mux2_1 _10804_ (.A0(\core.registers[4][21] ),
    .A1(\core.registers[5][21] ),
    .S(net1468),
    .X(_05792_));
 sky130_fd_sc_hd__o221a_1 _10805_ (.A1(net1644),
    .A2(\core.registers[7][21] ),
    .B1(net1467),
    .B2(\core.registers[6][21] ),
    .C1(net1542),
    .X(_05793_));
 sky130_fd_sc_hd__a211o_1 _10806_ (.A1(net1527),
    .A2(_05792_),
    .B1(_05793_),
    .C1(net1571),
    .X(_05794_));
 sky130_fd_sc_hd__a211o_1 _10807_ (.A1(net1526),
    .A2(_05787_),
    .B1(_05786_),
    .C1(net1571),
    .X(_05795_));
 sky130_fd_sc_hd__o211a_1 _10808_ (.A1(net1582),
    .A2(_05785_),
    .B1(_05795_),
    .C1(net1597),
    .X(_05796_));
 sky130_fd_sc_hd__a311o_4 _10809_ (.A1(net1593),
    .A2(_05791_),
    .A3(_05794_),
    .B1(_05796_),
    .C1(net1566),
    .X(_05797_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(\core.registers[8][21] ),
    .A1(\core.registers[9][21] ),
    .S(net1462),
    .X(_05798_));
 sky130_fd_sc_hd__mux2_1 _10811_ (.A0(\core.registers[10][21] ),
    .A1(\core.registers[11][21] ),
    .S(net1462),
    .X(_05799_));
 sky130_fd_sc_hd__mux2_1 _10812_ (.A0(\core.registers[28][21] ),
    .A1(\core.registers[29][21] ),
    .S(net1463),
    .X(_05800_));
 sky130_fd_sc_hd__a221o_1 _10813_ (.A1(net1641),
    .A2(\core.registers[30][21] ),
    .B1(\core.registers[31][21] ),
    .B2(net1464),
    .C1(net1663),
    .X(_05801_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(_05798_),
    .A1(_05799_),
    .S(net1543),
    .X(_05802_));
 sky130_fd_sc_hd__or2_1 _10815_ (.A(\core.registers[24][21] ),
    .B(net1463),
    .X(_05803_));
 sky130_fd_sc_hd__o21a_1 _10816_ (.A1(\core.registers[25][21] ),
    .A2(net1459),
    .B1(net1663),
    .X(_05804_));
 sky130_fd_sc_hd__a22o_1 _10817_ (.A1(net1646),
    .A2(\core.registers[26][21] ),
    .B1(\core.registers[27][21] ),
    .B2(net1464),
    .X(_05805_));
 sky130_fd_sc_hd__a221o_1 _10818_ (.A1(_05803_),
    .A2(_05804_),
    .B1(_05805_),
    .B2(net1787),
    .C1(net1674),
    .X(_05806_));
 sky130_fd_sc_hd__o211a_1 _10819_ (.A1(net1778),
    .A2(_05802_),
    .B1(_05806_),
    .C1(net1668),
    .X(_05807_));
 sky130_fd_sc_hd__mux2_1 _10820_ (.A0(\core.registers[12][21] ),
    .A1(\core.registers[13][21] ),
    .S(net1462),
    .X(_05808_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(\core.registers[14][21] ),
    .A1(\core.registers[15][21] ),
    .S(net1462),
    .X(_05809_));
 sky130_fd_sc_hd__mux2_1 _10822_ (.A0(_05808_),
    .A1(_05809_),
    .S(net1543),
    .X(_05810_));
 sky130_fd_sc_hd__o21a_1 _10823_ (.A1(net1787),
    .A2(_05800_),
    .B1(_05801_),
    .X(_05811_));
 sky130_fd_sc_hd__mux2_1 _10824_ (.A0(_05810_),
    .A1(_05811_),
    .S(net1778),
    .X(_05812_));
 sky130_fd_sc_hd__a21o_1 _10825_ (.A1(net1784),
    .A2(_05812_),
    .B1(net1561),
    .X(_05813_));
 sky130_fd_sc_hd__o21ai_4 _10826_ (.A1(_05807_),
    .A2(_05813_),
    .B1(_05797_),
    .Y(_05814_));
 sky130_fd_sc_hd__o2bb2a_2 _10827_ (.A1_N(net1094),
    .A2_N(net854),
    .B1(_05814_),
    .B2(net1045),
    .X(_05815_));
 sky130_fd_sc_hd__inv_2 _10828_ (.A(_05815_),
    .Y(_05816_));
 sky130_fd_sc_hd__mux2_4 _10829_ (.A0(net463),
    .A1(_05816_),
    .S(net1256),
    .X(_05817_));
 sky130_fd_sc_hd__or2_2 _10830_ (.A(_05782_),
    .B(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__clkinv_2 _10831_ (.A(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__and2_4 _10832_ (.A(_05782_),
    .B(_05817_),
    .X(_05820_));
 sky130_fd_sc_hd__a21oi_1 _10833_ (.A1(net1243),
    .A2(_04646_),
    .B1(_04022_),
    .Y(_05821_));
 sky130_fd_sc_hd__nor2_1 _10834_ (.A(_04002_),
    .B(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__a21o_1 _10835_ (.A1(\core.pipe1_csrData[20] ),
    .A2(net1247),
    .B1(net1238),
    .X(_05823_));
 sky130_fd_sc_hd__o21a_1 _10836_ (.A1(net1186),
    .A2(_05822_),
    .B1(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__o22a_4 _10837_ (.A1(\core.pipe1_resultRegister[20] ),
    .A2(net1188),
    .B1(_05824_),
    .B2(net1246),
    .X(_05825_));
 sky130_fd_sc_hd__or2_1 _10838_ (.A(\core.registers[5][20] ),
    .B(net1358),
    .X(_05826_));
 sky130_fd_sc_hd__o211a_1 _10839_ (.A1(\core.registers[4][20] ),
    .A2(net1389),
    .B1(_05826_),
    .C1(net1449),
    .X(_05827_));
 sky130_fd_sc_hd__mux2_1 _10840_ (.A0(\core.registers[0][20] ),
    .A1(\core.registers[1][20] ),
    .S(net1389),
    .X(_05828_));
 sky130_fd_sc_hd__a211o_1 _10841_ (.A1(net1435),
    .A2(_05828_),
    .B1(_05827_),
    .C1(net1356),
    .X(_05829_));
 sky130_fd_sc_hd__o221a_1 _10842_ (.A1(net1677),
    .A2(\core.registers[7][20] ),
    .B1(net1379),
    .B2(\core.registers[6][20] ),
    .C1(net1449),
    .X(_05830_));
 sky130_fd_sc_hd__o221a_1 _10843_ (.A1(net1679),
    .A2(\core.registers[3][20] ),
    .B1(net1379),
    .B2(\core.registers[2][20] ),
    .C1(net1435),
    .X(_05831_));
 sky130_fd_sc_hd__o31a_1 _10844_ (.A1(net1330),
    .A2(_05830_),
    .A3(_05831_),
    .B1(net1320),
    .X(_05832_));
 sky130_fd_sc_hd__or2_1 _10845_ (.A(\core.registers[16][20] ),
    .B(net1368),
    .X(_05833_));
 sky130_fd_sc_hd__o211a_1 _10846_ (.A1(\core.registers[17][20] ),
    .A2(net1357),
    .B1(_05833_),
    .C1(net1436),
    .X(_05834_));
 sky130_fd_sc_hd__mux2_1 _10847_ (.A0(\core.registers[20][20] ),
    .A1(\core.registers[21][20] ),
    .S(net1368),
    .X(_05835_));
 sky130_fd_sc_hd__a211o_1 _10848_ (.A1(net1447),
    .A2(_05835_),
    .B1(_05834_),
    .C1(net1341),
    .X(_05836_));
 sky130_fd_sc_hd__o221a_1 _10849_ (.A1(net1677),
    .A2(\core.registers[23][20] ),
    .B1(net1368),
    .B2(\core.registers[22][20] ),
    .C1(net1447),
    .X(_05837_));
 sky130_fd_sc_hd__o221a_1 _10850_ (.A1(net1677),
    .A2(\core.registers[19][20] ),
    .B1(net1368),
    .B2(\core.registers[18][20] ),
    .C1(net1436),
    .X(_05838_));
 sky130_fd_sc_hd__o31a_1 _10851_ (.A1(net1328),
    .A2(_05837_),
    .A3(_05838_),
    .B1(net1324),
    .X(_05839_));
 sky130_fd_sc_hd__mux2_1 _10852_ (.A0(\core.registers[12][20] ),
    .A1(\core.registers[13][20] ),
    .S(net1368),
    .X(_05840_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(\core.registers[14][20] ),
    .A1(\core.registers[15][20] ),
    .S(net1368),
    .X(_05841_));
 sky130_fd_sc_hd__mux2_1 _10854_ (.A0(_05840_),
    .A1(_05841_),
    .S(net1341),
    .X(_05842_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(\core.registers[28][20] ),
    .A1(\core.registers[29][20] ),
    .S(net1364),
    .X(_05843_));
 sky130_fd_sc_hd__and3_1 _10856_ (.A(net1769),
    .B(\core.registers[31][20] ),
    .C(net1371),
    .X(_05844_));
 sky130_fd_sc_hd__a211o_1 _10857_ (.A1(\core.registers[30][20] ),
    .A2(net1319),
    .B1(_05844_),
    .C1(net1708),
    .X(_05845_));
 sky130_fd_sc_hd__a21o_1 _10858_ (.A1(net1699),
    .A2(_05843_),
    .B1(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__o211a_1 _10859_ (.A1(net1753),
    .A2(_05842_),
    .B1(_05846_),
    .C1(net1763),
    .X(_05847_));
 sky130_fd_sc_hd__or2_1 _10860_ (.A(\core.registers[9][20] ),
    .B(net1357),
    .X(_05848_));
 sky130_fd_sc_hd__o211a_1 _10861_ (.A1(\core.registers[8][20] ),
    .A2(net1368),
    .B1(net1328),
    .C1(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__a22o_1 _10862_ (.A1(net1676),
    .A2(\core.registers[10][20] ),
    .B1(\core.registers[11][20] ),
    .B2(net1364),
    .X(_05850_));
 sky130_fd_sc_hd__a21o_1 _10863_ (.A1(net1341),
    .A2(_05850_),
    .B1(net1753),
    .X(_05851_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(\core.registers[24][20] ),
    .A1(\core.registers[25][20] ),
    .S(net1364),
    .X(_05852_));
 sky130_fd_sc_hd__a22o_1 _10865_ (.A1(net1679),
    .A2(\core.registers[26][20] ),
    .B1(\core.registers[27][20] ),
    .B2(net1364),
    .X(_05853_));
 sky130_fd_sc_hd__mux2_1 _10866_ (.A0(_05852_),
    .A1(_05853_),
    .S(net1769),
    .X(_05854_));
 sky130_fd_sc_hd__o221a_1 _10867_ (.A1(_05849_),
    .A2(_05851_),
    .B1(_05854_),
    .B2(net1708),
    .C1(net1704),
    .X(_05855_));
 sky130_fd_sc_hd__a21o_1 _10868_ (.A1(_05829_),
    .A2(_05832_),
    .B1(net1429),
    .X(_05856_));
 sky130_fd_sc_hd__a21o_1 _10869_ (.A1(_05836_),
    .A2(_05839_),
    .B1(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__o31a_1 _10870_ (.A1(net1427),
    .A2(_05847_),
    .A3(_05855_),
    .B1(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__o21a_1 _10871_ (.A1(net1141),
    .A2(net849),
    .B1(net1239),
    .X(_05859_));
 sky130_fd_sc_hd__o21ai_1 _10872_ (.A1(net1148),
    .A2(_05858_),
    .B1(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__nor2_1 _10873_ (.A(net1039),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__o22a_4 _10874_ (.A1(net1776),
    .A2(net1252),
    .B1(net1005),
    .B2(_05861_),
    .X(_05862_));
 sky130_fd_sc_hd__mux4_1 _10875_ (.A0(\core.registers[8][20] ),
    .A1(\core.registers[9][20] ),
    .A2(\core.registers[12][20] ),
    .A3(\core.registers[13][20] ),
    .S0(net1467),
    .S1(net1582),
    .X(_05863_));
 sky130_fd_sc_hd__nand2_1 _10876_ (.A(net1527),
    .B(_05863_),
    .Y(_05864_));
 sky130_fd_sc_hd__a22o_1 _10877_ (.A1(net1642),
    .A2(\core.registers[14][20] ),
    .B1(\core.registers[15][20] ),
    .B2(net1467),
    .X(_05865_));
 sky130_fd_sc_hd__a22o_1 _10878_ (.A1(net1642),
    .A2(\core.registers[10][20] ),
    .B1(\core.registers[11][20] ),
    .B2(net1463),
    .X(_05866_));
 sky130_fd_sc_hd__mux2_1 _10879_ (.A0(_05865_),
    .A1(_05866_),
    .S(net1572),
    .X(_05867_));
 sky130_fd_sc_hd__a21oi_1 _10880_ (.A1(net1542),
    .A2(_05867_),
    .B1(net1562),
    .Y(_05868_));
 sky130_fd_sc_hd__mux4_1 _10881_ (.A0(\core.registers[0][20] ),
    .A1(\core.registers[1][20] ),
    .A2(\core.registers[4][20] ),
    .A3(\core.registers[5][20] ),
    .S0(net1486),
    .S1(net1584),
    .X(_05869_));
 sky130_fd_sc_hd__and2_1 _10882_ (.A(net1527),
    .B(_05869_),
    .X(_05870_));
 sky130_fd_sc_hd__a22o_1 _10883_ (.A1(net1644),
    .A2(\core.registers[6][20] ),
    .B1(\core.registers[7][20] ),
    .B2(net1478),
    .X(_05871_));
 sky130_fd_sc_hd__a22o_1 _10884_ (.A1(net1644),
    .A2(\core.registers[2][20] ),
    .B1(\core.registers[3][20] ),
    .B2(net1478),
    .X(_05872_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(_05871_),
    .A1(_05872_),
    .S(net1572),
    .X(_05873_));
 sky130_fd_sc_hd__a21o_1 _10886_ (.A1(net1546),
    .A2(_05873_),
    .B1(net1566),
    .X(_05874_));
 sky130_fd_sc_hd__nor2_1 _10887_ (.A(_05870_),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__a22o_1 _10888_ (.A1(net1642),
    .A2(\core.registers[30][20] ),
    .B1(\core.registers[31][20] ),
    .B2(net1463),
    .X(_05876_));
 sky130_fd_sc_hd__a22o_1 _10889_ (.A1(net1642),
    .A2(\core.registers[26][20] ),
    .B1(\core.registers[27][20] ),
    .B2(net1463),
    .X(_05877_));
 sky130_fd_sc_hd__mux2_1 _10890_ (.A0(_05876_),
    .A1(_05877_),
    .S(net1571),
    .X(_05878_));
 sky130_fd_sc_hd__mux4_1 _10891_ (.A0(\core.registers[24][20] ),
    .A1(\core.registers[25][20] ),
    .A2(\core.registers[28][20] ),
    .A3(\core.registers[29][20] ),
    .S0(net1463),
    .S1(net1582),
    .X(_05879_));
 sky130_fd_sc_hd__a21o_1 _10892_ (.A1(net1526),
    .A2(_05879_),
    .B1(net1561),
    .X(_05880_));
 sky130_fd_sc_hd__a21oi_1 _10893_ (.A1(net1543),
    .A2(_05878_),
    .B1(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__mux4_1 _10894_ (.A0(\core.registers[16][20] ),
    .A1(\core.registers[17][20] ),
    .A2(\core.registers[20][20] ),
    .A3(\core.registers[21][20] ),
    .S0(net1467),
    .S1(net1582),
    .X(_05882_));
 sky130_fd_sc_hd__a22o_1 _10895_ (.A1(net1644),
    .A2(\core.registers[22][20] ),
    .B1(\core.registers[23][20] ),
    .B2(net1468),
    .X(_05883_));
 sky130_fd_sc_hd__a22o_1 _10896_ (.A1(net1644),
    .A2(\core.registers[18][20] ),
    .B1(\core.registers[19][20] ),
    .B2(net1468),
    .X(_05884_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(_05883_),
    .A1(_05884_),
    .S(net1572),
    .X(_05885_));
 sky130_fd_sc_hd__a21o_1 _10898_ (.A1(net1543),
    .A2(_05885_),
    .B1(net1566),
    .X(_05886_));
 sky130_fd_sc_hd__a21oi_1 _10899_ (.A1(net1527),
    .A2(_05882_),
    .B1(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__a21o_1 _10900_ (.A1(_05864_),
    .A2(_05868_),
    .B1(net1597),
    .X(_05888_));
 sky130_fd_sc_hd__or3_1 _10901_ (.A(net1593),
    .B(_05881_),
    .C(_05887_),
    .X(_05889_));
 sky130_fd_sc_hd__o21a_1 _10902_ (.A1(_05875_),
    .A2(_05888_),
    .B1(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__o2bb2a_2 _10903_ (.A1_N(net1094),
    .A2_N(net849),
    .B1(_05890_),
    .B2(net1045),
    .X(_05891_));
 sky130_fd_sc_hd__inv_2 _10904_ (.A(_05891_),
    .Y(_05892_));
 sky130_fd_sc_hd__mux2_4 _10905_ (.A0(net462),
    .A1(_05892_),
    .S(net1256),
    .X(_05893_));
 sky130_fd_sc_hd__inv_2 _10906_ (.A(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__and2_4 _10907_ (.A(_05862_),
    .B(_05893_),
    .X(_05895_));
 sky130_fd_sc_hd__nor2_4 _10908_ (.A(_05862_),
    .B(_05893_),
    .Y(_05896_));
 sky130_fd_sc_hd__nor2_8 _10909_ (.A(_05895_),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__a21oi_1 _10910_ (.A1(net1617),
    .A2(_04025_),
    .B1(net1186),
    .Y(_05898_));
 sky130_fd_sc_hd__a21oi_1 _10911_ (.A1(\core.pipe1_csrData[19] ),
    .A2(net1247),
    .B1(net1238),
    .Y(_05899_));
 sky130_fd_sc_hd__nor2_1 _10912_ (.A(_05898_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__o22a_4 _10913_ (.A1(\core.pipe1_resultRegister[19] ),
    .A2(net1189),
    .B1(_05900_),
    .B2(net1246),
    .X(_05901_));
 sky130_fd_sc_hd__or2_1 _10914_ (.A(\core.registers[5][19] ),
    .B(net1357),
    .X(_05902_));
 sky130_fd_sc_hd__o211a_1 _10915_ (.A1(\core.registers[4][19] ),
    .A2(net1379),
    .B1(_05902_),
    .C1(net1448),
    .X(_05903_));
 sky130_fd_sc_hd__mux2_1 _10916_ (.A0(\core.registers[0][19] ),
    .A1(\core.registers[1][19] ),
    .S(net1379),
    .X(_05904_));
 sky130_fd_sc_hd__a211o_1 _10917_ (.A1(net1435),
    .A2(_05904_),
    .B1(_05903_),
    .C1(net1344),
    .X(_05905_));
 sky130_fd_sc_hd__o221a_1 _10918_ (.A1(net1678),
    .A2(\core.registers[7][19] ),
    .B1(net1378),
    .B2(\core.registers[6][19] ),
    .C1(net1449),
    .X(_05906_));
 sky130_fd_sc_hd__o221a_1 _10919_ (.A1(net1678),
    .A2(\core.registers[3][19] ),
    .B1(net1378),
    .B2(\core.registers[2][19] ),
    .C1(net1435),
    .X(_05907_));
 sky130_fd_sc_hd__o31a_1 _10920_ (.A1(net1328),
    .A2(_05906_),
    .A3(_05907_),
    .B1(net1320),
    .X(_05908_));
 sky130_fd_sc_hd__or2_1 _10921_ (.A(\core.registers[16][19] ),
    .B(net1367),
    .X(_05909_));
 sky130_fd_sc_hd__o211a_1 _10922_ (.A1(\core.registers[17][19] ),
    .A2(net1357),
    .B1(_05909_),
    .C1(net1434),
    .X(_05910_));
 sky130_fd_sc_hd__mux2_1 _10923_ (.A0(\core.registers[20][19] ),
    .A1(\core.registers[21][19] ),
    .S(net1367),
    .X(_05911_));
 sky130_fd_sc_hd__a211o_1 _10924_ (.A1(net1447),
    .A2(_05911_),
    .B1(_05910_),
    .C1(net1342),
    .X(_05912_));
 sky130_fd_sc_hd__o221a_1 _10925_ (.A1(net1675),
    .A2(\core.registers[23][19] ),
    .B1(net1366),
    .B2(\core.registers[22][19] ),
    .C1(net1447),
    .X(_05913_));
 sky130_fd_sc_hd__o221a_1 _10926_ (.A1(net1675),
    .A2(\core.registers[19][19] ),
    .B1(net1366),
    .B2(\core.registers[18][19] ),
    .C1(net1434),
    .X(_05914_));
 sky130_fd_sc_hd__o31a_1 _10927_ (.A1(net1328),
    .A2(_05913_),
    .A3(_05914_),
    .B1(net1324),
    .X(_05915_));
 sky130_fd_sc_hd__mux2_1 _10928_ (.A0(\core.registers[12][19] ),
    .A1(\core.registers[13][19] ),
    .S(net1366),
    .X(_05916_));
 sky130_fd_sc_hd__mux2_1 _10929_ (.A0(\core.registers[14][19] ),
    .A1(\core.registers[15][19] ),
    .S(net1370),
    .X(_05917_));
 sky130_fd_sc_hd__mux2_1 _10930_ (.A0(_05916_),
    .A1(_05917_),
    .S(net1342),
    .X(_05918_));
 sky130_fd_sc_hd__mux2_1 _10931_ (.A0(\core.registers[28][19] ),
    .A1(\core.registers[29][19] ),
    .S(net1366),
    .X(_05919_));
 sky130_fd_sc_hd__and3_1 _10932_ (.A(net1768),
    .B(\core.registers[31][19] ),
    .C(net1366),
    .X(_05920_));
 sky130_fd_sc_hd__a31o_1 _10933_ (.A1(net1768),
    .A2(net1675),
    .A3(\core.registers[30][19] ),
    .B1(net1708),
    .X(_05921_));
 sky130_fd_sc_hd__a211o_1 _10934_ (.A1(net1699),
    .A2(_05919_),
    .B1(_05920_),
    .C1(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__o211a_1 _10935_ (.A1(net1753),
    .A2(_05918_),
    .B1(_05922_),
    .C1(net1763),
    .X(_05923_));
 sky130_fd_sc_hd__or2_1 _10936_ (.A(\core.registers[9][19] ),
    .B(net1357),
    .X(_05924_));
 sky130_fd_sc_hd__o211a_1 _10937_ (.A1(\core.registers[8][19] ),
    .A2(net1366),
    .B1(net1329),
    .C1(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__a22o_1 _10938_ (.A1(net1678),
    .A2(\core.registers[10][19] ),
    .B1(\core.registers[11][19] ),
    .B2(net1370),
    .X(_05926_));
 sky130_fd_sc_hd__a21o_1 _10939_ (.A1(net1342),
    .A2(_05926_),
    .B1(net1753),
    .X(_05927_));
 sky130_fd_sc_hd__mux2_1 _10940_ (.A0(\core.registers[24][19] ),
    .A1(\core.registers[25][19] ),
    .S(net1366),
    .X(_05928_));
 sky130_fd_sc_hd__a22o_1 _10941_ (.A1(net1676),
    .A2(\core.registers[26][19] ),
    .B1(\core.registers[27][19] ),
    .B2(net1366),
    .X(_05929_));
 sky130_fd_sc_hd__mux2_1 _10942_ (.A0(_05928_),
    .A1(_05929_),
    .S(net1768),
    .X(_05930_));
 sky130_fd_sc_hd__o221a_1 _10943_ (.A1(_05925_),
    .A2(_05927_),
    .B1(_05930_),
    .B2(net1708),
    .C1(net1704),
    .X(_05931_));
 sky130_fd_sc_hd__a21o_1 _10944_ (.A1(_05905_),
    .A2(_05908_),
    .B1(net1429),
    .X(_05932_));
 sky130_fd_sc_hd__a21o_1 _10945_ (.A1(_05912_),
    .A2(_05915_),
    .B1(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__o31a_2 _10946_ (.A1(net1427),
    .A2(_05923_),
    .A3(_05931_),
    .B1(_05933_),
    .X(_05934_));
 sky130_fd_sc_hd__o21a_1 _10947_ (.A1(net1141),
    .A2(net845),
    .B1(net1239),
    .X(_05935_));
 sky130_fd_sc_hd__o21ai_1 _10948_ (.A1(net1148),
    .A2(_05934_),
    .B1(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__nor2_1 _10949_ (.A(net1039),
    .B(_05936_),
    .Y(_05937_));
 sky130_fd_sc_hd__o22a_1 _10950_ (.A1(net1780),
    .A2(net1252),
    .B1(net1005),
    .B2(_05937_),
    .X(_05938_));
 sky130_fd_sc_hd__mux4_1 _10951_ (.A0(\core.registers[8][19] ),
    .A1(\core.registers[9][19] ),
    .A2(\core.registers[12][19] ),
    .A3(\core.registers[13][19] ),
    .S0(net1465),
    .S1(net1582),
    .X(_05939_));
 sky130_fd_sc_hd__nand2_1 _10952_ (.A(net1526),
    .B(_05939_),
    .Y(_05940_));
 sky130_fd_sc_hd__a22o_1 _10953_ (.A1(net1643),
    .A2(\core.registers[14][19] ),
    .B1(\core.registers[15][19] ),
    .B2(net1465),
    .X(_05941_));
 sky130_fd_sc_hd__a22o_1 _10954_ (.A1(net1643),
    .A2(\core.registers[10][19] ),
    .B1(\core.registers[11][19] ),
    .B2(net1466),
    .X(_05942_));
 sky130_fd_sc_hd__mux2_1 _10955_ (.A0(_05941_),
    .A1(_05942_),
    .S(net1571),
    .X(_05943_));
 sky130_fd_sc_hd__a21oi_1 _10956_ (.A1(net1542),
    .A2(_05943_),
    .B1(net1561),
    .Y(_05944_));
 sky130_fd_sc_hd__mux4_1 _10957_ (.A0(\core.registers[0][19] ),
    .A1(\core.registers[1][19] ),
    .A2(\core.registers[4][19] ),
    .A3(\core.registers[5][19] ),
    .S0(net1478),
    .S1(net1583),
    .X(_05945_));
 sky130_fd_sc_hd__and2_1 _10958_ (.A(net1528),
    .B(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__a22o_1 _10959_ (.A1(net1644),
    .A2(\core.registers[6][19] ),
    .B1(\core.registers[7][19] ),
    .B2(net1477),
    .X(_05947_));
 sky130_fd_sc_hd__a22o_1 _10960_ (.A1(net1643),
    .A2(\core.registers[2][19] ),
    .B1(\core.registers[3][19] ),
    .B2(net1477),
    .X(_05948_));
 sky130_fd_sc_hd__mux2_1 _10961_ (.A0(_05947_),
    .A1(_05948_),
    .S(net1572),
    .X(_05949_));
 sky130_fd_sc_hd__a21o_1 _10962_ (.A1(net1546),
    .A2(_05949_),
    .B1(net1566),
    .X(_05950_));
 sky130_fd_sc_hd__nor2_1 _10963_ (.A(_05946_),
    .B(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__a22o_1 _10964_ (.A1(net1641),
    .A2(\core.registers[30][19] ),
    .B1(\core.registers[31][19] ),
    .B2(net1465),
    .X(_05952_));
 sky130_fd_sc_hd__a22o_1 _10965_ (.A1(net1642),
    .A2(\core.registers[26][19] ),
    .B1(\core.registers[27][19] ),
    .B2(net1465),
    .X(_05953_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(_05952_),
    .A1(_05953_),
    .S(net1571),
    .X(_05954_));
 sky130_fd_sc_hd__mux4_1 _10967_ (.A0(\core.registers[24][19] ),
    .A1(\core.registers[25][19] ),
    .A2(\core.registers[28][19] ),
    .A3(\core.registers[29][19] ),
    .S0(net1465),
    .S1(net1582),
    .X(_05955_));
 sky130_fd_sc_hd__a21o_1 _10968_ (.A1(net1526),
    .A2(_05955_),
    .B1(net1561),
    .X(_05956_));
 sky130_fd_sc_hd__a21oi_1 _10969_ (.A1(net1542),
    .A2(_05954_),
    .B1(_05956_),
    .Y(_05957_));
 sky130_fd_sc_hd__mux4_1 _10970_ (.A0(\core.registers[16][19] ),
    .A1(\core.registers[17][19] ),
    .A2(\core.registers[20][19] ),
    .A3(\core.registers[21][19] ),
    .S0(net1465),
    .S1(net1582),
    .X(_05958_));
 sky130_fd_sc_hd__a22o_1 _10971_ (.A1(net1641),
    .A2(\core.registers[22][19] ),
    .B1(\core.registers[23][19] ),
    .B2(net1465),
    .X(_05959_));
 sky130_fd_sc_hd__a22o_1 _10972_ (.A1(net1641),
    .A2(\core.registers[18][19] ),
    .B1(\core.registers[19][19] ),
    .B2(net1465),
    .X(_05960_));
 sky130_fd_sc_hd__mux2_1 _10973_ (.A0(_05959_),
    .A1(_05960_),
    .S(net1571),
    .X(_05961_));
 sky130_fd_sc_hd__a21o_1 _10974_ (.A1(net1542),
    .A2(_05961_),
    .B1(net1566),
    .X(_05962_));
 sky130_fd_sc_hd__a21oi_1 _10975_ (.A1(net1526),
    .A2(_05958_),
    .B1(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__a21o_1 _10976_ (.A1(_05940_),
    .A2(_05944_),
    .B1(net1597),
    .X(_05964_));
 sky130_fd_sc_hd__or3_1 _10977_ (.A(net1593),
    .B(_05957_),
    .C(_05963_),
    .X(_05965_));
 sky130_fd_sc_hd__o21a_2 _10978_ (.A1(_05951_),
    .A2(_05964_),
    .B1(_05965_),
    .X(_05966_));
 sky130_fd_sc_hd__o2bb2a_2 _10979_ (.A1_N(net1094),
    .A2_N(net845),
    .B1(_05966_),
    .B2(net1045),
    .X(_05967_));
 sky130_fd_sc_hd__inv_2 _10980_ (.A(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__mux2_2 _10981_ (.A0(net460),
    .A1(_05968_),
    .S(net1252),
    .X(_05969_));
 sky130_fd_sc_hd__inv_2 _10982_ (.A(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__and2_1 _10983_ (.A(_05938_),
    .B(_05969_),
    .X(_05971_));
 sky130_fd_sc_hd__inv_2 _10984_ (.A(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__or2_4 _10985_ (.A(_05938_),
    .B(_05969_),
    .X(_05973_));
 sky130_fd_sc_hd__a21oi_1 _10986_ (.A1(net1618),
    .A2(_04139_),
    .B1(net1186),
    .Y(_05974_));
 sky130_fd_sc_hd__a21oi_1 _10987_ (.A1(\core.pipe1_csrData[18] ),
    .A2(net1250),
    .B1(net1237),
    .Y(_05975_));
 sky130_fd_sc_hd__nor2_1 _10988_ (.A(_05974_),
    .B(_05975_),
    .Y(_05976_));
 sky130_fd_sc_hd__o22a_4 _10989_ (.A1(\core.pipe1_resultRegister[18] ),
    .A2(net1188),
    .B1(_05976_),
    .B2(net1245),
    .X(_05977_));
 sky130_fd_sc_hd__or2_1 _10990_ (.A(\core.registers[5][18] ),
    .B(net1360),
    .X(_05978_));
 sky130_fd_sc_hd__o211a_1 _10991_ (.A1(\core.registers[4][18] ),
    .A2(net1420),
    .B1(_05978_),
    .C1(net1455),
    .X(_05979_));
 sky130_fd_sc_hd__mux2_1 _10992_ (.A0(\core.registers[0][18] ),
    .A1(\core.registers[1][18] ),
    .S(net1420),
    .X(_05980_));
 sky130_fd_sc_hd__a211o_1 _10993_ (.A1(net1444),
    .A2(_05980_),
    .B1(_05979_),
    .C1(net1352),
    .X(_05981_));
 sky130_fd_sc_hd__o221a_1 _10994_ (.A1(net1692),
    .A2(\core.registers[7][18] ),
    .B1(net1420),
    .B2(\core.registers[6][18] ),
    .C1(net1455),
    .X(_05982_));
 sky130_fd_sc_hd__o221a_1 _10995_ (.A1(net1692),
    .A2(\core.registers[3][18] ),
    .B1(net1420),
    .B2(\core.registers[2][18] ),
    .C1(net1444),
    .X(_05983_));
 sky130_fd_sc_hd__o31a_1 _10996_ (.A1(net1337),
    .A2(_05982_),
    .A3(_05983_),
    .B1(net1323),
    .X(_05984_));
 sky130_fd_sc_hd__or2_1 _10997_ (.A(\core.registers[16][18] ),
    .B(net1420),
    .X(_05985_));
 sky130_fd_sc_hd__o211a_1 _10998_ (.A1(\core.registers[17][18] ),
    .A2(net1360),
    .B1(_05985_),
    .C1(net1446),
    .X(_05986_));
 sky130_fd_sc_hd__mux2_1 _10999_ (.A0(\core.registers[20][18] ),
    .A1(\core.registers[21][18] ),
    .S(net1420),
    .X(_05987_));
 sky130_fd_sc_hd__a211o_1 _11000_ (.A1(net1454),
    .A2(_05987_),
    .B1(_05986_),
    .C1(net1352),
    .X(_05988_));
 sky130_fd_sc_hd__o221a_1 _11001_ (.A1(net1692),
    .A2(\core.registers[23][18] ),
    .B1(net1420),
    .B2(\core.registers[22][18] ),
    .C1(net1454),
    .X(_05989_));
 sky130_fd_sc_hd__o221a_1 _11002_ (.A1(net1693),
    .A2(\core.registers[19][18] ),
    .B1(net1420),
    .B2(\core.registers[18][18] ),
    .C1(net1446),
    .X(_05990_));
 sky130_fd_sc_hd__o31a_1 _11003_ (.A1(net1337),
    .A2(_05989_),
    .A3(_05990_),
    .B1(net1326),
    .X(_05991_));
 sky130_fd_sc_hd__mux2_1 _11004_ (.A0(\core.registers[12][18] ),
    .A1(\core.registers[13][18] ),
    .S(net1421),
    .X(_05992_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(\core.registers[14][18] ),
    .A1(\core.registers[15][18] ),
    .S(net1421),
    .X(_05993_));
 sky130_fd_sc_hd__mux2_1 _11006_ (.A0(_05992_),
    .A1(_05993_),
    .S(net1352),
    .X(_05994_));
 sky130_fd_sc_hd__mux2_1 _11007_ (.A0(\core.registers[28][18] ),
    .A1(\core.registers[29][18] ),
    .S(net1416),
    .X(_05995_));
 sky130_fd_sc_hd__and3_1 _11008_ (.A(net1774),
    .B(\core.registers[31][18] ),
    .C(net1416),
    .X(_05996_));
 sky130_fd_sc_hd__a31o_1 _11009_ (.A1(net1774),
    .A2(net1691),
    .A3(\core.registers[30][18] ),
    .B1(net1710),
    .X(_05997_));
 sky130_fd_sc_hd__a211o_1 _11010_ (.A1(net1701),
    .A2(_05995_),
    .B1(_05996_),
    .C1(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__o211a_1 _11011_ (.A1(net1759),
    .A2(_05994_),
    .B1(_05998_),
    .C1(net1766),
    .X(_05999_));
 sky130_fd_sc_hd__or2_1 _11012_ (.A(\core.registers[9][18] ),
    .B(net1360),
    .X(_06000_));
 sky130_fd_sc_hd__o211a_1 _11013_ (.A1(\core.registers[8][18] ),
    .A2(net1416),
    .B1(net1337),
    .C1(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__a22o_1 _11014_ (.A1(net1692),
    .A2(\core.registers[10][18] ),
    .B1(\core.registers[11][18] ),
    .B2(net1421),
    .X(_06002_));
 sky130_fd_sc_hd__a21o_1 _11015_ (.A1(net1352),
    .A2(_06002_),
    .B1(net1759),
    .X(_06003_));
 sky130_fd_sc_hd__mux2_1 _11016_ (.A0(\core.registers[24][18] ),
    .A1(\core.registers[25][18] ),
    .S(net1416),
    .X(_06004_));
 sky130_fd_sc_hd__a22o_1 _11017_ (.A1(net1691),
    .A2(\core.registers[26][18] ),
    .B1(\core.registers[27][18] ),
    .B2(net1417),
    .X(_06005_));
 sky130_fd_sc_hd__mux2_1 _11018_ (.A0(_06004_),
    .A1(_06005_),
    .S(net1774),
    .X(_06006_));
 sky130_fd_sc_hd__o221a_1 _11019_ (.A1(_06001_),
    .A2(_06003_),
    .B1(_06006_),
    .B2(net1710),
    .C1(net1706),
    .X(_06007_));
 sky130_fd_sc_hd__a21o_1 _11020_ (.A1(_05981_),
    .A2(_05984_),
    .B1(net1433),
    .X(_06008_));
 sky130_fd_sc_hd__a21o_1 _11021_ (.A1(_05988_),
    .A2(_05991_),
    .B1(_06008_),
    .X(_06009_));
 sky130_fd_sc_hd__o31a_4 _11022_ (.A1(_04077_),
    .A2(_05999_),
    .A3(_06007_),
    .B1(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__o21a_1 _11023_ (.A1(net1144),
    .A2(net841),
    .B1(net1241),
    .X(_06011_));
 sky130_fd_sc_hd__o21ai_4 _11024_ (.A1(net1149),
    .A2(_06010_),
    .B1(_06011_),
    .Y(_06012_));
 sky130_fd_sc_hd__nor2_1 _11025_ (.A(net1039),
    .B(_06012_),
    .Y(_06013_));
 sky130_fd_sc_hd__o22a_2 _11026_ (.A1(\core.pipe0_currentInstruction[18] ),
    .A2(net1252),
    .B1(net1005),
    .B2(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__mux4_1 _11027_ (.A0(\core.registers[8][18] ),
    .A1(\core.registers[9][18] ),
    .A2(\core.registers[12][18] ),
    .A3(\core.registers[13][18] ),
    .S0(net1520),
    .S1(net1590),
    .X(_06015_));
 sky130_fd_sc_hd__nand2_1 _11028_ (.A(net1538),
    .B(_06015_),
    .Y(_06016_));
 sky130_fd_sc_hd__a22o_1 _11029_ (.A1(net1658),
    .A2(\core.registers[14][18] ),
    .B1(\core.registers[15][18] ),
    .B2(net1520),
    .X(_06017_));
 sky130_fd_sc_hd__a22o_1 _11030_ (.A1(net1658),
    .A2(\core.registers[10][18] ),
    .B1(\core.registers[11][18] ),
    .B2(net1520),
    .X(_06018_));
 sky130_fd_sc_hd__mux2_1 _11031_ (.A0(_06017_),
    .A1(_06018_),
    .S(net1578),
    .X(_06019_));
 sky130_fd_sc_hd__a21oi_1 _11032_ (.A1(net1557),
    .A2(_06019_),
    .B1(net1564),
    .Y(_06020_));
 sky130_fd_sc_hd__mux4_1 _11033_ (.A0(\core.registers[0][18] ),
    .A1(\core.registers[1][18] ),
    .A2(\core.registers[4][18] ),
    .A3(\core.registers[5][18] ),
    .S0(net1519),
    .S1(net1590),
    .X(_06021_));
 sky130_fd_sc_hd__and2_1 _11034_ (.A(net1538),
    .B(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__a22o_1 _11035_ (.A1(net1660),
    .A2(\core.registers[6][18] ),
    .B1(\core.registers[7][18] ),
    .B2(net1519),
    .X(_06023_));
 sky130_fd_sc_hd__a22o_1 _11036_ (.A1(net1658),
    .A2(\core.registers[2][18] ),
    .B1(\core.registers[3][18] ),
    .B2(net1519),
    .X(_06024_));
 sky130_fd_sc_hd__mux2_1 _11037_ (.A0(_06023_),
    .A1(_06024_),
    .S(net1578),
    .X(_06025_));
 sky130_fd_sc_hd__a21o_1 _11038_ (.A1(net1557),
    .A2(_06025_),
    .B1(net1570),
    .X(_06026_));
 sky130_fd_sc_hd__nor2_1 _11039_ (.A(_06022_),
    .B(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__a22o_1 _11040_ (.A1(net1661),
    .A2(\core.registers[30][18] ),
    .B1(\core.registers[31][18] ),
    .B2(net1515),
    .X(_06028_));
 sky130_fd_sc_hd__a22o_1 _11041_ (.A1(net1661),
    .A2(\core.registers[26][18] ),
    .B1(\core.registers[27][18] ),
    .B2(net1515),
    .X(_06029_));
 sky130_fd_sc_hd__mux2_1 _11042_ (.A0(_06028_),
    .A1(_06029_),
    .S(net1579),
    .X(_06030_));
 sky130_fd_sc_hd__mux4_1 _11043_ (.A0(\core.registers[24][18] ),
    .A1(\core.registers[25][18] ),
    .A2(\core.registers[28][18] ),
    .A3(\core.registers[29][18] ),
    .S0(net1516),
    .S1(net1591),
    .X(_06031_));
 sky130_fd_sc_hd__a21o_1 _11044_ (.A1(net1540),
    .A2(_06031_),
    .B1(net1564),
    .X(_06032_));
 sky130_fd_sc_hd__a21oi_1 _11045_ (.A1(net1559),
    .A2(_06030_),
    .B1(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__mux4_1 _11046_ (.A0(\core.registers[16][18] ),
    .A1(\core.registers[17][18] ),
    .A2(\core.registers[20][18] ),
    .A3(\core.registers[21][18] ),
    .S0(net1519),
    .S1(net1589),
    .X(_06034_));
 sky130_fd_sc_hd__a22o_1 _11047_ (.A1(net1658),
    .A2(\core.registers[22][18] ),
    .B1(\core.registers[23][18] ),
    .B2(net1519),
    .X(_06035_));
 sky130_fd_sc_hd__a22o_1 _11048_ (.A1(net1658),
    .A2(\core.registers[18][18] ),
    .B1(\core.registers[19][18] ),
    .B2(net1519),
    .X(_06036_));
 sky130_fd_sc_hd__mux2_1 _11049_ (.A0(_06035_),
    .A1(_06036_),
    .S(net1578),
    .X(_06037_));
 sky130_fd_sc_hd__a21o_1 _11050_ (.A1(net1557),
    .A2(_06037_),
    .B1(net1568),
    .X(_06038_));
 sky130_fd_sc_hd__a21oi_1 _11051_ (.A1(net1538),
    .A2(_06034_),
    .B1(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__a21o_1 _11052_ (.A1(_06016_),
    .A2(_06020_),
    .B1(net1599),
    .X(_06040_));
 sky130_fd_sc_hd__or3_1 _11053_ (.A(net1595),
    .B(_06033_),
    .C(_06039_),
    .X(_06041_));
 sky130_fd_sc_hd__o21a_4 _11054_ (.A1(_06027_),
    .A2(_06040_),
    .B1(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__o2bb2a_4 _11055_ (.A1_N(net1095),
    .A2_N(net841),
    .B1(_06042_),
    .B2(net1044),
    .X(_06043_));
 sky130_fd_sc_hd__inv_2 _11056_ (.A(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__mux2_4 _11057_ (.A0(net459),
    .A1(_06044_),
    .S(net1253),
    .X(_06045_));
 sky130_fd_sc_hd__inv_2 _11058_ (.A(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__and2_4 _11059_ (.A(_06014_),
    .B(_06045_),
    .X(_06047_));
 sky130_fd_sc_hd__clkinv_2 _11060_ (.A(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__nor2_4 _11061_ (.A(_06014_),
    .B(_06045_),
    .Y(_06049_));
 sky130_fd_sc_hd__nor2_8 _11062_ (.A(_06047_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__inv_2 _11063_ (.A(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__a21oi_1 _11064_ (.A1(net1618),
    .A2(_04227_),
    .B1(net1187),
    .Y(_06052_));
 sky130_fd_sc_hd__a21oi_1 _11065_ (.A1(\core.pipe1_csrData[17] ),
    .A2(net1249),
    .B1(net1238),
    .Y(_06053_));
 sky130_fd_sc_hd__nor2_1 _11066_ (.A(_06052_),
    .B(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__o22a_4 _11067_ (.A1(\core.pipe1_resultRegister[17] ),
    .A2(net1188),
    .B1(_06054_),
    .B2(net1246),
    .X(_06055_));
 sky130_fd_sc_hd__or2_1 _11068_ (.A(\core.registers[5][17] ),
    .B(net1357),
    .X(_06056_));
 sky130_fd_sc_hd__o211a_1 _11069_ (.A1(\core.registers[4][17] ),
    .A2(net1380),
    .B1(_06056_),
    .C1(net1448),
    .X(_06057_));
 sky130_fd_sc_hd__mux2_1 _11070_ (.A0(\core.registers[0][17] ),
    .A1(\core.registers[1][17] ),
    .S(net1380),
    .X(_06058_));
 sky130_fd_sc_hd__a211o_1 _11071_ (.A1(net1435),
    .A2(_06058_),
    .B1(_06057_),
    .C1(net1344),
    .X(_06059_));
 sky130_fd_sc_hd__o221a_1 _11072_ (.A1(net1680),
    .A2(\core.registers[7][17] ),
    .B1(net1378),
    .B2(\core.registers[6][17] ),
    .C1(net1448),
    .X(_06060_));
 sky130_fd_sc_hd__o221a_1 _11073_ (.A1(net1680),
    .A2(\core.registers[3][17] ),
    .B1(net1381),
    .B2(\core.registers[2][17] ),
    .C1(net1435),
    .X(_06061_));
 sky130_fd_sc_hd__o31a_1 _11074_ (.A1(net1330),
    .A2(_06060_),
    .A3(_06061_),
    .B1(net1320),
    .X(_06062_));
 sky130_fd_sc_hd__or2_1 _11075_ (.A(\core.registers[16][17] ),
    .B(net1378),
    .X(_06063_));
 sky130_fd_sc_hd__o211a_1 _11076_ (.A1(\core.registers[17][17] ),
    .A2(net1357),
    .B1(_06063_),
    .C1(net1435),
    .X(_06064_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(\core.registers[20][17] ),
    .A1(\core.registers[21][17] ),
    .S(net1378),
    .X(_06065_));
 sky130_fd_sc_hd__a211o_1 _11078_ (.A1(net1448),
    .A2(_06065_),
    .B1(_06064_),
    .C1(net1344),
    .X(_06066_));
 sky130_fd_sc_hd__o221a_1 _11079_ (.A1(net1678),
    .A2(\core.registers[23][17] ),
    .B1(net1367),
    .B2(\core.registers[22][17] ),
    .C1(net1447),
    .X(_06067_));
 sky130_fd_sc_hd__o221a_1 _11080_ (.A1(net1678),
    .A2(\core.registers[19][17] ),
    .B1(net1367),
    .B2(\core.registers[18][17] ),
    .C1(net1434),
    .X(_06068_));
 sky130_fd_sc_hd__o31a_1 _11081_ (.A1(net1329),
    .A2(_06067_),
    .A3(_06068_),
    .B1(net1324),
    .X(_06069_));
 sky130_fd_sc_hd__mux2_1 _11082_ (.A0(\core.registers[12][17] ),
    .A1(\core.registers[13][17] ),
    .S(net1367),
    .X(_06070_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(\core.registers[14][17] ),
    .A1(\core.registers[15][17] ),
    .S(net1378),
    .X(_06071_));
 sky130_fd_sc_hd__mux2_1 _11084_ (.A0(_06070_),
    .A1(_06071_),
    .S(net1344),
    .X(_06072_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(\core.registers[28][17] ),
    .A1(\core.registers[29][17] ),
    .S(net1378),
    .X(_06073_));
 sky130_fd_sc_hd__and3_1 _11086_ (.A(net1770),
    .B(\core.registers[31][17] ),
    .C(net1378),
    .X(_06074_));
 sky130_fd_sc_hd__a211o_1 _11087_ (.A1(\core.registers[30][17] ),
    .A2(net1319),
    .B1(_06074_),
    .C1(net1708),
    .X(_06075_));
 sky130_fd_sc_hd__a21o_1 _11088_ (.A1(net1703),
    .A2(_06073_),
    .B1(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__o211a_1 _11089_ (.A1(net1754),
    .A2(_06072_),
    .B1(_06076_),
    .C1(net1763),
    .X(_06077_));
 sky130_fd_sc_hd__or2_1 _11090_ (.A(\core.registers[9][17] ),
    .B(net1357),
    .X(_06078_));
 sky130_fd_sc_hd__o211a_1 _11091_ (.A1(\core.registers[8][17] ),
    .A2(net1370),
    .B1(net1328),
    .C1(_06078_),
    .X(_06079_));
 sky130_fd_sc_hd__a22o_1 _11092_ (.A1(net1678),
    .A2(\core.registers[10][17] ),
    .B1(\core.registers[11][17] ),
    .B2(net1367),
    .X(_06080_));
 sky130_fd_sc_hd__a21o_1 _11093_ (.A1(net1342),
    .A2(_06080_),
    .B1(net1754),
    .X(_06081_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(\core.registers[24][17] ),
    .A1(\core.registers[25][17] ),
    .S(net1378),
    .X(_06082_));
 sky130_fd_sc_hd__a22o_1 _11095_ (.A1(net1678),
    .A2(\core.registers[26][17] ),
    .B1(\core.registers[27][17] ),
    .B2(net1378),
    .X(_06083_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(_06082_),
    .A1(_06083_),
    .S(net1770),
    .X(_06084_));
 sky130_fd_sc_hd__o221a_1 _11097_ (.A1(_06079_),
    .A2(_06081_),
    .B1(_06084_),
    .B2(net1708),
    .C1(net1704),
    .X(_06085_));
 sky130_fd_sc_hd__a21o_1 _11098_ (.A1(_06059_),
    .A2(_06062_),
    .B1(net1429),
    .X(_06086_));
 sky130_fd_sc_hd__a21o_1 _11099_ (.A1(_06066_),
    .A2(_06069_),
    .B1(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__o31a_2 _11100_ (.A1(net1427),
    .A2(_06077_),
    .A3(_06085_),
    .B1(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__o21a_1 _11101_ (.A1(net1141),
    .A2(_06055_),
    .B1(net1239),
    .X(_06089_));
 sky130_fd_sc_hd__o21ai_2 _11102_ (.A1(net1148),
    .A2(_06088_),
    .B1(_06089_),
    .Y(_06090_));
 sky130_fd_sc_hd__nor2_1 _11103_ (.A(net1039),
    .B(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__o22a_2 _11104_ (.A1(net1784),
    .A2(net1252),
    .B1(net1005),
    .B2(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__mux4_1 _11105_ (.A0(\core.registers[8][17] ),
    .A1(\core.registers[9][17] ),
    .A2(\core.registers[12][17] ),
    .A3(\core.registers[13][17] ),
    .S0(net1466),
    .S1(net1583),
    .X(_06093_));
 sky130_fd_sc_hd__nand2_1 _11106_ (.A(net1528),
    .B(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__a22o_1 _11107_ (.A1(net1643),
    .A2(\core.registers[14][17] ),
    .B1(\core.registers[15][17] ),
    .B2(net1477),
    .X(_06095_));
 sky130_fd_sc_hd__a22o_1 _11108_ (.A1(net1643),
    .A2(\core.registers[10][17] ),
    .B1(\core.registers[11][17] ),
    .B2(net1466),
    .X(_06096_));
 sky130_fd_sc_hd__mux2_1 _11109_ (.A0(_06095_),
    .A1(_06096_),
    .S(net1572),
    .X(_06097_));
 sky130_fd_sc_hd__a21oi_1 _11110_ (.A1(net1542),
    .A2(_06097_),
    .B1(net1561),
    .Y(_06098_));
 sky130_fd_sc_hd__mux4_1 _11111_ (.A0(\core.registers[0][17] ),
    .A1(\core.registers[1][17] ),
    .A2(\core.registers[4][17] ),
    .A3(\core.registers[5][17] ),
    .S0(net1479),
    .S1(net1585),
    .X(_06099_));
 sky130_fd_sc_hd__and2_1 _11112_ (.A(net1527),
    .B(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__a22o_1 _11113_ (.A1(net1647),
    .A2(\core.registers[6][17] ),
    .B1(\core.registers[7][17] ),
    .B2(net1477),
    .X(_06101_));
 sky130_fd_sc_hd__a22o_1 _11114_ (.A1(net1647),
    .A2(\core.registers[2][17] ),
    .B1(\core.registers[3][17] ),
    .B2(net1480),
    .X(_06102_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(_06101_),
    .A1(_06102_),
    .S(net1572),
    .X(_06103_));
 sky130_fd_sc_hd__a21o_1 _11116_ (.A1(net1546),
    .A2(_06103_),
    .B1(net1566),
    .X(_06104_));
 sky130_fd_sc_hd__nor2_1 _11117_ (.A(_06100_),
    .B(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__a22o_1 _11118_ (.A1(net1643),
    .A2(\core.registers[30][17] ),
    .B1(\core.registers[31][17] ),
    .B2(net1477),
    .X(_06106_));
 sky130_fd_sc_hd__a22o_1 _11119_ (.A1(net1643),
    .A2(\core.registers[26][17] ),
    .B1(\core.registers[27][17] ),
    .B2(net1477),
    .X(_06107_));
 sky130_fd_sc_hd__mux2_1 _11120_ (.A0(_06106_),
    .A1(_06107_),
    .S(net1572),
    .X(_06108_));
 sky130_fd_sc_hd__mux4_1 _11121_ (.A0(\core.registers[24][17] ),
    .A1(\core.registers[25][17] ),
    .A2(\core.registers[28][17] ),
    .A3(\core.registers[29][17] ),
    .S0(net1477),
    .S1(net1583),
    .X(_06109_));
 sky130_fd_sc_hd__a21o_1 _11122_ (.A1(net1527),
    .A2(_06109_),
    .B1(net1561),
    .X(_06110_));
 sky130_fd_sc_hd__a21oi_1 _11123_ (.A1(net1546),
    .A2(_06108_),
    .B1(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__mux4_1 _11124_ (.A0(\core.registers[16][17] ),
    .A1(\core.registers[17][17] ),
    .A2(\core.registers[20][17] ),
    .A3(\core.registers[21][17] ),
    .S0(net1477),
    .S1(net1583),
    .X(_06112_));
 sky130_fd_sc_hd__a22o_1 _11125_ (.A1(net1643),
    .A2(\core.registers[22][17] ),
    .B1(\core.registers[23][17] ),
    .B2(net1477),
    .X(_06113_));
 sky130_fd_sc_hd__a22o_1 _11126_ (.A1(net1643),
    .A2(\core.registers[18][17] ),
    .B1(\core.registers[19][17] ),
    .B2(net1466),
    .X(_06114_));
 sky130_fd_sc_hd__mux2_1 _11127_ (.A0(_06113_),
    .A1(_06114_),
    .S(net1572),
    .X(_06115_));
 sky130_fd_sc_hd__a21o_1 _11128_ (.A1(net1546),
    .A2(_06115_),
    .B1(net1566),
    .X(_06116_));
 sky130_fd_sc_hd__a21oi_1 _11129_ (.A1(net1527),
    .A2(_06112_),
    .B1(_06116_),
    .Y(_06117_));
 sky130_fd_sc_hd__a21o_1 _11130_ (.A1(_06094_),
    .A2(_06098_),
    .B1(net1597),
    .X(_06118_));
 sky130_fd_sc_hd__or3_1 _11131_ (.A(net1593),
    .B(_06111_),
    .C(_06117_),
    .X(_06119_));
 sky130_fd_sc_hd__o21a_2 _11132_ (.A1(_06105_),
    .A2(_06118_),
    .B1(_06119_),
    .X(_06120_));
 sky130_fd_sc_hd__o2bb2a_2 _11133_ (.A1_N(net1094),
    .A2_N(_06055_),
    .B1(_06120_),
    .B2(net1045),
    .X(_06121_));
 sky130_fd_sc_hd__inv_2 _11134_ (.A(_06121_),
    .Y(_06122_));
 sky130_fd_sc_hd__mux2_2 _11135_ (.A0(net458),
    .A1(_06122_),
    .S(net1252),
    .X(_06123_));
 sky130_fd_sc_hd__clkinv_2 _11136_ (.A(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__and2_4 _11137_ (.A(_06092_),
    .B(_06123_),
    .X(_06125_));
 sky130_fd_sc_hd__nor2_2 _11138_ (.A(_06092_),
    .B(_06123_),
    .Y(_06126_));
 sky130_fd_sc_hd__nor2_4 _11139_ (.A(_06125_),
    .B(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__inv_2 _11140_ (.A(_06127_),
    .Y(_06128_));
 sky130_fd_sc_hd__nor2_1 _11141_ (.A(_04002_),
    .B(_04314_),
    .Y(_06129_));
 sky130_fd_sc_hd__a21o_1 _11142_ (.A1(\core.pipe1_csrData[16] ),
    .A2(net1249),
    .B1(net1238),
    .X(_06130_));
 sky130_fd_sc_hd__o21a_1 _11143_ (.A1(net1186),
    .A2(_06129_),
    .B1(_06130_),
    .X(_06131_));
 sky130_fd_sc_hd__o22a_4 _11144_ (.A1(\core.pipe1_resultRegister[16] ),
    .A2(net1189),
    .B1(_06131_),
    .B2(net1246),
    .X(_06132_));
 sky130_fd_sc_hd__or2_1 _11145_ (.A(\core.registers[5][16] ),
    .B(net1359),
    .X(_06133_));
 sky130_fd_sc_hd__o211a_1 _11146_ (.A1(\core.registers[4][16] ),
    .A2(net1388),
    .B1(_06133_),
    .C1(net1451),
    .X(_06134_));
 sky130_fd_sc_hd__mux2_1 _11147_ (.A0(\core.registers[0][16] ),
    .A1(\core.registers[1][16] ),
    .S(net1388),
    .X(_06135_));
 sky130_fd_sc_hd__a211o_1 _11148_ (.A1(net1438),
    .A2(_06135_),
    .B1(_06134_),
    .C1(net1349),
    .X(_06136_));
 sky130_fd_sc_hd__o221a_1 _11149_ (.A1(net1686),
    .A2(\core.registers[7][16] ),
    .B1(net1401),
    .B2(\core.registers[6][16] ),
    .C1(net1451),
    .X(_06137_));
 sky130_fd_sc_hd__o221a_1 _11150_ (.A1(net1683),
    .A2(\core.registers[3][16] ),
    .B1(net1401),
    .B2(\core.registers[2][16] ),
    .C1(net1440),
    .X(_06138_));
 sky130_fd_sc_hd__o31a_1 _11151_ (.A1(net1333),
    .A2(_06137_),
    .A3(_06138_),
    .B1(net1321),
    .X(_06139_));
 sky130_fd_sc_hd__or2_1 _11152_ (.A(\core.registers[16][16] ),
    .B(net1384),
    .X(_06140_));
 sky130_fd_sc_hd__o211a_1 _11153_ (.A1(\core.registers[17][16] ),
    .A2(net1359),
    .B1(_06140_),
    .C1(net1439),
    .X(_06141_));
 sky130_fd_sc_hd__mux2_1 _11154_ (.A0(\core.registers[20][16] ),
    .A1(\core.registers[21][16] ),
    .S(net1385),
    .X(_06142_));
 sky130_fd_sc_hd__a211o_1 _11155_ (.A1(net1451),
    .A2(_06142_),
    .B1(_06141_),
    .C1(net1347),
    .X(_06143_));
 sky130_fd_sc_hd__o221a_1 _11156_ (.A1(net1683),
    .A2(\core.registers[23][16] ),
    .B1(net1385),
    .B2(\core.registers[22][16] ),
    .C1(net1451),
    .X(_06144_));
 sky130_fd_sc_hd__o221a_1 _11157_ (.A1(net1683),
    .A2(\core.registers[19][16] ),
    .B1(net1385),
    .B2(\core.registers[18][16] ),
    .C1(net1439),
    .X(_06145_));
 sky130_fd_sc_hd__o31a_1 _11158_ (.A1(net1331),
    .A2(_06144_),
    .A3(_06145_),
    .B1(net1325),
    .X(_06146_));
 sky130_fd_sc_hd__mux2_1 _11159_ (.A0(\core.registers[12][16] ),
    .A1(\core.registers[13][16] ),
    .S(net1393),
    .X(_06147_));
 sky130_fd_sc_hd__mux2_1 _11160_ (.A0(\core.registers[14][16] ),
    .A1(\core.registers[15][16] ),
    .S(net1401),
    .X(_06148_));
 sky130_fd_sc_hd__mux2_1 _11161_ (.A0(_06147_),
    .A1(_06148_),
    .S(net1347),
    .X(_06149_));
 sky130_fd_sc_hd__mux2_1 _11162_ (.A0(\core.registers[28][16] ),
    .A1(\core.registers[29][16] ),
    .S(net1393),
    .X(_06150_));
 sky130_fd_sc_hd__and3_1 _11163_ (.A(net1772),
    .B(\core.registers[31][16] ),
    .C(net1393),
    .X(_06151_));
 sky130_fd_sc_hd__a211o_1 _11164_ (.A1(\core.registers[30][16] ),
    .A2(net1319),
    .B1(_06151_),
    .C1(net1710),
    .X(_06152_));
 sky130_fd_sc_hd__a21o_1 _11165_ (.A1(net1702),
    .A2(_06150_),
    .B1(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__o211a_1 _11166_ (.A1(net1757),
    .A2(_06149_),
    .B1(_06153_),
    .C1(net1765),
    .X(_06154_));
 sky130_fd_sc_hd__or2_1 _11167_ (.A(\core.registers[9][16] ),
    .B(net1362),
    .X(_06155_));
 sky130_fd_sc_hd__o211a_1 _11168_ (.A1(\core.registers[8][16] ),
    .A2(net1393),
    .B1(net1333),
    .C1(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__a22o_1 _11169_ (.A1(net1686),
    .A2(\core.registers[10][16] ),
    .B1(\core.registers[11][16] ),
    .B2(net1401),
    .X(_06157_));
 sky130_fd_sc_hd__a21o_1 _11170_ (.A1(net1349),
    .A2(_06157_),
    .B1(net1757),
    .X(_06158_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(\core.registers[24][16] ),
    .A1(\core.registers[25][16] ),
    .S(net1393),
    .X(_06159_));
 sky130_fd_sc_hd__a22o_1 _11172_ (.A1(net1686),
    .A2(\core.registers[26][16] ),
    .B1(\core.registers[27][16] ),
    .B2(net1393),
    .X(_06160_));
 sky130_fd_sc_hd__mux2_1 _11173_ (.A0(_06159_),
    .A1(_06160_),
    .S(net1772),
    .X(_06161_));
 sky130_fd_sc_hd__o221a_1 _11174_ (.A1(_06156_),
    .A2(_06158_),
    .B1(_06161_),
    .B2(net1710),
    .C1(net1707),
    .X(_06162_));
 sky130_fd_sc_hd__a21o_1 _11175_ (.A1(_06136_),
    .A2(_06139_),
    .B1(net1431),
    .X(_06163_));
 sky130_fd_sc_hd__a21o_1 _11176_ (.A1(_06143_),
    .A2(_06146_),
    .B1(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__o31a_2 _11177_ (.A1(net1428),
    .A2(_06154_),
    .A3(_06162_),
    .B1(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__o21a_1 _11178_ (.A1(net1146),
    .A2(_06132_),
    .B1(net1240),
    .X(_06166_));
 sky130_fd_sc_hd__o21ai_4 _11179_ (.A1(net1148),
    .A2(_06165_),
    .B1(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__nor2_1 _11180_ (.A(net1040),
    .B(_06167_),
    .Y(_06168_));
 sky130_fd_sc_hd__o22a_4 _11181_ (.A1(net1789),
    .A2(net1253),
    .B1(net1005),
    .B2(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__mux4_1 _11182_ (.A0(\core.registers[8][16] ),
    .A1(\core.registers[9][16] ),
    .A2(\core.registers[12][16] ),
    .A3(\core.registers[13][16] ),
    .S0(net1492),
    .S1(net1587),
    .X(_06170_));
 sky130_fd_sc_hd__nand2_1 _11183_ (.A(net1532),
    .B(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__a22o_1 _11184_ (.A1(net1650),
    .A2(\core.registers[14][16] ),
    .B1(\core.registers[15][16] ),
    .B2(net1500),
    .X(_06172_));
 sky130_fd_sc_hd__a22o_1 _11185_ (.A1(net1653),
    .A2(\core.registers[10][16] ),
    .B1(\core.registers[11][16] ),
    .B2(net1500),
    .X(_06173_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(_06172_),
    .A1(_06173_),
    .S(net1575),
    .X(_06174_));
 sky130_fd_sc_hd__a21oi_1 _11187_ (.A1(net1552),
    .A2(_06174_),
    .B1(net1565),
    .Y(_06175_));
 sky130_fd_sc_hd__mux4_1 _11188_ (.A0(\core.registers[0][16] ),
    .A1(\core.registers[1][16] ),
    .A2(\core.registers[4][16] ),
    .A3(\core.registers[5][16] ),
    .S0(net1488),
    .S1(net1586),
    .X(_06176_));
 sky130_fd_sc_hd__and2_1 _11189_ (.A(net1532),
    .B(_06176_),
    .X(_06177_));
 sky130_fd_sc_hd__a22o_1 _11190_ (.A1(net1653),
    .A2(\core.registers[6][16] ),
    .B1(\core.registers[7][16] ),
    .B2(net1500),
    .X(_06178_));
 sky130_fd_sc_hd__a22o_1 _11191_ (.A1(net1650),
    .A2(\core.registers[2][16] ),
    .B1(\core.registers[3][16] ),
    .B2(net1500),
    .X(_06179_));
 sky130_fd_sc_hd__mux2_1 _11192_ (.A0(_06178_),
    .A1(_06179_),
    .S(net1575),
    .X(_06180_));
 sky130_fd_sc_hd__a21o_1 _11193_ (.A1(net1552),
    .A2(_06180_),
    .B1(net1570),
    .X(_06181_));
 sky130_fd_sc_hd__nor2_1 _11194_ (.A(_06177_),
    .B(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__a21oi_1 _11195_ (.A1(_06171_),
    .A2(_06175_),
    .B1(_06182_),
    .Y(_06183_));
 sky130_fd_sc_hd__a22o_1 _11196_ (.A1(net1648),
    .A2(\core.registers[30][16] ),
    .B1(\core.registers[31][16] ),
    .B2(net1492),
    .X(_06184_));
 sky130_fd_sc_hd__a22o_1 _11197_ (.A1(net1648),
    .A2(\core.registers[26][16] ),
    .B1(\core.registers[27][16] ),
    .B2(net1492),
    .X(_06185_));
 sky130_fd_sc_hd__mux2_1 _11198_ (.A0(_06184_),
    .A1(_06185_),
    .S(net1575),
    .X(_06186_));
 sky130_fd_sc_hd__mux4_1 _11199_ (.A0(\core.registers[24][16] ),
    .A1(\core.registers[25][16] ),
    .A2(\core.registers[28][16] ),
    .A3(\core.registers[29][16] ),
    .S0(net1492),
    .S1(net1587),
    .X(_06187_));
 sky130_fd_sc_hd__a21o_1 _11200_ (.A1(net1533),
    .A2(_06187_),
    .B1(net1563),
    .X(_06188_));
 sky130_fd_sc_hd__a21o_1 _11201_ (.A1(net1551),
    .A2(_06186_),
    .B1(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__mux4_1 _11202_ (.A0(\core.registers[16][16] ),
    .A1(\core.registers[17][16] ),
    .A2(\core.registers[20][16] ),
    .A3(\core.registers[21][16] ),
    .S0(net1484),
    .S1(net1586),
    .X(_06190_));
 sky130_fd_sc_hd__a22o_1 _11203_ (.A1(net1649),
    .A2(\core.registers[22][16] ),
    .B1(\core.registers[23][16] ),
    .B2(net1484),
    .X(_06191_));
 sky130_fd_sc_hd__a22o_1 _11204_ (.A1(net1649),
    .A2(\core.registers[18][16] ),
    .B1(\core.registers[19][16] ),
    .B2(net1484),
    .X(_06192_));
 sky130_fd_sc_hd__mux2_1 _11205_ (.A0(_06191_),
    .A1(_06192_),
    .S(net1574),
    .X(_06193_));
 sky130_fd_sc_hd__a21o_1 _11206_ (.A1(net1548),
    .A2(_06193_),
    .B1(net1570),
    .X(_06194_));
 sky130_fd_sc_hd__a21o_1 _11207_ (.A1(net1531),
    .A2(_06190_),
    .B1(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__a21o_1 _11208_ (.A1(_06189_),
    .A2(_06195_),
    .B1(net1594),
    .X(_06196_));
 sky130_fd_sc_hd__o211a_2 _11209_ (.A1(net1598),
    .A2(_06183_),
    .B1(_06196_),
    .C1(net1046),
    .X(_06197_));
 sky130_fd_sc_hd__a21o_4 _11210_ (.A1(net1096),
    .A2(_06132_),
    .B1(_06197_),
    .X(_06198_));
 sky130_fd_sc_hd__mux2_4 _11211_ (.A0(net1747),
    .A1(_06198_),
    .S(net1253),
    .X(_06199_));
 sky130_fd_sc_hd__inv_2 _11212_ (.A(_06199_),
    .Y(_06200_));
 sky130_fd_sc_hd__and2_2 _11213_ (.A(_06169_),
    .B(_06199_),
    .X(_06201_));
 sky130_fd_sc_hd__nor2_4 _11214_ (.A(_06169_),
    .B(_06199_),
    .Y(_06202_));
 sky130_fd_sc_hd__nor2_4 _11215_ (.A(_06201_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__a21o_1 _11216_ (.A1(\core.pipe1_csrData[15] ),
    .A2(net1247),
    .B1(net1238),
    .X(_06204_));
 sky130_fd_sc_hd__and3_1 _11217_ (.A(_03982_),
    .B(_03984_),
    .C(_03991_),
    .X(_06205_));
 sky130_fd_sc_hd__nor2_1 _11218_ (.A(_03986_),
    .B(_03993_),
    .Y(_06206_));
 sky130_fd_sc_hd__nor2_1 _11219_ (.A(_04015_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__a21o_1 _11220_ (.A1(_04007_),
    .A2(_05593_),
    .B1(_04018_),
    .X(_06208_));
 sky130_fd_sc_hd__o22a_1 _11221_ (.A1(_04038_),
    .A2(_06205_),
    .B1(_06207_),
    .B2(_06208_),
    .X(_06209_));
 sky130_fd_sc_hd__o21a_1 _11222_ (.A1(net1242),
    .A2(_06209_),
    .B1(_06204_),
    .X(_06210_));
 sky130_fd_sc_hd__o22a_4 _11223_ (.A1(\core.pipe1_resultRegister[15] ),
    .A2(net1189),
    .B1(_06210_),
    .B2(net1246),
    .X(_06211_));
 sky130_fd_sc_hd__or2_1 _11224_ (.A(\core.registers[5][15] ),
    .B(net1359),
    .X(_06212_));
 sky130_fd_sc_hd__o211a_1 _11225_ (.A1(\core.registers[4][15] ),
    .A2(net1384),
    .B1(_06212_),
    .C1(net1450),
    .X(_06213_));
 sky130_fd_sc_hd__mux2_1 _11226_ (.A0(\core.registers[0][15] ),
    .A1(\core.registers[1][15] ),
    .S(net1384),
    .X(_06214_));
 sky130_fd_sc_hd__a211o_1 _11227_ (.A1(net1438),
    .A2(_06214_),
    .B1(_06213_),
    .C1(net1345),
    .X(_06215_));
 sky130_fd_sc_hd__o221a_1 _11228_ (.A1(net1682),
    .A2(\core.registers[7][15] ),
    .B1(net1385),
    .B2(\core.registers[6][15] ),
    .C1(net1450),
    .X(_06216_));
 sky130_fd_sc_hd__o221a_1 _11229_ (.A1(net1682),
    .A2(\core.registers[3][15] ),
    .B1(net1384),
    .B2(\core.registers[2][15] ),
    .C1(net1438),
    .X(_06217_));
 sky130_fd_sc_hd__o31a_1 _11230_ (.A1(net1330),
    .A2(_06216_),
    .A3(_06217_),
    .B1(_04087_),
    .X(_06218_));
 sky130_fd_sc_hd__or2_1 _11231_ (.A(\core.registers[16][15] ),
    .B(net1382),
    .X(_06219_));
 sky130_fd_sc_hd__o211a_1 _11232_ (.A1(\core.registers[17][15] ),
    .A2(net1359),
    .B1(_06219_),
    .C1(net1438),
    .X(_06220_));
 sky130_fd_sc_hd__mux2_1 _11233_ (.A0(\core.registers[20][15] ),
    .A1(\core.registers[21][15] ),
    .S(net1382),
    .X(_06221_));
 sky130_fd_sc_hd__a211o_1 _11234_ (.A1(net1450),
    .A2(_06221_),
    .B1(_06220_),
    .C1(net1345),
    .X(_06222_));
 sky130_fd_sc_hd__o221a_1 _11235_ (.A1(net1682),
    .A2(\core.registers[23][15] ),
    .B1(net1382),
    .B2(\core.registers[22][15] ),
    .C1(net1450),
    .X(_06223_));
 sky130_fd_sc_hd__o221a_1 _11236_ (.A1(net1680),
    .A2(\core.registers[19][15] ),
    .B1(net1382),
    .B2(\core.registers[18][15] ),
    .C1(net1438),
    .X(_06224_));
 sky130_fd_sc_hd__o31a_1 _11237_ (.A1(net1330),
    .A2(_06223_),
    .A3(_06224_),
    .B1(net1325),
    .X(_06225_));
 sky130_fd_sc_hd__mux2_1 _11238_ (.A0(\core.registers[12][15] ),
    .A1(\core.registers[13][15] ),
    .S(net1382),
    .X(_06226_));
 sky130_fd_sc_hd__mux2_1 _11239_ (.A0(\core.registers[14][15] ),
    .A1(\core.registers[15][15] ),
    .S(net1382),
    .X(_06227_));
 sky130_fd_sc_hd__mux2_1 _11240_ (.A0(_06226_),
    .A1(_06227_),
    .S(net1345),
    .X(_06228_));
 sky130_fd_sc_hd__mux2_1 _11241_ (.A0(\core.registers[28][15] ),
    .A1(\core.registers[29][15] ),
    .S(net1382),
    .X(_06229_));
 sky130_fd_sc_hd__and3_1 _11242_ (.A(net1770),
    .B(\core.registers[31][15] ),
    .C(net1382),
    .X(_06230_));
 sky130_fd_sc_hd__a31o_1 _11243_ (.A1(net1770),
    .A2(net1682),
    .A3(\core.registers[30][15] ),
    .B1(net1709),
    .X(_06231_));
 sky130_fd_sc_hd__a211o_1 _11244_ (.A1(net1700),
    .A2(_06229_),
    .B1(_06230_),
    .C1(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__o211a_1 _11245_ (.A1(net1755),
    .A2(_06228_),
    .B1(_06232_),
    .C1(net1763),
    .X(_06233_));
 sky130_fd_sc_hd__mux2_1 _11246_ (.A0(\core.registers[8][15] ),
    .A1(\core.registers[9][15] ),
    .S(net1382),
    .X(_06234_));
 sky130_fd_sc_hd__mux2_1 _11247_ (.A0(\core.registers[10][15] ),
    .A1(\core.registers[11][15] ),
    .S(net1382),
    .X(_06235_));
 sky130_fd_sc_hd__mux2_1 _11248_ (.A0(_06234_),
    .A1(_06235_),
    .S(net1345),
    .X(_06236_));
 sky130_fd_sc_hd__mux2_1 _11249_ (.A0(\core.registers[24][15] ),
    .A1(\core.registers[25][15] ),
    .S(net1383),
    .X(_06237_));
 sky130_fd_sc_hd__a22o_1 _11250_ (.A1(net1682),
    .A2(\core.registers[26][15] ),
    .B1(\core.registers[27][15] ),
    .B2(net1383),
    .X(_06238_));
 sky130_fd_sc_hd__mux2_1 _11251_ (.A0(_06237_),
    .A1(_06238_),
    .S(net1770),
    .X(_06239_));
 sky130_fd_sc_hd__mux2_1 _11252_ (.A0(_06236_),
    .A1(_06239_),
    .S(net1755),
    .X(_06240_));
 sky130_fd_sc_hd__a21o_1 _11253_ (.A1(_06215_),
    .A2(_06218_),
    .B1(net1431),
    .X(_06241_));
 sky130_fd_sc_hd__a21o_1 _11254_ (.A1(_06222_),
    .A2(_06225_),
    .B1(_06241_),
    .X(_06242_));
 sky130_fd_sc_hd__a211o_1 _11255_ (.A1(net1705),
    .A2(_06240_),
    .B1(_06233_),
    .C1(net1428),
    .X(_06243_));
 sky130_fd_sc_hd__a21o_2 _11256_ (.A1(_06242_),
    .A2(_06243_),
    .B1(net1148),
    .X(_06244_));
 sky130_fd_sc_hd__o211ai_4 _11257_ (.A1(net1143),
    .A2(net743),
    .B1(_06244_),
    .C1(net1240),
    .Y(_06245_));
 sky130_fd_sc_hd__nor2_1 _11258_ (.A(net1040),
    .B(_06245_),
    .Y(_06246_));
 sky130_fd_sc_hd__o22a_2 _11259_ (.A1(net1793),
    .A2(net1257),
    .B1(net1006),
    .B2(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__inv_2 _11260_ (.A(_06247_),
    .Y(_06248_));
 sky130_fd_sc_hd__or2_2 _11261_ (.A(net456),
    .B(net1253),
    .X(_06249_));
 sky130_fd_sc_hd__mux4_1 _11262_ (.A0(\core.registers[16][15] ),
    .A1(\core.registers[17][15] ),
    .A2(\core.registers[20][15] ),
    .A3(\core.registers[21][15] ),
    .S0(net1481),
    .S1(net1585),
    .X(_06250_));
 sky130_fd_sc_hd__a22o_1 _11263_ (.A1(net1648),
    .A2(\core.registers[22][15] ),
    .B1(\core.registers[23][15] ),
    .B2(net1481),
    .X(_06251_));
 sky130_fd_sc_hd__a22o_1 _11264_ (.A1(net1647),
    .A2(\core.registers[18][15] ),
    .B1(\core.registers[19][15] ),
    .B2(net1481),
    .X(_06252_));
 sky130_fd_sc_hd__mux2_1 _11265_ (.A0(_06251_),
    .A1(_06252_),
    .S(net1574),
    .X(_06253_));
 sky130_fd_sc_hd__a21o_1 _11266_ (.A1(net1547),
    .A2(_06253_),
    .B1(net1567),
    .X(_06254_));
 sky130_fd_sc_hd__a21oi_1 _11267_ (.A1(net1530),
    .A2(_06250_),
    .B1(_06254_),
    .Y(_06255_));
 sky130_fd_sc_hd__a22o_1 _11268_ (.A1(net1648),
    .A2(\core.registers[30][15] ),
    .B1(\core.registers[31][15] ),
    .B2(net1481),
    .X(_06256_));
 sky130_fd_sc_hd__a22o_1 _11269_ (.A1(net1648),
    .A2(\core.registers[26][15] ),
    .B1(\core.registers[27][15] ),
    .B2(net1482),
    .X(_06257_));
 sky130_fd_sc_hd__mux2_1 _11270_ (.A0(_06256_),
    .A1(_06257_),
    .S(net1574),
    .X(_06258_));
 sky130_fd_sc_hd__mux4_1 _11271_ (.A0(\core.registers[24][15] ),
    .A1(\core.registers[25][15] ),
    .A2(\core.registers[28][15] ),
    .A3(\core.registers[29][15] ),
    .S0(net1481),
    .S1(net1585),
    .X(_06259_));
 sky130_fd_sc_hd__a21o_1 _11272_ (.A1(net1530),
    .A2(_06259_),
    .B1(net1562),
    .X(_06260_));
 sky130_fd_sc_hd__a21oi_2 _11273_ (.A1(net1547),
    .A2(_06258_),
    .B1(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__mux4_1 _11274_ (.A0(\core.registers[0][15] ),
    .A1(\core.registers[1][15] ),
    .A2(\core.registers[4][15] ),
    .A3(\core.registers[5][15] ),
    .S0(net1483),
    .S1(net1586),
    .X(_06262_));
 sky130_fd_sc_hd__and2_1 _11275_ (.A(net1530),
    .B(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__a22o_1 _11276_ (.A1(net1648),
    .A2(\core.registers[6][15] ),
    .B1(\core.registers[7][15] ),
    .B2(net1481),
    .X(_06264_));
 sky130_fd_sc_hd__a22o_1 _11277_ (.A1(net1648),
    .A2(\core.registers[2][15] ),
    .B1(\core.registers[3][15] ),
    .B2(net1483),
    .X(_06265_));
 sky130_fd_sc_hd__mux2_1 _11278_ (.A0(_06264_),
    .A1(_06265_),
    .S(net1574),
    .X(_06266_));
 sky130_fd_sc_hd__a21o_1 _11279_ (.A1(net1547),
    .A2(_06266_),
    .B1(net1567),
    .X(_06267_));
 sky130_fd_sc_hd__nor2_1 _11280_ (.A(_06263_),
    .B(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__mux4_1 _11281_ (.A0(\core.registers[8][15] ),
    .A1(\core.registers[9][15] ),
    .A2(\core.registers[12][15] ),
    .A3(\core.registers[13][15] ),
    .S0(net1481),
    .S1(net1585),
    .X(_06269_));
 sky130_fd_sc_hd__nand2_1 _11282_ (.A(net1530),
    .B(_06269_),
    .Y(_06270_));
 sky130_fd_sc_hd__a22o_1 _11283_ (.A1(net1647),
    .A2(\core.registers[14][15] ),
    .B1(\core.registers[15][15] ),
    .B2(net1481),
    .X(_06271_));
 sky130_fd_sc_hd__a22o_1 _11284_ (.A1(net1647),
    .A2(\core.registers[10][15] ),
    .B1(\core.registers[11][15] ),
    .B2(net1481),
    .X(_06272_));
 sky130_fd_sc_hd__mux2_1 _11285_ (.A0(_06271_),
    .A1(_06272_),
    .S(net1574),
    .X(_06273_));
 sky130_fd_sc_hd__a21oi_1 _11286_ (.A1(net1547),
    .A2(_06273_),
    .B1(net1562),
    .Y(_06274_));
 sky130_fd_sc_hd__a21o_1 _11287_ (.A1(_06270_),
    .A2(_06274_),
    .B1(net1598),
    .X(_06275_));
 sky130_fd_sc_hd__o32a_4 _11288_ (.A1(net1593),
    .A2(_06255_),
    .A3(_06261_),
    .B1(_06268_),
    .B2(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__a2bb2o_4 _11289_ (.A1_N(net1045),
    .A2_N(_06276_),
    .B1(net743),
    .B2(net1097),
    .X(_06277_));
 sky130_fd_sc_hd__o21ai_4 _11290_ (.A1(net1263),
    .A2(_06277_),
    .B1(_06249_),
    .Y(_06278_));
 sky130_fd_sc_hd__nor2_4 _11291_ (.A(_06248_),
    .B(_06278_),
    .Y(_06279_));
 sky130_fd_sc_hd__and2_2 _11292_ (.A(_06248_),
    .B(_06278_),
    .X(_06280_));
 sky130_fd_sc_hd__nor2_4 _11293_ (.A(_06279_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__inv_4 _11294_ (.A(_06281_),
    .Y(_06282_));
 sky130_fd_sc_hd__a21o_1 _11295_ (.A1(\core.pipe1_csrData[14] ),
    .A2(net1249),
    .B1(net1237),
    .X(_06283_));
 sky130_fd_sc_hd__o22ai_1 _11296_ (.A1(_04015_),
    .A2(_05072_),
    .B1(_05666_),
    .B2(_04008_),
    .Y(_06284_));
 sky130_fd_sc_hd__o22a_1 _11297_ (.A1(_04038_),
    .A2(_04470_),
    .B1(_06284_),
    .B2(_04018_),
    .X(_06285_));
 sky130_fd_sc_hd__o21a_1 _11298_ (.A1(net1242),
    .A2(_06285_),
    .B1(_06283_),
    .X(_06286_));
 sky130_fd_sc_hd__o22a_4 _11299_ (.A1(\core.pipe1_resultRegister[14] ),
    .A2(_03934_),
    .B1(_06286_),
    .B2(net1245),
    .X(_06287_));
 sky130_fd_sc_hd__or2_1 _11300_ (.A(\core.registers[5][14] ),
    .B(net1357),
    .X(_06288_));
 sky130_fd_sc_hd__o211a_1 _11301_ (.A1(\core.registers[4][14] ),
    .A2(net1369),
    .B1(_06288_),
    .C1(net1447),
    .X(_06289_));
 sky130_fd_sc_hd__mux2_1 _11302_ (.A0(\core.registers[0][14] ),
    .A1(\core.registers[1][14] ),
    .S(net1369),
    .X(_06290_));
 sky130_fd_sc_hd__a211o_1 _11303_ (.A1(net1434),
    .A2(_06290_),
    .B1(_06289_),
    .C1(net1342),
    .X(_06291_));
 sky130_fd_sc_hd__o221a_1 _11304_ (.A1(net1678),
    .A2(\core.registers[7][14] ),
    .B1(net1367),
    .B2(\core.registers[6][14] ),
    .C1(net1447),
    .X(_06292_));
 sky130_fd_sc_hd__o221a_1 _11305_ (.A1(net1678),
    .A2(\core.registers[3][14] ),
    .B1(net1369),
    .B2(\core.registers[2][14] ),
    .C1(net1434),
    .X(_06293_));
 sky130_fd_sc_hd__o31a_1 _11306_ (.A1(net1328),
    .A2(_06292_),
    .A3(_06293_),
    .B1(net1320),
    .X(_06294_));
 sky130_fd_sc_hd__or2_1 _11307_ (.A(\core.registers[16][14] ),
    .B(net1367),
    .X(_06295_));
 sky130_fd_sc_hd__o211a_1 _11308_ (.A1(\core.registers[17][14] ),
    .A2(net1357),
    .B1(_06295_),
    .C1(net1434),
    .X(_06296_));
 sky130_fd_sc_hd__mux2_1 _11309_ (.A0(\core.registers[20][14] ),
    .A1(\core.registers[21][14] ),
    .S(net1367),
    .X(_06297_));
 sky130_fd_sc_hd__a211o_1 _11310_ (.A1(net1447),
    .A2(_06297_),
    .B1(_06296_),
    .C1(net1342),
    .X(_06298_));
 sky130_fd_sc_hd__o221a_1 _11311_ (.A1(net1675),
    .A2(\core.registers[23][14] ),
    .B1(net1366),
    .B2(\core.registers[22][14] ),
    .C1(net1447),
    .X(_06299_));
 sky130_fd_sc_hd__o221a_1 _11312_ (.A1(net1676),
    .A2(\core.registers[19][14] ),
    .B1(net1366),
    .B2(\core.registers[18][14] ),
    .C1(net1434),
    .X(_06300_));
 sky130_fd_sc_hd__o31a_1 _11313_ (.A1(net1328),
    .A2(_06299_),
    .A3(_06300_),
    .B1(net1324),
    .X(_06301_));
 sky130_fd_sc_hd__mux2_1 _11314_ (.A0(\core.registers[12][14] ),
    .A1(\core.registers[13][14] ),
    .S(net1365),
    .X(_06302_));
 sky130_fd_sc_hd__mux2_1 _11315_ (.A0(\core.registers[14][14] ),
    .A1(\core.registers[15][14] ),
    .S(net1365),
    .X(_06303_));
 sky130_fd_sc_hd__mux2_1 _11316_ (.A0(_06302_),
    .A1(_06303_),
    .S(net1341),
    .X(_06304_));
 sky130_fd_sc_hd__mux2_1 _11317_ (.A0(\core.registers[28][14] ),
    .A1(\core.registers[29][14] ),
    .S(net1365),
    .X(_06305_));
 sky130_fd_sc_hd__and3_1 _11318_ (.A(net1768),
    .B(\core.registers[31][14] ),
    .C(net1365),
    .X(_06306_));
 sky130_fd_sc_hd__a31o_1 _11319_ (.A1(net1768),
    .A2(net1675),
    .A3(\core.registers[30][14] ),
    .B1(net1708),
    .X(_06307_));
 sky130_fd_sc_hd__a211o_1 _11320_ (.A1(net1699),
    .A2(_06305_),
    .B1(_06306_),
    .C1(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__o211a_1 _11321_ (.A1(net1753),
    .A2(_06304_),
    .B1(_06308_),
    .C1(net1763),
    .X(_06309_));
 sky130_fd_sc_hd__mux2_1 _11322_ (.A0(\core.registers[8][14] ),
    .A1(\core.registers[9][14] ),
    .S(net1365),
    .X(_06310_));
 sky130_fd_sc_hd__mux2_1 _11323_ (.A0(\core.registers[10][14] ),
    .A1(\core.registers[11][14] ),
    .S(net1365),
    .X(_06311_));
 sky130_fd_sc_hd__mux2_1 _11324_ (.A0(_06310_),
    .A1(_06311_),
    .S(net1341),
    .X(_06312_));
 sky130_fd_sc_hd__mux2_1 _11325_ (.A0(\core.registers[24][14] ),
    .A1(\core.registers[25][14] ),
    .S(net1365),
    .X(_06313_));
 sky130_fd_sc_hd__a22o_1 _11326_ (.A1(net1675),
    .A2(\core.registers[26][14] ),
    .B1(\core.registers[27][14] ),
    .B2(net1365),
    .X(_06314_));
 sky130_fd_sc_hd__mux2_1 _11327_ (.A0(_06313_),
    .A1(_06314_),
    .S(net1768),
    .X(_06315_));
 sky130_fd_sc_hd__mux2_1 _11328_ (.A0(_06312_),
    .A1(_06315_),
    .S(net1753),
    .X(_06316_));
 sky130_fd_sc_hd__a21o_1 _11329_ (.A1(_06291_),
    .A2(_06294_),
    .B1(net1429),
    .X(_06317_));
 sky130_fd_sc_hd__a21o_1 _11330_ (.A1(_06298_),
    .A2(_06301_),
    .B1(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__a211o_2 _11331_ (.A1(net1704),
    .A2(_06316_),
    .B1(_06309_),
    .C1(net1427),
    .X(_06319_));
 sky130_fd_sc_hd__a21o_4 _11332_ (.A1(_06318_),
    .A2(_06319_),
    .B1(net1148),
    .X(_06320_));
 sky130_fd_sc_hd__o211ai_4 _11333_ (.A1(net1142),
    .A2(_06287_),
    .B1(_06320_),
    .C1(net1239),
    .Y(_06321_));
 sky130_fd_sc_hd__nor2_1 _11334_ (.A(net1040),
    .B(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__o22a_1 _11335_ (.A1(net1794),
    .A2(net1253),
    .B1(net1006),
    .B2(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__inv_2 _11336_ (.A(_06323_),
    .Y(_06324_));
 sky130_fd_sc_hd__or2_2 _11337_ (.A(net455),
    .B(net1253),
    .X(_06325_));
 sky130_fd_sc_hd__mux4_1 _11338_ (.A0(\core.registers[16][14] ),
    .A1(\core.registers[17][14] ),
    .A2(\core.registers[20][14] ),
    .A3(\core.registers[21][14] ),
    .S0(net1466),
    .S1(net1583),
    .X(_06326_));
 sky130_fd_sc_hd__a22o_1 _11339_ (.A1(net1641),
    .A2(\core.registers[22][14] ),
    .B1(\core.registers[23][14] ),
    .B2(net1465),
    .X(_06327_));
 sky130_fd_sc_hd__a22o_1 _11340_ (.A1(net1641),
    .A2(\core.registers[18][14] ),
    .B1(\core.registers[19][14] ),
    .B2(net1465),
    .X(_06328_));
 sky130_fd_sc_hd__mux2_1 _11341_ (.A0(_06327_),
    .A1(_06328_),
    .S(net1571),
    .X(_06329_));
 sky130_fd_sc_hd__a21o_1 _11342_ (.A1(net1542),
    .A2(_06329_),
    .B1(net1566),
    .X(_06330_));
 sky130_fd_sc_hd__a21oi_1 _11343_ (.A1(net1526),
    .A2(_06326_),
    .B1(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__a22o_1 _11344_ (.A1(net1641),
    .A2(\core.registers[30][14] ),
    .B1(\core.registers[31][14] ),
    .B2(net1464),
    .X(_06332_));
 sky130_fd_sc_hd__a22o_1 _11345_ (.A1(net1641),
    .A2(\core.registers[26][14] ),
    .B1(\core.registers[27][14] ),
    .B2(net1464),
    .X(_06333_));
 sky130_fd_sc_hd__mux2_1 _11346_ (.A0(_06332_),
    .A1(_06333_),
    .S(net1571),
    .X(_06334_));
 sky130_fd_sc_hd__mux4_1 _11347_ (.A0(\core.registers[24][14] ),
    .A1(\core.registers[25][14] ),
    .A2(\core.registers[28][14] ),
    .A3(\core.registers[29][14] ),
    .S0(net1464),
    .S1(net1582),
    .X(_06335_));
 sky130_fd_sc_hd__a21o_1 _11348_ (.A1(net1526),
    .A2(_06335_),
    .B1(net1561),
    .X(_06336_));
 sky130_fd_sc_hd__a21oi_2 _11349_ (.A1(net1543),
    .A2(_06334_),
    .B1(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__mux4_2 _11350_ (.A0(\core.registers[0][14] ),
    .A1(\core.registers[1][14] ),
    .A2(\core.registers[4][14] ),
    .A3(\core.registers[5][14] ),
    .S0(net1467),
    .S1(net1582),
    .X(_06338_));
 sky130_fd_sc_hd__and2_1 _11351_ (.A(net1526),
    .B(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__a22o_1 _11352_ (.A1(net1643),
    .A2(\core.registers[6][14] ),
    .B1(\core.registers[7][14] ),
    .B2(net1466),
    .X(_06340_));
 sky130_fd_sc_hd__a22o_1 _11353_ (.A1(net1644),
    .A2(\core.registers[2][14] ),
    .B1(\core.registers[3][14] ),
    .B2(net1466),
    .X(_06341_));
 sky130_fd_sc_hd__mux2_1 _11354_ (.A0(_06340_),
    .A1(_06341_),
    .S(net1571),
    .X(_06342_));
 sky130_fd_sc_hd__a21o_1 _11355_ (.A1(net1542),
    .A2(_06342_),
    .B1(net1566),
    .X(_06343_));
 sky130_fd_sc_hd__nor2_1 _11356_ (.A(_06339_),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__mux4_2 _11357_ (.A0(\core.registers[8][14] ),
    .A1(\core.registers[9][14] ),
    .A2(\core.registers[12][14] ),
    .A3(\core.registers[13][14] ),
    .S0(net1464),
    .S1(net1582),
    .X(_06345_));
 sky130_fd_sc_hd__nand2_1 _11358_ (.A(net1526),
    .B(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__a22o_1 _11359_ (.A1(net1641),
    .A2(\core.registers[14][14] ),
    .B1(\core.registers[15][14] ),
    .B2(net1464),
    .X(_06347_));
 sky130_fd_sc_hd__a22o_1 _11360_ (.A1(net1641),
    .A2(\core.registers[10][14] ),
    .B1(\core.registers[11][14] ),
    .B2(net1464),
    .X(_06348_));
 sky130_fd_sc_hd__mux2_1 _11361_ (.A0(_06347_),
    .A1(_06348_),
    .S(net1571),
    .X(_06349_));
 sky130_fd_sc_hd__a21oi_1 _11362_ (.A1(net1543),
    .A2(_06349_),
    .B1(net1561),
    .Y(_06350_));
 sky130_fd_sc_hd__a21o_1 _11363_ (.A1(_06346_),
    .A2(_06350_),
    .B1(net1597),
    .X(_06351_));
 sky130_fd_sc_hd__o32a_4 _11364_ (.A1(net1593),
    .A2(_06331_),
    .A3(_06337_),
    .B1(_06344_),
    .B2(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__a2bb2o_4 _11365_ (.A1_N(net1045),
    .A2_N(_06352_),
    .B1(_06287_),
    .B2(net1094),
    .X(_06353_));
 sky130_fd_sc_hd__o21ai_4 _11366_ (.A1(net1263),
    .A2(_06353_),
    .B1(_06325_),
    .Y(_06354_));
 sky130_fd_sc_hd__nor2_2 _11367_ (.A(_06324_),
    .B(_06354_),
    .Y(_06355_));
 sky130_fd_sc_hd__and2_2 _11368_ (.A(_06324_),
    .B(_06354_),
    .X(_06356_));
 sky130_fd_sc_hd__nor2_4 _11369_ (.A(_06355_),
    .B(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__inv_2 _11370_ (.A(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__a21o_1 _11371_ (.A1(\core.pipe1_csrData[13] ),
    .A2(net1250),
    .B1(net1237),
    .X(_06359_));
 sky130_fd_sc_hd__o22ai_1 _11372_ (.A1(_04015_),
    .A2(_05150_),
    .B1(_05744_),
    .B2(_04008_),
    .Y(_06360_));
 sky130_fd_sc_hd__o22a_1 _11373_ (.A1(_04038_),
    .A2(_04556_),
    .B1(_06360_),
    .B2(_04018_),
    .X(_06361_));
 sky130_fd_sc_hd__o21a_1 _11374_ (.A1(net1242),
    .A2(_06361_),
    .B1(_06359_),
    .X(_06362_));
 sky130_fd_sc_hd__o22a_2 _11375_ (.A1(\core.pipe1_resultRegister[13] ),
    .A2(net1188),
    .B1(_06362_),
    .B2(net1245),
    .X(_06363_));
 sky130_fd_sc_hd__nor2_1 _11376_ (.A(net1144),
    .B(net735),
    .Y(_06364_));
 sky130_fd_sc_hd__or2_1 _11377_ (.A(\core.registers[5][13] ),
    .B(net1360),
    .X(_06365_));
 sky130_fd_sc_hd__o211a_1 _11378_ (.A1(\core.registers[4][13] ),
    .A2(net1423),
    .B1(_06365_),
    .C1(net1455),
    .X(_06366_));
 sky130_fd_sc_hd__mux2_1 _11379_ (.A0(\core.registers[0][13] ),
    .A1(\core.registers[1][13] ),
    .S(net1425),
    .X(_06367_));
 sky130_fd_sc_hd__a211o_1 _11380_ (.A1(net1444),
    .A2(_06367_),
    .B1(_06366_),
    .C1(net1353),
    .X(_06368_));
 sky130_fd_sc_hd__o221a_1 _11381_ (.A1(net1696),
    .A2(\core.registers[7][13] ),
    .B1(net1422),
    .B2(\core.registers[6][13] ),
    .C1(net1455),
    .X(_06369_));
 sky130_fd_sc_hd__o221a_1 _11382_ (.A1(net1696),
    .A2(\core.registers[3][13] ),
    .B1(net1422),
    .B2(\core.registers[2][13] ),
    .C1(net1444),
    .X(_06370_));
 sky130_fd_sc_hd__o31a_1 _11383_ (.A1(net1339),
    .A2(_06369_),
    .A3(_06370_),
    .B1(net1322),
    .X(_06371_));
 sky130_fd_sc_hd__or2_1 _11384_ (.A(\core.registers[16][13] ),
    .B(net1422),
    .X(_06372_));
 sky130_fd_sc_hd__o211a_1 _11385_ (.A1(\core.registers[17][13] ),
    .A2(net1361),
    .B1(_06372_),
    .C1(net1444),
    .X(_06373_));
 sky130_fd_sc_hd__mux2_1 _11386_ (.A0(\core.registers[20][13] ),
    .A1(\core.registers[21][13] ),
    .S(net1420),
    .X(_06374_));
 sky130_fd_sc_hd__a211o_1 _11387_ (.A1(net1455),
    .A2(_06374_),
    .B1(_06373_),
    .C1(net1352),
    .X(_06375_));
 sky130_fd_sc_hd__o221a_1 _11388_ (.A1(net1693),
    .A2(\core.registers[23][13] ),
    .B1(net1422),
    .B2(\core.registers[22][13] ),
    .C1(net1455),
    .X(_06376_));
 sky130_fd_sc_hd__o221a_1 _11389_ (.A1(net1693),
    .A2(\core.registers[19][13] ),
    .B1(net1420),
    .B2(\core.registers[18][13] ),
    .C1(net1444),
    .X(_06377_));
 sky130_fd_sc_hd__o31a_1 _11390_ (.A1(net1337),
    .A2(_06376_),
    .A3(_06377_),
    .B1(net1326),
    .X(_06378_));
 sky130_fd_sc_hd__mux2_1 _11391_ (.A0(\core.registers[12][13] ),
    .A1(\core.registers[13][13] ),
    .S(net1421),
    .X(_06379_));
 sky130_fd_sc_hd__mux2_1 _11392_ (.A0(\core.registers[14][13] ),
    .A1(\core.registers[15][13] ),
    .S(net1421),
    .X(_06380_));
 sky130_fd_sc_hd__mux2_1 _11393_ (.A0(_06379_),
    .A1(_06380_),
    .S(net1352),
    .X(_06381_));
 sky130_fd_sc_hd__mux2_1 _11394_ (.A0(\core.registers[28][13] ),
    .A1(\core.registers[29][13] ),
    .S(net1416),
    .X(_06382_));
 sky130_fd_sc_hd__and3_1 _11395_ (.A(net1774),
    .B(\core.registers[31][13] ),
    .C(net1416),
    .X(_06383_));
 sky130_fd_sc_hd__a31o_1 _11396_ (.A1(net1774),
    .A2(net1695),
    .A3(\core.registers[30][13] ),
    .B1(net1710),
    .X(_06384_));
 sky130_fd_sc_hd__a211o_1 _11397_ (.A1(net1701),
    .A2(_06382_),
    .B1(_06383_),
    .C1(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__o211a_1 _11398_ (.A1(net1760),
    .A2(_06381_),
    .B1(_06385_),
    .C1(net1766),
    .X(_06386_));
 sky130_fd_sc_hd__or2_1 _11399_ (.A(\core.registers[9][13] ),
    .B(net1360),
    .X(_06387_));
 sky130_fd_sc_hd__o211a_1 _11400_ (.A1(\core.registers[8][13] ),
    .A2(net1416),
    .B1(net1338),
    .C1(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__a22o_1 _11401_ (.A1(net1692),
    .A2(\core.registers[10][13] ),
    .B1(\core.registers[11][13] ),
    .B2(net1421),
    .X(_06389_));
 sky130_fd_sc_hd__a21o_1 _11402_ (.A1(net1352),
    .A2(_06389_),
    .B1(net1760),
    .X(_06390_));
 sky130_fd_sc_hd__mux2_1 _11403_ (.A0(\core.registers[24][13] ),
    .A1(\core.registers[25][13] ),
    .S(net1426),
    .X(_06391_));
 sky130_fd_sc_hd__a22o_1 _11404_ (.A1(net1695),
    .A2(\core.registers[26][13] ),
    .B1(\core.registers[27][13] ),
    .B2(net1417),
    .X(_06392_));
 sky130_fd_sc_hd__mux2_1 _11405_ (.A0(_06391_),
    .A1(_06392_),
    .S(net1774),
    .X(_06393_));
 sky130_fd_sc_hd__o221a_2 _11406_ (.A1(_06388_),
    .A2(_06390_),
    .B1(_06393_),
    .B2(net1710),
    .C1(net1707),
    .X(_06394_));
 sky130_fd_sc_hd__a21o_1 _11407_ (.A1(_06368_),
    .A2(_06371_),
    .B1(net1433),
    .X(_06395_));
 sky130_fd_sc_hd__a21o_2 _11408_ (.A1(_06375_),
    .A2(_06378_),
    .B1(_06395_),
    .X(_06396_));
 sky130_fd_sc_hd__o31ai_4 _11409_ (.A1(_04077_),
    .A2(_06386_),
    .A3(_06394_),
    .B1(_06396_),
    .Y(_06397_));
 sky130_fd_sc_hd__a211o_4 _11410_ (.A1(net1145),
    .A2(_06397_),
    .B1(_06364_),
    .C1(_04095_),
    .X(_06398_));
 sky130_fd_sc_hd__nor2_1 _11411_ (.A(net1041),
    .B(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__o22a_2 _11412_ (.A1(\core.pipe0_currentInstruction[13] ),
    .A2(net1257),
    .B1(net1006),
    .B2(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__mux4_1 _11413_ (.A0(\core.registers[16][13] ),
    .A1(\core.registers[17][13] ),
    .A2(\core.registers[20][13] ),
    .A3(\core.registers[21][13] ),
    .S0(net1519),
    .S1(net1590),
    .X(_06401_));
 sky130_fd_sc_hd__a22o_1 _11414_ (.A1(net1658),
    .A2(\core.registers[22][13] ),
    .B1(\core.registers[23][13] ),
    .B2(net1519),
    .X(_06402_));
 sky130_fd_sc_hd__a22o_1 _11415_ (.A1(net1658),
    .A2(\core.registers[18][13] ),
    .B1(\core.registers[19][13] ),
    .B2(net1519),
    .X(_06403_));
 sky130_fd_sc_hd__mux2_1 _11416_ (.A0(_06402_),
    .A1(_06403_),
    .S(net1578),
    .X(_06404_));
 sky130_fd_sc_hd__a21o_1 _11417_ (.A1(net1557),
    .A2(_06404_),
    .B1(net1568),
    .X(_06405_));
 sky130_fd_sc_hd__a21oi_2 _11418_ (.A1(net1538),
    .A2(_06401_),
    .B1(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__mux4_1 _11419_ (.A0(\core.registers[24][13] ),
    .A1(\core.registers[25][13] ),
    .A2(\core.registers[28][13] ),
    .A3(\core.registers[29][13] ),
    .S0(net1516),
    .S1(net1591),
    .X(_06407_));
 sky130_fd_sc_hd__a22o_1 _11420_ (.A1(net1661),
    .A2(\core.registers[30][13] ),
    .B1(\core.registers[31][13] ),
    .B2(net1516),
    .X(_06408_));
 sky130_fd_sc_hd__a22o_1 _11421_ (.A1(net1661),
    .A2(\core.registers[26][13] ),
    .B1(\core.registers[27][13] ),
    .B2(net1515),
    .X(_06409_));
 sky130_fd_sc_hd__mux2_1 _11422_ (.A0(_06408_),
    .A1(_06409_),
    .S(net1579),
    .X(_06410_));
 sky130_fd_sc_hd__a21o_1 _11423_ (.A1(net1559),
    .A2(_06410_),
    .B1(net1564),
    .X(_06411_));
 sky130_fd_sc_hd__a21oi_2 _11424_ (.A1(net1540),
    .A2(_06407_),
    .B1(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__a22o_1 _11425_ (.A1(net1660),
    .A2(\core.registers[6][13] ),
    .B1(\core.registers[7][13] ),
    .B2(net1523),
    .X(_06413_));
 sky130_fd_sc_hd__a22o_1 _11426_ (.A1(net1660),
    .A2(\core.registers[2][13] ),
    .B1(\core.registers[3][13] ),
    .B2(net1519),
    .X(_06414_));
 sky130_fd_sc_hd__mux2_1 _11427_ (.A0(_06413_),
    .A1(_06414_),
    .S(net1578),
    .X(_06415_));
 sky130_fd_sc_hd__and2_1 _11428_ (.A(net1557),
    .B(_06415_),
    .X(_06416_));
 sky130_fd_sc_hd__mux4_1 _11429_ (.A0(\core.registers[0][13] ),
    .A1(\core.registers[1][13] ),
    .A2(\core.registers[4][13] ),
    .A3(\core.registers[5][13] ),
    .S0(net1522),
    .S1(net1591),
    .X(_06417_));
 sky130_fd_sc_hd__a21o_1 _11430_ (.A1(net1538),
    .A2(_06417_),
    .B1(net1569),
    .X(_06418_));
 sky130_fd_sc_hd__nor2_1 _11431_ (.A(_06416_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__mux4_1 _11432_ (.A0(\core.registers[8][13] ),
    .A1(\core.registers[9][13] ),
    .A2(\core.registers[12][13] ),
    .A3(\core.registers[13][13] ),
    .S0(net1520),
    .S1(net1590),
    .X(_06420_));
 sky130_fd_sc_hd__nand2_1 _11433_ (.A(net1538),
    .B(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__a22o_1 _11434_ (.A1(net1658),
    .A2(\core.registers[14][13] ),
    .B1(\core.registers[15][13] ),
    .B2(net1520),
    .X(_06422_));
 sky130_fd_sc_hd__a22o_1 _11435_ (.A1(net1658),
    .A2(\core.registers[10][13] ),
    .B1(\core.registers[11][13] ),
    .B2(net1520),
    .X(_06423_));
 sky130_fd_sc_hd__mux2_1 _11436_ (.A0(_06422_),
    .A1(_06423_),
    .S(net1578),
    .X(_06424_));
 sky130_fd_sc_hd__a21oi_1 _11437_ (.A1(net1557),
    .A2(_06424_),
    .B1(net1565),
    .Y(_06425_));
 sky130_fd_sc_hd__a21o_1 _11438_ (.A1(_06421_),
    .A2(_06425_),
    .B1(net1599),
    .X(_06426_));
 sky130_fd_sc_hd__o32a_4 _11439_ (.A1(net1595),
    .A2(_06406_),
    .A3(_06412_),
    .B1(_06419_),
    .B2(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__a2bb2o_4 _11440_ (.A1_N(_03946_),
    .A2_N(_06427_),
    .B1(net735),
    .B2(net1095),
    .X(_06428_));
 sky130_fd_sc_hd__or2_2 _11441_ (.A(net454),
    .B(net1258),
    .X(_06429_));
 sky130_fd_sc_hd__o21ai_4 _11442_ (.A1(net1263),
    .A2(_06428_),
    .B1(_06429_),
    .Y(_06430_));
 sky130_fd_sc_hd__clkinv_2 _11443_ (.A(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__and2_4 _11444_ (.A(_06400_),
    .B(_06431_),
    .X(_06432_));
 sky130_fd_sc_hd__nor2_4 _11445_ (.A(_06400_),
    .B(_06431_),
    .Y(_06433_));
 sky130_fd_sc_hd__nor2_8 _11446_ (.A(_06432_),
    .B(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__a21o_1 _11447_ (.A1(\core.pipe1_csrData[12] ),
    .A2(net1250),
    .B1(_04887_),
    .X(_06435_));
 sky130_fd_sc_hd__o22ai_1 _11448_ (.A1(_04015_),
    .A2(_05222_),
    .B1(_05821_),
    .B2(_04008_),
    .Y(_06436_));
 sky130_fd_sc_hd__o22a_1 _11449_ (.A1(_04038_),
    .A2(_04642_),
    .B1(_06436_),
    .B2(_04018_),
    .X(_06437_));
 sky130_fd_sc_hd__o21a_1 _11450_ (.A1(net1242),
    .A2(_06437_),
    .B1(_06435_),
    .X(_06438_));
 sky130_fd_sc_hd__o22a_2 _11451_ (.A1(\core.pipe1_resultRegister[12] ),
    .A2(net1188),
    .B1(_06438_),
    .B2(net1245),
    .X(_06439_));
 sky130_fd_sc_hd__nor2_1 _11452_ (.A(net1144),
    .B(net731),
    .Y(_06440_));
 sky130_fd_sc_hd__or2_1 _11453_ (.A(\core.registers[5][12] ),
    .B(net1360),
    .X(_06441_));
 sky130_fd_sc_hd__o211a_1 _11454_ (.A1(\core.registers[4][12] ),
    .A2(net1424),
    .B1(_06441_),
    .C1(net1455),
    .X(_06442_));
 sky130_fd_sc_hd__mux2_1 _11455_ (.A0(\core.registers[0][12] ),
    .A1(\core.registers[1][12] ),
    .S(net1424),
    .X(_06443_));
 sky130_fd_sc_hd__a211o_1 _11456_ (.A1(net1444),
    .A2(_06443_),
    .B1(_06442_),
    .C1(net1353),
    .X(_06444_));
 sky130_fd_sc_hd__o221a_1 _11457_ (.A1(net1696),
    .A2(\core.registers[7][12] ),
    .B1(net1423),
    .B2(\core.registers[6][12] ),
    .C1(net1455),
    .X(_06445_));
 sky130_fd_sc_hd__o221a_1 _11458_ (.A1(net1697),
    .A2(\core.registers[3][12] ),
    .B1(net1423),
    .B2(\core.registers[2][12] ),
    .C1(net1444),
    .X(_06446_));
 sky130_fd_sc_hd__o31a_1 _11459_ (.A1(net1339),
    .A2(_06445_),
    .A3(_06446_),
    .B1(net1322),
    .X(_06447_));
 sky130_fd_sc_hd__or2_1 _11460_ (.A(\core.registers[16][12] ),
    .B(net1423),
    .X(_06448_));
 sky130_fd_sc_hd__o211a_1 _11461_ (.A1(\core.registers[17][12] ),
    .A2(net1360),
    .B1(_06448_),
    .C1(net1444),
    .X(_06449_));
 sky130_fd_sc_hd__mux2_1 _11462_ (.A0(\core.registers[20][12] ),
    .A1(\core.registers[21][12] ),
    .S(net1423),
    .X(_06450_));
 sky130_fd_sc_hd__a211o_1 _11463_ (.A1(net1455),
    .A2(_06450_),
    .B1(_06449_),
    .C1(net1353),
    .X(_06451_));
 sky130_fd_sc_hd__o221a_1 _11464_ (.A1(net1696),
    .A2(\core.registers[23][12] ),
    .B1(net1423),
    .B2(\core.registers[22][12] ),
    .C1(net1455),
    .X(_06452_));
 sky130_fd_sc_hd__o221a_1 _11465_ (.A1(net1696),
    .A2(\core.registers[19][12] ),
    .B1(net1423),
    .B2(\core.registers[18][12] ),
    .C1(net1445),
    .X(_06453_));
 sky130_fd_sc_hd__o31a_1 _11466_ (.A1(net1337),
    .A2(_06452_),
    .A3(_06453_),
    .B1(net1326),
    .X(_06454_));
 sky130_fd_sc_hd__o21a_1 _11467_ (.A1(\core.registers[12][12] ),
    .A2(net1421),
    .B1(net1337),
    .X(_06455_));
 sky130_fd_sc_hd__o21ai_1 _11468_ (.A1(\core.registers[13][12] ),
    .A2(net1361),
    .B1(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__a22o_1 _11469_ (.A1(net1692),
    .A2(\core.registers[14][12] ),
    .B1(\core.registers[15][12] ),
    .B2(net1421),
    .X(_06457_));
 sky130_fd_sc_hd__nand2_1 _11470_ (.A(net1352),
    .B(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__mux2_1 _11471_ (.A0(\core.registers[28][12] ),
    .A1(\core.registers[29][12] ),
    .S(net1417),
    .X(_06459_));
 sky130_fd_sc_hd__and3_1 _11472_ (.A(net1774),
    .B(\core.registers[31][12] ),
    .C(net1405),
    .X(_06460_));
 sky130_fd_sc_hd__a211o_1 _11473_ (.A1(\core.registers[30][12] ),
    .A2(net1319),
    .B1(_06460_),
    .C1(net1711),
    .X(_06461_));
 sky130_fd_sc_hd__a21oi_2 _11474_ (.A1(net1703),
    .A2(_06459_),
    .B1(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__a311o_1 _11475_ (.A1(net1711),
    .A2(_06456_),
    .A3(_06458_),
    .B1(_06462_),
    .C1(_03835_),
    .X(_06463_));
 sky130_fd_sc_hd__mux2_1 _11476_ (.A0(\core.registers[8][12] ),
    .A1(\core.registers[9][12] ),
    .S(net1421),
    .X(_06464_));
 sky130_fd_sc_hd__mux2_1 _11477_ (.A0(\core.registers[10][12] ),
    .A1(\core.registers[11][12] ),
    .S(net1421),
    .X(_06465_));
 sky130_fd_sc_hd__mux2_2 _11478_ (.A0(_06464_),
    .A1(_06465_),
    .S(net1352),
    .X(_06466_));
 sky130_fd_sc_hd__or2_1 _11479_ (.A(\core.registers[25][12] ),
    .B(net1360),
    .X(_06467_));
 sky130_fd_sc_hd__o211a_2 _11480_ (.A1(\core.registers[24][12] ),
    .A2(net1417),
    .B1(_06467_),
    .C1(net1702),
    .X(_06468_));
 sky130_fd_sc_hd__and3_1 _11481_ (.A(net1774),
    .B(\core.registers[27][12] ),
    .C(net1417),
    .X(_06469_));
 sky130_fd_sc_hd__a211o_2 _11482_ (.A1(\core.registers[26][12] ),
    .A2(net1319),
    .B1(_06469_),
    .C1(net1711),
    .X(_06470_));
 sky130_fd_sc_hd__o221ai_4 _11483_ (.A1(net1760),
    .A2(_06466_),
    .B1(_06468_),
    .B2(_06470_),
    .C1(_03835_),
    .Y(_06471_));
 sky130_fd_sc_hd__a21o_1 _11484_ (.A1(_06444_),
    .A2(_06447_),
    .B1(net1433),
    .X(_06472_));
 sky130_fd_sc_hd__a21oi_2 _11485_ (.A1(_06451_),
    .A2(_06454_),
    .B1(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__a31o_2 _11486_ (.A1(_04076_),
    .A2(_06463_),
    .A3(_06471_),
    .B1(_06473_),
    .X(_06474_));
 sky130_fd_sc_hd__a211o_4 _11487_ (.A1(net1145),
    .A2(_06474_),
    .B1(_06440_),
    .C1(_04095_),
    .X(_06475_));
 sky130_fd_sc_hd__nor2_1 _11488_ (.A(net1040),
    .B(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__o22a_2 _11489_ (.A1(\core.pipe0_currentInstruction[12] ),
    .A2(net1257),
    .B1(net1006),
    .B2(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__or2_2 _11490_ (.A(net453),
    .B(net1257),
    .X(_06478_));
 sky130_fd_sc_hd__mux4_2 _11491_ (.A0(\core.registers[16][12] ),
    .A1(\core.registers[17][12] ),
    .A2(\core.registers[20][12] ),
    .A3(\core.registers[21][12] ),
    .S0(net1521),
    .S1(net1590),
    .X(_06479_));
 sky130_fd_sc_hd__a22o_1 _11492_ (.A1(net1659),
    .A2(\core.registers[22][12] ),
    .B1(\core.registers[23][12] ),
    .B2(net1521),
    .X(_06480_));
 sky130_fd_sc_hd__a22o_1 _11493_ (.A1(net1659),
    .A2(\core.registers[18][12] ),
    .B1(\core.registers[19][12] ),
    .B2(net1521),
    .X(_06481_));
 sky130_fd_sc_hd__mux2_1 _11494_ (.A0(_06480_),
    .A1(_06481_),
    .S(net1578),
    .X(_06482_));
 sky130_fd_sc_hd__a21o_1 _11495_ (.A1(net1557),
    .A2(_06482_),
    .B1(net1569),
    .X(_06483_));
 sky130_fd_sc_hd__a21oi_2 _11496_ (.A1(net1539),
    .A2(_06479_),
    .B1(_06483_),
    .Y(_06484_));
 sky130_fd_sc_hd__a22o_1 _11497_ (.A1(net1654),
    .A2(\core.registers[30][12] ),
    .B1(\core.registers[31][12] ),
    .B2(net1504),
    .X(_06485_));
 sky130_fd_sc_hd__a22o_1 _11498_ (.A1(net1661),
    .A2(\core.registers[26][12] ),
    .B1(\core.registers[27][12] ),
    .B2(net1515),
    .X(_06486_));
 sky130_fd_sc_hd__mux2_2 _11499_ (.A0(_06485_),
    .A1(_06486_),
    .S(net1579),
    .X(_06487_));
 sky130_fd_sc_hd__mux4_1 _11500_ (.A0(\core.registers[24][12] ),
    .A1(\core.registers[25][12] ),
    .A2(\core.registers[28][12] ),
    .A3(\core.registers[29][12] ),
    .S0(net1515),
    .S1(net1591),
    .X(_06488_));
 sky130_fd_sc_hd__a21o_1 _11501_ (.A1(net1540),
    .A2(_06488_),
    .B1(net1564),
    .X(_06489_));
 sky130_fd_sc_hd__a21oi_4 _11502_ (.A1(net1559),
    .A2(_06487_),
    .B1(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__mux4_1 _11503_ (.A0(\core.registers[0][12] ),
    .A1(\core.registers[1][12] ),
    .A2(\core.registers[4][12] ),
    .A3(\core.registers[5][12] ),
    .S0(net1522),
    .S1(net1591),
    .X(_06491_));
 sky130_fd_sc_hd__and2_1 _11504_ (.A(net1538),
    .B(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__a22o_1 _11505_ (.A1(net1660),
    .A2(\core.registers[6][12] ),
    .B1(\core.registers[7][12] ),
    .B2(net1521),
    .X(_06493_));
 sky130_fd_sc_hd__a22o_1 _11506_ (.A1(net1660),
    .A2(\core.registers[2][12] ),
    .B1(\core.registers[3][12] ),
    .B2(net1521),
    .X(_06494_));
 sky130_fd_sc_hd__mux2_1 _11507_ (.A0(_06493_),
    .A1(_06494_),
    .S(net1579),
    .X(_06495_));
 sky130_fd_sc_hd__a21o_1 _11508_ (.A1(net1557),
    .A2(_06495_),
    .B1(net1570),
    .X(_06496_));
 sky130_fd_sc_hd__nor2_1 _11509_ (.A(_06492_),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__mux4_1 _11510_ (.A0(\core.registers[8][12] ),
    .A1(\core.registers[9][12] ),
    .A2(\core.registers[12][12] ),
    .A3(\core.registers[13][12] ),
    .S0(net1520),
    .S1(net1590),
    .X(_06498_));
 sky130_fd_sc_hd__nand2_1 _11511_ (.A(net1538),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__a22o_1 _11512_ (.A1(net1658),
    .A2(\core.registers[14][12] ),
    .B1(\core.registers[15][12] ),
    .B2(net1520),
    .X(_06500_));
 sky130_fd_sc_hd__a22o_1 _11513_ (.A1(net1659),
    .A2(\core.registers[10][12] ),
    .B1(\core.registers[11][12] ),
    .B2(net1520),
    .X(_06501_));
 sky130_fd_sc_hd__mux2_1 _11514_ (.A0(_06500_),
    .A1(_06501_),
    .S(net1578),
    .X(_06502_));
 sky130_fd_sc_hd__a21oi_1 _11515_ (.A1(net1557),
    .A2(_06502_),
    .B1(net1565),
    .Y(_06503_));
 sky130_fd_sc_hd__a21o_1 _11516_ (.A1(_06499_),
    .A2(_06503_),
    .B1(net1600),
    .X(_06504_));
 sky130_fd_sc_hd__o32a_4 _11517_ (.A1(net1595),
    .A2(_06484_),
    .A3(_06490_),
    .B1(_06497_),
    .B2(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__a2bb2o_4 _11518_ (.A1_N(net1044),
    .A2_N(_06505_),
    .B1(net731),
    .B2(net1095),
    .X(_06506_));
 sky130_fd_sc_hd__o21ai_4 _11519_ (.A1(net1263),
    .A2(_06506_),
    .B1(_06478_),
    .Y(_06507_));
 sky130_fd_sc_hd__clkinv_2 _11520_ (.A(_06507_),
    .Y(_06508_));
 sky130_fd_sc_hd__and2_2 _11521_ (.A(_06477_),
    .B(_06508_),
    .X(_06509_));
 sky130_fd_sc_hd__nor2_2 _11522_ (.A(_06477_),
    .B(_06508_),
    .Y(_06510_));
 sky130_fd_sc_hd__nor2_4 _11523_ (.A(_06509_),
    .B(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__clkinv_4 _11524_ (.A(_06511_),
    .Y(_06512_));
 sky130_fd_sc_hd__o21ba_4 _11525_ (.A1(_04131_),
    .A2(_05067_),
    .B1_N(_04132_),
    .X(_06513_));
 sky130_fd_sc_hd__o21bai_4 _11526_ (.A1(_06512_),
    .A2(_06513_),
    .B1_N(_06509_),
    .Y(_06514_));
 sky130_fd_sc_hd__a21oi_4 _11527_ (.A1(_06434_),
    .A2(_06514_),
    .B1(_06432_),
    .Y(_06515_));
 sky130_fd_sc_hd__o21bai_4 _11528_ (.A1(_06358_),
    .A2(_06515_),
    .B1_N(_06355_),
    .Y(_06516_));
 sky130_fd_sc_hd__a21oi_4 _11529_ (.A1(_06281_),
    .A2(_06516_),
    .B1(_06279_),
    .Y(_06517_));
 sky130_fd_sc_hd__o21bai_4 _11530_ (.A1(_06202_),
    .A2(_06517_),
    .B1_N(_06201_),
    .Y(_06518_));
 sky130_fd_sc_hd__a21oi_4 _11531_ (.A1(_06127_),
    .A2(_06518_),
    .B1(_06125_),
    .Y(_06519_));
 sky130_fd_sc_hd__o21ai_4 _11532_ (.A1(_06051_),
    .A2(_06519_),
    .B1(_06048_),
    .Y(_06520_));
 sky130_fd_sc_hd__o211ai_4 _11533_ (.A1(_06051_),
    .A2(_06519_),
    .B1(_05972_),
    .C1(_06048_),
    .Y(_06521_));
 sky130_fd_sc_hd__nand2_2 _11534_ (.A(_05973_),
    .B(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__a31o_2 _11535_ (.A1(_05897_),
    .A2(_05973_),
    .A3(_06521_),
    .B1(_05895_),
    .X(_06523_));
 sky130_fd_sc_hd__o21a_1 _11536_ (.A1(_05820_),
    .A2(_05895_),
    .B1(_05818_),
    .X(_06524_));
 sky130_fd_sc_hd__nor2_8 _11537_ (.A(_05819_),
    .B(_05820_),
    .Y(_06525_));
 sky130_fd_sc_hd__a41o_4 _11538_ (.A1(_05897_),
    .A2(_05973_),
    .A3(_06521_),
    .A4(_06525_),
    .B1(_06524_),
    .X(_06526_));
 sky130_fd_sc_hd__a21o_2 _11539_ (.A1(_05742_),
    .A2(_06526_),
    .B1(_05740_),
    .X(_06527_));
 sky130_fd_sc_hd__o21ba_1 _11540_ (.A1(_05664_),
    .A2(_05740_),
    .B1_N(_05665_),
    .X(_06528_));
 sky130_fd_sc_hd__nor2_8 _11541_ (.A(_05664_),
    .B(_05665_),
    .Y(_06529_));
 sky130_fd_sc_hd__a31o_4 _11542_ (.A1(_05742_),
    .A2(_06526_),
    .A3(_06529_),
    .B1(_06528_),
    .X(_06530_));
 sky130_fd_sc_hd__a21o_2 _11543_ (.A1(_05591_),
    .A2(_06530_),
    .B1(_05589_),
    .X(_06531_));
 sky130_fd_sc_hd__o21ba_1 _11544_ (.A1(_05515_),
    .A2(_05589_),
    .B1_N(_05514_),
    .X(_06532_));
 sky130_fd_sc_hd__nor2_4 _11545_ (.A(_05514_),
    .B(_05515_),
    .Y(_06533_));
 sky130_fd_sc_hd__inv_2 _11546_ (.A(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__a31o_4 _11547_ (.A1(_05591_),
    .A2(_06530_),
    .A3(_06533_),
    .B1(_06532_),
    .X(_06535_));
 sky130_fd_sc_hd__a21oi_4 _11548_ (.A1(_05443_),
    .A2(_06535_),
    .B1(_05440_),
    .Y(_06536_));
 sky130_fd_sc_hd__o21a_1 _11549_ (.A1(_05369_),
    .A2(_05440_),
    .B1(_05368_),
    .X(_06537_));
 sky130_fd_sc_hd__nor2_8 _11550_ (.A(_05367_),
    .B(_05369_),
    .Y(_06538_));
 sky130_fd_sc_hd__a31o_4 _11551_ (.A1(_05443_),
    .A2(_06535_),
    .A3(_06538_),
    .B1(_06537_),
    .X(_06539_));
 sky130_fd_sc_hd__a311o_2 _11552_ (.A1(_05443_),
    .A2(_06535_),
    .A3(_06538_),
    .B1(_06537_),
    .C1(_05295_),
    .X(_06540_));
 sky130_fd_sc_hd__nand2_2 _11553_ (.A(_05294_),
    .B(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__a31o_4 _11554_ (.A1(_05220_),
    .A2(_05294_),
    .A3(_06540_),
    .B1(_05221_),
    .X(_06542_));
 sky130_fd_sc_hd__xnor2_4 _11555_ (.A(_05149_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__or3_1 _11556_ (.A(_03894_),
    .B(_03981_),
    .C(net1616),
    .X(_06544_));
 sky130_fd_sc_hd__a211oi_2 _11557_ (.A1(_04013_),
    .A2(_06544_),
    .B1(_06206_),
    .C1(net1242),
    .Y(_06545_));
 sky130_fd_sc_hd__a221o_4 _11558_ (.A1(\core.pipe1_csrData[31] ),
    .A2(net1248),
    .B1(_03935_),
    .B2(\core.pipe1_resultRegister[31] ),
    .C1(_06545_),
    .X(_06546_));
 sky130_fd_sc_hd__mux4_1 _11559_ (.A0(\core.registers[16][31] ),
    .A1(\core.registers[17][31] ),
    .A2(\core.registers[20][31] ),
    .A3(\core.registers[21][31] ),
    .S0(net1379),
    .S1(net1448),
    .X(_06547_));
 sky130_fd_sc_hd__o22a_1 _11560_ (.A1(net1681),
    .A2(\core.registers[23][31] ),
    .B1(net1379),
    .B2(\core.registers[22][31] ),
    .X(_06548_));
 sky130_fd_sc_hd__o22a_1 _11561_ (.A1(net1681),
    .A2(\core.registers[19][31] ),
    .B1(net1380),
    .B2(\core.registers[18][31] ),
    .X(_06549_));
 sky130_fd_sc_hd__mux2_1 _11562_ (.A0(_06548_),
    .A1(_06549_),
    .S(net1435),
    .X(_06550_));
 sky130_fd_sc_hd__o21a_1 _11563_ (.A1(net1330),
    .A2(_06550_),
    .B1(net1324),
    .X(_06551_));
 sky130_fd_sc_hd__o21a_1 _11564_ (.A1(net1344),
    .A2(_06547_),
    .B1(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__o22a_1 _11565_ (.A1(net1680),
    .A2(\core.registers[7][31] ),
    .B1(net1380),
    .B2(\core.registers[6][31] ),
    .X(_06553_));
 sky130_fd_sc_hd__o22a_1 _11566_ (.A1(net1681),
    .A2(\core.registers[3][31] ),
    .B1(net1384),
    .B2(\core.registers[2][31] ),
    .X(_06554_));
 sky130_fd_sc_hd__mux2_1 _11567_ (.A0(_06553_),
    .A1(_06554_),
    .S(net1438),
    .X(_06555_));
 sky130_fd_sc_hd__or2_1 _11568_ (.A(net1330),
    .B(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__mux4_1 _11569_ (.A0(\core.registers[0][31] ),
    .A1(\core.registers[1][31] ),
    .A2(\core.registers[4][31] ),
    .A3(\core.registers[5][31] ),
    .S0(net1384),
    .S1(net1450),
    .X(_06557_));
 sky130_fd_sc_hd__o21a_1 _11570_ (.A1(net1344),
    .A2(_06557_),
    .B1(net1320),
    .X(_06558_));
 sky130_fd_sc_hd__a21oi_2 _11571_ (.A1(_06556_),
    .A2(_06558_),
    .B1(_06552_),
    .Y(_06559_));
 sky130_fd_sc_hd__a221o_1 _11572_ (.A1(net1675),
    .A2(\core.registers[26][31] ),
    .B1(\core.registers[27][31] ),
    .B2(net1371),
    .C1(net1699),
    .X(_06560_));
 sky130_fd_sc_hd__mux2_1 _11573_ (.A0(\core.registers[24][31] ),
    .A1(\core.registers[25][31] ),
    .S(net1363),
    .X(_06561_));
 sky130_fd_sc_hd__o21a_1 _11574_ (.A1(net1768),
    .A2(_06561_),
    .B1(_06560_),
    .X(_06562_));
 sky130_fd_sc_hd__mux2_1 _11575_ (.A0(\core.registers[8][31] ),
    .A1(\core.registers[9][31] ),
    .S(net1363),
    .X(_06563_));
 sky130_fd_sc_hd__mux2_1 _11576_ (.A0(\core.registers[10][31] ),
    .A1(\core.registers[11][31] ),
    .S(net1363),
    .X(_06564_));
 sky130_fd_sc_hd__mux2_1 _11577_ (.A0(_06563_),
    .A1(_06564_),
    .S(net1341),
    .X(_06565_));
 sky130_fd_sc_hd__mux2_1 _11578_ (.A0(_06562_),
    .A1(_06565_),
    .S(net1708),
    .X(_06566_));
 sky130_fd_sc_hd__nor2_1 _11579_ (.A(net1763),
    .B(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__a221o_1 _11580_ (.A1(net1679),
    .A2(\core.registers[30][31] ),
    .B1(\core.registers[31][31] ),
    .B2(net1379),
    .C1(net1700),
    .X(_06568_));
 sky130_fd_sc_hd__mux2_1 _11581_ (.A0(\core.registers[28][31] ),
    .A1(\core.registers[29][31] ),
    .S(net1379),
    .X(_06569_));
 sky130_fd_sc_hd__o21ai_1 _11582_ (.A1(net1771),
    .A2(_06569_),
    .B1(_06568_),
    .Y(_06570_));
 sky130_fd_sc_hd__nand2_1 _11583_ (.A(net1754),
    .B(_06570_),
    .Y(_06571_));
 sky130_fd_sc_hd__a221o_1 _11584_ (.A1(net1679),
    .A2(\core.registers[14][31] ),
    .B1(\core.registers[15][31] ),
    .B2(net1369),
    .C1(net1699),
    .X(_06572_));
 sky130_fd_sc_hd__a31o_1 _11585_ (.A1(net1776),
    .A2(\core.registers[13][31] ),
    .A3(net1629),
    .B1(net1768),
    .X(_06573_));
 sky130_fd_sc_hd__a21o_1 _11586_ (.A1(\core.registers[12][31] ),
    .A2(net1358),
    .B1(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__a21o_1 _11587_ (.A1(_06572_),
    .A2(_06574_),
    .B1(net1754),
    .X(_06575_));
 sky130_fd_sc_hd__a21oi_1 _11588_ (.A1(_06571_),
    .A2(_06575_),
    .B1(net1704),
    .Y(_06576_));
 sky130_fd_sc_hd__o31a_1 _11589_ (.A1(net1427),
    .A2(_06567_),
    .A3(_06576_),
    .B1(net1143),
    .X(_06577_));
 sky130_fd_sc_hd__o21ai_2 _11590_ (.A1(net1429),
    .A2(_06559_),
    .B1(_06577_),
    .Y(_06578_));
 sky130_fd_sc_hd__o211a_2 _11591_ (.A1(net1141),
    .A2(net1025),
    .B1(_06578_),
    .C1(net1239),
    .X(_06579_));
 sky130_fd_sc_hd__mux2_4 _11592_ (.A0(net1751),
    .A1(_06579_),
    .S(_04129_),
    .X(_06580_));
 sky130_fd_sc_hd__mux2_1 _11593_ (.A0(\core.registers[28][31] ),
    .A1(\core.registers[29][31] ),
    .S(net1478),
    .X(_06581_));
 sky130_fd_sc_hd__a221o_1 _11594_ (.A1(net1644),
    .A2(\core.registers[30][31] ),
    .B1(\core.registers[31][31] ),
    .B2(net1478),
    .C1(net1663),
    .X(_06582_));
 sky130_fd_sc_hd__mux2_1 _11595_ (.A0(\core.registers[24][31] ),
    .A1(\core.registers[25][31] ),
    .S(net1462),
    .X(_06583_));
 sky130_fd_sc_hd__a221o_1 _11596_ (.A1(net1642),
    .A2(\core.registers[26][31] ),
    .B1(\core.registers[27][31] ),
    .B2(net1463),
    .C1(net1663),
    .X(_06584_));
 sky130_fd_sc_hd__mux2_1 _11597_ (.A0(\core.registers[8][31] ),
    .A1(\core.registers[9][31] ),
    .S(net1462),
    .X(_06585_));
 sky130_fd_sc_hd__mux2_1 _11598_ (.A0(\core.registers[10][31] ),
    .A1(\core.registers[11][31] ),
    .S(net1462),
    .X(_06586_));
 sky130_fd_sc_hd__mux2_1 _11599_ (.A0(_06585_),
    .A1(_06586_),
    .S(net1543),
    .X(_06587_));
 sky130_fd_sc_hd__o21ai_1 _11600_ (.A1(net1787),
    .A2(_06583_),
    .B1(_06584_),
    .Y(_06588_));
 sky130_fd_sc_hd__nand2_1 _11601_ (.A(net1778),
    .B(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__o211a_2 _11602_ (.A1(net1778),
    .A2(_06587_),
    .B1(_06589_),
    .C1(net1668),
    .X(_06590_));
 sky130_fd_sc_hd__o21a_1 _11603_ (.A1(net1788),
    .A2(_06581_),
    .B1(_06582_),
    .X(_06591_));
 sky130_fd_sc_hd__mux2_1 _11604_ (.A0(\core.registers[12][31] ),
    .A1(\core.registers[13][31] ),
    .S(net1467),
    .X(_06592_));
 sky130_fd_sc_hd__mux2_1 _11605_ (.A0(\core.registers[14][31] ),
    .A1(\core.registers[15][31] ),
    .S(net1468),
    .X(_06593_));
 sky130_fd_sc_hd__mux2_1 _11606_ (.A0(_06592_),
    .A1(_06593_),
    .S(net1543),
    .X(_06594_));
 sky130_fd_sc_hd__mux2_1 _11607_ (.A0(_06591_),
    .A1(_06594_),
    .S(net1674),
    .X(_06595_));
 sky130_fd_sc_hd__a211o_1 _11608_ (.A1(net1784),
    .A2(_06595_),
    .B1(_06590_),
    .C1(net1561),
    .X(_06596_));
 sky130_fd_sc_hd__mux2_1 _11609_ (.A0(\core.registers[18][31] ),
    .A1(\core.registers[19][31] ),
    .S(net1479),
    .X(_06597_));
 sky130_fd_sc_hd__mux2_1 _11610_ (.A0(\core.registers[16][31] ),
    .A1(\core.registers[17][31] ),
    .S(net1478),
    .X(_06598_));
 sky130_fd_sc_hd__mux2_1 _11611_ (.A0(_06597_),
    .A1(_06598_),
    .S(net1528),
    .X(_06599_));
 sky130_fd_sc_hd__o221a_1 _11612_ (.A1(net1649),
    .A2(\core.registers[23][31] ),
    .B1(net1479),
    .B2(\core.registers[22][31] ),
    .C1(net1548),
    .X(_06600_));
 sky130_fd_sc_hd__mux2_1 _11613_ (.A0(\core.registers[20][31] ),
    .A1(\core.registers[21][31] ),
    .S(net1478),
    .X(_06601_));
 sky130_fd_sc_hd__mux2_1 _11614_ (.A0(\core.registers[0][31] ),
    .A1(\core.registers[1][31] ),
    .S(net1483),
    .X(_06602_));
 sky130_fd_sc_hd__mux2_1 _11615_ (.A0(\core.registers[2][31] ),
    .A1(\core.registers[3][31] ),
    .S(net1483),
    .X(_06603_));
 sky130_fd_sc_hd__mux2_1 _11616_ (.A0(_06602_),
    .A1(_06603_),
    .S(net1548),
    .X(_06604_));
 sky130_fd_sc_hd__mux2_1 _11617_ (.A0(\core.registers[4][31] ),
    .A1(\core.registers[5][31] ),
    .S(net1483),
    .X(_06605_));
 sky130_fd_sc_hd__o221a_1 _11618_ (.A1(net1649),
    .A2(\core.registers[7][31] ),
    .B1(net1478),
    .B2(\core.registers[6][31] ),
    .C1(net1548),
    .X(_06606_));
 sky130_fd_sc_hd__a211o_1 _11619_ (.A1(net1530),
    .A2(_06605_),
    .B1(_06606_),
    .C1(net1574),
    .X(_06607_));
 sky130_fd_sc_hd__a211o_1 _11620_ (.A1(net1528),
    .A2(_06601_),
    .B1(_06600_),
    .C1(net1572),
    .X(_06608_));
 sky130_fd_sc_hd__o211a_1 _11621_ (.A1(net1585),
    .A2(_06599_),
    .B1(_06608_),
    .C1(net1597),
    .X(_06609_));
 sky130_fd_sc_hd__o211a_1 _11622_ (.A1(net1585),
    .A2(_06604_),
    .B1(_06607_),
    .C1(net1594),
    .X(_06610_));
 sky130_fd_sc_hd__o31a_2 _11623_ (.A1(net1566),
    .A2(_06609_),
    .A3(_06610_),
    .B1(_06596_),
    .X(_06611_));
 sky130_fd_sc_hd__a22oi_4 _11624_ (.A1(net1097),
    .A2(net1025),
    .B1(_06611_),
    .B2(net1046),
    .Y(_06612_));
 sky130_fd_sc_hd__mux2_8 _11625_ (.A0(_03823_),
    .A1(_06612_),
    .S(net1254),
    .X(_06613_));
 sky130_fd_sc_hd__inv_2 _11626_ (.A(_06613_),
    .Y(_06614_));
 sky130_fd_sc_hd__nor2_4 _11627_ (.A(_06580_),
    .B(_06613_),
    .Y(_06615_));
 sky130_fd_sc_hd__nand2_2 _11628_ (.A(_06580_),
    .B(_06613_),
    .Y(_06616_));
 sky130_fd_sc_hd__and2b_4 _11629_ (.A_N(_06615_),
    .B(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__a21oi_4 _11630_ (.A1(_05149_),
    .A2(_06542_),
    .B1(_05146_),
    .Y(_06618_));
 sky130_fd_sc_hd__xnor2_4 _11631_ (.A(_06617_),
    .B(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__and2_1 _11632_ (.A(_06543_),
    .B(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__nor2_1 _11633_ (.A(_05219_),
    .B(_05221_),
    .Y(_06621_));
 sky130_fd_sc_hd__or2_4 _11634_ (.A(_05219_),
    .B(_05221_),
    .X(_06622_));
 sky130_fd_sc_hd__xnor2_4 _11635_ (.A(_06541_),
    .B(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__nand2_8 _11636_ (.A(_05294_),
    .B(_05296_),
    .Y(_06624_));
 sky130_fd_sc_hd__xor2_4 _11637_ (.A(_06539_),
    .B(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__xor2_4 _11638_ (.A(_06536_),
    .B(_06538_),
    .X(_06626_));
 sky130_fd_sc_hd__xnor2_4 _11639_ (.A(_05442_),
    .B(_06535_),
    .Y(_06627_));
 sky130_fd_sc_hd__xnor2_4 _11640_ (.A(_06531_),
    .B(_06533_),
    .Y(_06628_));
 sky130_fd_sc_hd__clkinv_2 _11641_ (.A(_06628_),
    .Y(_06629_));
 sky130_fd_sc_hd__xnor2_4 _11642_ (.A(_05591_),
    .B(_06530_),
    .Y(_06630_));
 sky130_fd_sc_hd__clkinv_2 _11643_ (.A(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__and4b_1 _11644_ (.A_N(_06627_),
    .B(_06628_),
    .C(_06630_),
    .D(_06626_),
    .X(_06632_));
 sky130_fd_sc_hd__and4_4 _11645_ (.A(_06620_),
    .B(_06623_),
    .C(_06625_),
    .D(_06632_),
    .X(_06633_));
 sky130_fd_sc_hd__nor2_4 _11646_ (.A(_04053_),
    .B(net1043),
    .Y(_06634_));
 sky130_fd_sc_hd__or2_2 _11647_ (.A(_04053_),
    .B(net1043),
    .X(_06635_));
 sky130_fd_sc_hd__and2b_1 _11648_ (.A_N(_05050_),
    .B(net885),
    .X(_06636_));
 sky130_fd_sc_hd__nor2_1 _11649_ (.A(_05051_),
    .B(_06636_),
    .Y(_06637_));
 sky130_fd_sc_hd__or2_4 _11650_ (.A(_05051_),
    .B(_06636_),
    .X(_06638_));
 sky130_fd_sc_hd__nor2_1 _11651_ (.A(_04971_),
    .B(_05051_),
    .Y(_06639_));
 sky130_fd_sc_hd__nor2_1 _11652_ (.A(_05053_),
    .B(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__or2_4 _11653_ (.A(_05053_),
    .B(_06639_),
    .X(_06641_));
 sky130_fd_sc_hd__nor2_1 _11654_ (.A(net671),
    .B(net635),
    .Y(_06642_));
 sky130_fd_sc_hd__nand2_8 _11655_ (.A(net667),
    .B(net633),
    .Y(_06643_));
 sky130_fd_sc_hd__and2_4 _11656_ (.A(_04047_),
    .B(_04048_),
    .X(_06644_));
 sky130_fd_sc_hd__nand2_8 _11657_ (.A(_04047_),
    .B(_04048_),
    .Y(_06645_));
 sky130_fd_sc_hd__nand2_8 _11658_ (.A(_04071_),
    .B(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__mux2_1 _11659_ (.A0(_04060_),
    .A1(_06646_),
    .S(_04971_),
    .X(_06647_));
 sky130_fd_sc_hd__o22a_4 _11660_ (.A1(net991),
    .A2(net611),
    .B1(_06647_),
    .B2(_06638_),
    .X(_06648_));
 sky130_fd_sc_hd__and2_4 _11661_ (.A(_04071_),
    .B(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__nand2_4 _11662_ (.A(_04071_),
    .B(_06648_),
    .Y(_06650_));
 sky130_fd_sc_hd__nor2_1 _11663_ (.A(net1601),
    .B(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__and2_4 _11664_ (.A(_06633_),
    .B(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__a22o_4 _11665_ (.A1(\core.fetchProgramCounter[11] ),
    .A2(net1601),
    .B1(_05068_),
    .B2(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__nor2_2 _11666_ (.A(_06633_),
    .B(_06650_),
    .Y(_06654_));
 sky130_fd_sc_hd__xnor2_4 _11667_ (.A(_06527_),
    .B(_06529_),
    .Y(_06655_));
 sky130_fd_sc_hd__clkinv_4 _11668_ (.A(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__xnor2_4 _11669_ (.A(_05742_),
    .B(_06526_),
    .Y(_06657_));
 sky130_fd_sc_hd__clkinv_2 _11670_ (.A(_06657_),
    .Y(_06658_));
 sky130_fd_sc_hd__xor2_4 _11671_ (.A(_06523_),
    .B(_06525_),
    .X(_06659_));
 sky130_fd_sc_hd__xnor2_4 _11672_ (.A(_05897_),
    .B(_06522_),
    .Y(_06660_));
 sky130_fd_sc_hd__and2_4 _11673_ (.A(_05972_),
    .B(_05973_),
    .X(_06661_));
 sky130_fd_sc_hd__xor2_4 _11674_ (.A(_06520_),
    .B(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__xnor2_4 _11675_ (.A(_06050_),
    .B(_06519_),
    .Y(_06663_));
 sky130_fd_sc_hd__xnor2_4 _11676_ (.A(_06128_),
    .B(_06518_),
    .Y(_06664_));
 sky130_fd_sc_hd__xnor2_4 _11677_ (.A(_06203_),
    .B(_06517_),
    .Y(_06665_));
 sky130_fd_sc_hd__xnor2_4 _11678_ (.A(_06282_),
    .B(_06516_),
    .Y(_06666_));
 sky130_fd_sc_hd__xnor2_4 _11679_ (.A(_06357_),
    .B(_06515_),
    .Y(_06667_));
 sky130_fd_sc_hd__xor2_4 _11680_ (.A(_06434_),
    .B(_06514_),
    .X(_06668_));
 sky130_fd_sc_hd__xnor2_4 _11681_ (.A(_06512_),
    .B(_06513_),
    .Y(_06669_));
 sky130_fd_sc_hd__inv_2 _11682_ (.A(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__or3b_1 _11683_ (.A(_06668_),
    .B(_06670_),
    .C_N(_06651_),
    .X(_06671_));
 sky130_fd_sc_hd__or4_1 _11684_ (.A(_06665_),
    .B(_06666_),
    .C(_06667_),
    .D(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__or4_1 _11685_ (.A(_06662_),
    .B(_06663_),
    .C(_06664_),
    .D(_06672_),
    .X(_06673_));
 sky130_fd_sc_hd__or4_1 _11686_ (.A(_06658_),
    .B(_06659_),
    .C(_06660_),
    .D(_06673_),
    .X(_06674_));
 sky130_fd_sc_hd__nor2_2 _11687_ (.A(_04029_),
    .B(_06649_),
    .Y(_06675_));
 sky130_fd_sc_hd__nand2b_4 _11688_ (.A_N(\coreWBInterface.state[0] ),
    .B(\coreWBInterface.state[1] ),
    .Y(_06676_));
 sky130_fd_sc_hd__nand2_8 _11689_ (.A(_03854_),
    .B(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__nor2_1 _11690_ (.A(\memoryController.last_instruction_enableWB ),
    .B(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__a21o_1 _11691_ (.A1(\localMemoryInterface.coreReadReady ),
    .A2(net1635),
    .B1(net1638),
    .X(_06679_));
 sky130_fd_sc_hd__o21a_2 _11692_ (.A1(net1625),
    .A2(_06678_),
    .B1(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__nand2_1 _11693_ (.A(\memoryController.last_instruction_enableWB ),
    .B(net1635),
    .Y(_06681_));
 sky130_fd_sc_hd__nand2b_2 _11694_ (.A_N(net1315),
    .B(_06677_),
    .Y(_06682_));
 sky130_fd_sc_hd__or2_2 _11695_ (.A(\localMemoryInterface.coreReadReady ),
    .B(net1635),
    .X(_06683_));
 sky130_fd_sc_hd__o2111a_1 _11696_ (.A1(_06675_),
    .A2(_06680_),
    .B1(_06682_),
    .C1(_06683_),
    .D1(net1719),
    .X(_06684_));
 sky130_fd_sc_hd__o2111ai_4 _11697_ (.A1(_06675_),
    .A2(_06680_),
    .B1(_06682_),
    .C1(_06683_),
    .D1(net1719),
    .Y(_06685_));
 sky130_fd_sc_hd__or4_2 _11698_ (.A(\core.fetchProgramCounter[15] ),
    .B(\core.fetchProgramCounter[14] ),
    .C(\core.fetchProgramCounter[13] ),
    .D(\core.fetchProgramCounter[12] ),
    .X(_06686_));
 sky130_fd_sc_hd__or4_1 _11699_ (.A(\core.fetchProgramCounter[19] ),
    .B(\core.fetchProgramCounter[18] ),
    .C(\core.fetchProgramCounter[17] ),
    .D(\core.fetchProgramCounter[16] ),
    .X(_06687_));
 sky130_fd_sc_hd__or4_1 _11700_ (.A(\core.fetchProgramCounter[23] ),
    .B(\core.fetchProgramCounter[22] ),
    .C(\core.fetchProgramCounter[21] ),
    .D(\core.fetchProgramCounter[20] ),
    .X(_06688_));
 sky130_fd_sc_hd__or4_2 _11701_ (.A(_03876_),
    .B(_06686_),
    .C(_06687_),
    .D(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__o32a_4 _11702_ (.A1(_06654_),
    .A2(_06656_),
    .A3(_06674_),
    .B1(net598),
    .B2(_06689_),
    .X(_06690_));
 sky130_fd_sc_hd__a211oi_4 _11703_ (.A1(_04057_),
    .A2(net532),
    .B1(_06690_),
    .C1(\localMemoryInterface.coreReadReady ),
    .Y(_06691_));
 sky130_fd_sc_hd__nand2_1 _11704_ (.A(_06653_),
    .B(_06691_),
    .Y(net375));
 sky130_fd_sc_hd__nand2b_1 _11705_ (.A_N(_06653_),
    .B(_06691_),
    .Y(net374));
 sky130_fd_sc_hd__and3b_4 _11706_ (.A_N(_06690_),
    .B(net532),
    .C(_04057_),
    .X(_06692_));
 sky130_fd_sc_hd__or2_1 _11707_ (.A(\wbSRAMInterface.state[1] ),
    .B(\wbSRAMInterface.state[0] ),
    .X(_06693_));
 sky130_fd_sc_hd__or4_1 _11708_ (.A(\wbSRAMInterface.currentAddress[12] ),
    .B(\wbSRAMInterface.currentAddress[13] ),
    .C(\wbSRAMInterface.currentAddress[16] ),
    .D(\wbSRAMInterface.currentAddress[15] ),
    .X(_06694_));
 sky130_fd_sc_hd__o21a_1 _11709_ (.A1(\wbSRAMInterface.currentAddress[14] ),
    .A2(_06694_),
    .B1(net1615),
    .X(_06695_));
 sky130_fd_sc_hd__nand2_2 _11710_ (.A(\wbSRAMInterface.state[1] ),
    .B(\wbSRAMInterface.state[0] ),
    .Y(_06696_));
 sky130_fd_sc_hd__nand2_4 _11711_ (.A(net1615),
    .B(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__or2_1 _11712_ (.A(net1910),
    .B(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__o31a_4 _11713_ (.A1(\wbSRAMInterface.currentAddress[17] ),
    .A2(\wbSRAMInterface.currentAddress[18] ),
    .A3(\wbSRAMInterface.currentAddress[19] ),
    .B1(net1615),
    .X(_06699_));
 sky130_fd_sc_hd__or4_4 _11714_ (.A(\wbSRAMInterface.currentAddress[20] ),
    .B(\wbSRAMInterface.currentAddress[21] ),
    .C(\wbSRAMInterface.currentAddress[22] ),
    .D(\wbSRAMInterface.currentAddress[23] ),
    .X(_06700_));
 sky130_fd_sc_hd__nor4_4 _11715_ (.A(_06695_),
    .B(net1279),
    .C(_06699_),
    .D(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__and2b_4 _11716_ (.A_N(\wbSRAMInterface.state[1] ),
    .B(\wbSRAMInterface.state[0] ),
    .X(_06702_));
 sky130_fd_sc_hd__nand2b_4 _11717_ (.A_N(\wbSRAMInterface.state[1] ),
    .B(\wbSRAMInterface.state[0] ),
    .Y(_06703_));
 sky130_fd_sc_hd__a21oi_4 _11718_ (.A1(net1236),
    .A2(_06702_),
    .B1(net500),
    .Y(net483));
 sky130_fd_sc_hd__or3b_4 _11719_ (.A(net1738),
    .B(_06702_),
    .C_N(_06701_),
    .X(_06704_));
 sky130_fd_sc_hd__and2b_4 _11720_ (.A_N(net500),
    .B(net1236),
    .X(_06705_));
 sky130_fd_sc_hd__a22oi_4 _11721_ (.A1(_06653_),
    .A2(net500),
    .B1(_06705_),
    .B2(\wbSRAMInterface.currentAddress[11] ),
    .Y(_06706_));
 sky130_fd_sc_hd__a21o_1 _11722_ (.A1(net483),
    .A2(_06704_),
    .B1(_06706_),
    .X(net373));
 sky130_fd_sc_hd__a21bo_1 _11723_ (.A1(net483),
    .A2(_06704_),
    .B1_N(_06706_),
    .X(net372));
 sky130_fd_sc_hd__nor2_4 _11724_ (.A(_03821_),
    .B(_03873_),
    .Y(_06707_));
 sky130_fd_sc_hd__and2_2 _11725_ (.A(\core.fetchProgramCounter[0] ),
    .B(net1310),
    .X(net305));
 sky130_fd_sc_hd__and2_1 _11726_ (.A(\core.fetchProgramCounter[1] ),
    .B(net1310),
    .X(net316));
 sky130_fd_sc_hd__nor2_1 _11727_ (.A(_06625_),
    .B(_06650_),
    .Y(_06708_));
 sky130_fd_sc_hd__and3_4 _11728_ (.A(_06620_),
    .B(_06623_),
    .C(_06708_),
    .X(_06709_));
 sky130_fd_sc_hd__and2b_2 _11729_ (.A_N(net1310),
    .B(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__nand2b_1 _11730_ (.A_N(net1311),
    .B(_06709_),
    .Y(_06711_));
 sky130_fd_sc_hd__and2b_4 _11731_ (.A_N(_04885_),
    .B(_04886_),
    .X(_06712_));
 sky130_fd_sc_hd__xnor2_4 _11732_ (.A(_05054_),
    .B(_06712_),
    .Y(_06713_));
 sky130_fd_sc_hd__a22o_2 _11733_ (.A1(\core.fetchProgramCounter[2] ),
    .A2(net1312),
    .B1(net527),
    .B2(_06713_),
    .X(net325));
 sky130_fd_sc_hd__nor2_8 _11734_ (.A(_04804_),
    .B(_04806_),
    .Y(_06714_));
 sky130_fd_sc_hd__xnor2_4 _11735_ (.A(_05056_),
    .B(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__a22o_2 _11736_ (.A1(\core.fetchProgramCounter[3] ),
    .A2(net1312),
    .B1(net527),
    .B2(_06715_),
    .X(net326));
 sky130_fd_sc_hd__xor2_4 _11737_ (.A(_04724_),
    .B(_05058_),
    .X(_06716_));
 sky130_fd_sc_hd__a22o_1 _11738_ (.A1(\core.fetchProgramCounter[4] ),
    .A2(net1312),
    .B1(net527),
    .B2(_06716_),
    .X(net327));
 sky130_fd_sc_hd__xnor2_4 _11739_ (.A(_04635_),
    .B(_05059_),
    .Y(_06717_));
 sky130_fd_sc_hd__inv_6 _11740_ (.A(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__a22o_1 _11741_ (.A1(\core.fetchProgramCounter[5] ),
    .A2(net1312),
    .B1(net526),
    .B2(_06718_),
    .X(net328));
 sky130_fd_sc_hd__and2b_4 _11742_ (.A_N(_04548_),
    .B(_04549_),
    .X(_06719_));
 sky130_fd_sc_hd__xnor2_4 _11743_ (.A(_05060_),
    .B(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__a22o_1 _11744_ (.A1(\core.fetchProgramCounter[6] ),
    .A2(net1311),
    .B1(net526),
    .B2(_06720_),
    .X(net329));
 sky130_fd_sc_hd__nor2_8 _11745_ (.A(_04462_),
    .B(_04463_),
    .Y(_06721_));
 sky130_fd_sc_hd__xnor2_4 _11746_ (.A(_05062_),
    .B(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__a22o_2 _11747_ (.A1(\core.fetchProgramCounter[7] ),
    .A2(net1314),
    .B1(net529),
    .B2(_06722_),
    .X(net330));
 sky130_fd_sc_hd__xnor2_4 _11748_ (.A(_04391_),
    .B(_05064_),
    .Y(_06723_));
 sky130_fd_sc_hd__a22o_1 _11749_ (.A1(\core.fetchProgramCounter[8] ),
    .A2(net1311),
    .B1(net525),
    .B2(_06723_),
    .X(net331));
 sky130_fd_sc_hd__xnor2_4 _11750_ (.A(_04307_),
    .B(_05065_),
    .Y(_06724_));
 sky130_fd_sc_hd__clkinv_4 _11751_ (.A(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__a22o_1 _11752_ (.A1(\core.fetchProgramCounter[9] ),
    .A2(net1314),
    .B1(net528),
    .B2(_06725_),
    .X(net332));
 sky130_fd_sc_hd__xor2_4 _11753_ (.A(_04218_),
    .B(_05066_),
    .X(_06726_));
 sky130_fd_sc_hd__a22o_1 _11754_ (.A1(\core.fetchProgramCounter[10] ),
    .A2(net1310),
    .B1(net526),
    .B2(_06726_),
    .X(net306));
 sky130_fd_sc_hd__a22o_1 _11755_ (.A1(\core.fetchProgramCounter[11] ),
    .A2(net1311),
    .B1(net525),
    .B2(_05068_),
    .X(net307));
 sky130_fd_sc_hd__a22o_1 _11756_ (.A1(\core.fetchProgramCounter[12] ),
    .A2(net1314),
    .B1(net528),
    .B2(_06670_),
    .X(net308));
 sky130_fd_sc_hd__a22o_1 _11757_ (.A1(\core.fetchProgramCounter[13] ),
    .A2(net1314),
    .B1(net528),
    .B2(_06668_),
    .X(net309));
 sky130_fd_sc_hd__a22o_1 _11758_ (.A1(\core.fetchProgramCounter[14] ),
    .A2(net1314),
    .B1(net528),
    .B2(_06667_),
    .X(net310));
 sky130_fd_sc_hd__a22o_1 _11759_ (.A1(\core.fetchProgramCounter[15] ),
    .A2(net1314),
    .B1(net528),
    .B2(_06666_),
    .X(net311));
 sky130_fd_sc_hd__a22o_2 _11760_ (.A1(\core.fetchProgramCounter[16] ),
    .A2(net1313),
    .B1(net530),
    .B2(_06665_),
    .X(net312));
 sky130_fd_sc_hd__a22o_2 _11761_ (.A1(\core.fetchProgramCounter[17] ),
    .A2(net1313),
    .B1(net530),
    .B2(_06664_),
    .X(net313));
 sky130_fd_sc_hd__a22o_2 _11762_ (.A1(\core.fetchProgramCounter[18] ),
    .A2(net1313),
    .B1(net527),
    .B2(_06663_),
    .X(net314));
 sky130_fd_sc_hd__a22o_4 _11763_ (.A1(\core.fetchProgramCounter[19] ),
    .A2(net1313),
    .B1(net527),
    .B2(_06662_),
    .X(net315));
 sky130_fd_sc_hd__a22o_4 _11764_ (.A1(\core.fetchProgramCounter[20] ),
    .A2(net1313),
    .B1(net527),
    .B2(_06660_),
    .X(net317));
 sky130_fd_sc_hd__a22o_4 _11765_ (.A1(\core.fetchProgramCounter[21] ),
    .A2(net1313),
    .B1(net530),
    .B2(_06659_),
    .X(net318));
 sky130_fd_sc_hd__a22o_4 _11766_ (.A1(\core.fetchProgramCounter[22] ),
    .A2(net1313),
    .B1(net527),
    .B2(_06658_),
    .X(net319));
 sky130_fd_sc_hd__a22o_4 _11767_ (.A1(\core.fetchProgramCounter[23] ),
    .A2(net1313),
    .B1(net527),
    .B2(_06656_),
    .X(net320));
 sky130_fd_sc_hd__a22o_2 _11768_ (.A1(\core.fetchProgramCounter[24] ),
    .A2(net1310),
    .B1(net525),
    .B2(_06631_),
    .X(net321));
 sky130_fd_sc_hd__a22o_2 _11769_ (.A1(\core.fetchProgramCounter[25] ),
    .A2(net1310),
    .B1(net527),
    .B2(_06629_),
    .X(net322));
 sky130_fd_sc_hd__a22o_4 _11770_ (.A1(\core.fetchProgramCounter[26] ),
    .A2(net1313),
    .B1(net530),
    .B2(_06627_),
    .X(net323));
 sky130_fd_sc_hd__a2bb2o_4 _11771_ (.A1_N(_06626_),
    .A2_N(_06711_),
    .B1(net1311),
    .B2(\core.fetchProgramCounter[27] ),
    .X(net324));
 sky130_fd_sc_hd__a21o_1 _11772_ (.A1(net613),
    .A2(_06709_),
    .B1(net1310),
    .X(net366));
 sky130_fd_sc_hd__a21oi_1 _11773_ (.A1(net668),
    .A2(_06644_),
    .B1(net1043),
    .Y(_06727_));
 sky130_fd_sc_hd__and3_4 _11774_ (.A(net633),
    .B(_06649_),
    .C(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__a21o_1 _11775_ (.A1(_06709_),
    .A2(_06728_),
    .B1(net1310),
    .X(net367));
 sky130_fd_sc_hd__a21oi_4 _11776_ (.A1(_04972_),
    .A2(_06645_),
    .B1(net669),
    .Y(_06729_));
 sky130_fd_sc_hd__a211oi_4 _11777_ (.A1(_04053_),
    .A2(net611),
    .B1(_06650_),
    .C1(_06729_),
    .Y(_06730_));
 sky130_fd_sc_hd__a21o_1 _11778_ (.A1(_06709_),
    .A2(_06730_),
    .B1(net1310),
    .X(net368));
 sky130_fd_sc_hd__or2_1 _11779_ (.A(net633),
    .B(_06727_),
    .X(_06731_));
 sky130_fd_sc_hd__o211a_4 _11780_ (.A1(_06634_),
    .A2(net634),
    .B1(_06649_),
    .C1(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__a21o_1 _11781_ (.A1(_06709_),
    .A2(_06732_),
    .B1(net1310),
    .X(net369));
 sky130_fd_sc_hd__nor2_8 _11782_ (.A(net1043),
    .B(_05012_),
    .Y(_06733_));
 sky130_fd_sc_hd__nand2_1 _11783_ (.A(net669),
    .B(_06733_),
    .Y(_06734_));
 sky130_fd_sc_hd__and3_1 _11784_ (.A(net613),
    .B(net526),
    .C(_06733_),
    .X(net334));
 sky130_fd_sc_hd__nor2_8 _11785_ (.A(net1043),
    .B(_04930_),
    .Y(_06735_));
 sky130_fd_sc_hd__nand2_1 _11786_ (.A(net667),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__and3_1 _11787_ (.A(net613),
    .B(net526),
    .C(_06735_),
    .X(net345));
 sky130_fd_sc_hd__nor2_8 _11788_ (.A(net1043),
    .B(_04848_),
    .Y(_06737_));
 sky130_fd_sc_hd__and3_1 _11789_ (.A(net613),
    .B(net526),
    .C(_06737_),
    .X(net356));
 sky130_fd_sc_hd__nor4_2 _11790_ (.A(_04070_),
    .B(_04095_),
    .C(_04731_),
    .D(_04762_),
    .Y(_06738_));
 sky130_fd_sc_hd__nand2_1 _11791_ (.A(net667),
    .B(net989),
    .Y(_06739_));
 sky130_fd_sc_hd__and3_1 _11792_ (.A(net613),
    .B(net526),
    .C(net989),
    .X(net359));
 sky130_fd_sc_hd__nor2_8 _11793_ (.A(net1043),
    .B(_04682_),
    .Y(_06740_));
 sky130_fd_sc_hd__nand2_1 _11794_ (.A(net667),
    .B(_06740_),
    .Y(_06741_));
 sky130_fd_sc_hd__and3_1 _11795_ (.A(net613),
    .B(net526),
    .C(_06740_),
    .X(net360));
 sky130_fd_sc_hd__nor2_8 _11796_ (.A(net1043),
    .B(_04630_),
    .Y(_06742_));
 sky130_fd_sc_hd__and3_1 _11797_ (.A(net613),
    .B(net526),
    .C(_06742_),
    .X(net361));
 sky130_fd_sc_hd__nor2_8 _11798_ (.A(net1043),
    .B(_04545_),
    .Y(_06743_));
 sky130_fd_sc_hd__and3_1 _11799_ (.A(net613),
    .B(net526),
    .C(_06743_),
    .X(net362));
 sky130_fd_sc_hd__nand4_4 _11800_ (.A(_04071_),
    .B(net1239),
    .C(_04425_),
    .D(_04459_),
    .Y(_06744_));
 sky130_fd_sc_hd__nor2_8 _11801_ (.A(_06643_),
    .B(_06744_),
    .Y(_06745_));
 sky130_fd_sc_hd__and2_1 _11802_ (.A(net525),
    .B(_06745_),
    .X(net363));
 sky130_fd_sc_hd__nor2_2 _11803_ (.A(net667),
    .B(_06733_),
    .Y(_06746_));
 sky130_fd_sc_hd__or2_4 _11804_ (.A(_04352_),
    .B(_06646_),
    .X(_06747_));
 sky130_fd_sc_hd__a21oi_4 _11805_ (.A1(net667),
    .A2(_06747_),
    .B1(_06746_),
    .Y(_06748_));
 sky130_fd_sc_hd__and3_1 _11806_ (.A(net633),
    .B(net525),
    .C(_06748_),
    .X(net364));
 sky130_fd_sc_hd__nor2_2 _11807_ (.A(net667),
    .B(_06735_),
    .Y(_06749_));
 sky130_fd_sc_hd__or2_4 _11808_ (.A(_04266_),
    .B(_06646_),
    .X(_06750_));
 sky130_fd_sc_hd__a21oi_4 _11809_ (.A1(net667),
    .A2(_06750_),
    .B1(_06749_),
    .Y(_06751_));
 sky130_fd_sc_hd__and3_1 _11810_ (.A(net633),
    .B(net525),
    .C(_06751_),
    .X(net365));
 sky130_fd_sc_hd__nor2_2 _11811_ (.A(net669),
    .B(_06737_),
    .Y(_06752_));
 sky130_fd_sc_hd__or2_4 _11812_ (.A(_04178_),
    .B(_06646_),
    .X(_06753_));
 sky130_fd_sc_hd__a21oi_4 _11813_ (.A1(net669),
    .A2(_06753_),
    .B1(_06752_),
    .Y(_06754_));
 sky130_fd_sc_hd__and3_1 _11814_ (.A(_06641_),
    .B(net525),
    .C(_06754_),
    .X(net335));
 sky130_fd_sc_hd__nor2_4 _11815_ (.A(net668),
    .B(net989),
    .Y(_06755_));
 sky130_fd_sc_hd__or3b_4 _11816_ (.A(net1043),
    .B(_06644_),
    .C_N(_04127_),
    .X(_06756_));
 sky130_fd_sc_hd__a21oi_4 _11817_ (.A1(net668),
    .A2(_06756_),
    .B1(_06755_),
    .Y(_06757_));
 sky130_fd_sc_hd__and3_1 _11818_ (.A(_06641_),
    .B(net525),
    .C(_06757_),
    .X(net336));
 sky130_fd_sc_hd__or2_4 _11819_ (.A(_06475_),
    .B(_06646_),
    .X(_06758_));
 sky130_fd_sc_hd__nor2_2 _11820_ (.A(net667),
    .B(_06740_),
    .Y(_06759_));
 sky130_fd_sc_hd__a211oi_4 _11821_ (.A1(net667),
    .A2(_06758_),
    .B1(_06759_),
    .C1(net634),
    .Y(_06760_));
 sky130_fd_sc_hd__and2_1 _11822_ (.A(net528),
    .B(_06760_),
    .X(net337));
 sky130_fd_sc_hd__nor2_1 _11823_ (.A(_06398_),
    .B(_06646_),
    .Y(_06761_));
 sky130_fd_sc_hd__or2_2 _11824_ (.A(net671),
    .B(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__nor2_1 _11825_ (.A(_06638_),
    .B(_06742_),
    .Y(_06763_));
 sky130_fd_sc_hd__nor2_1 _11826_ (.A(net635),
    .B(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__and3_4 _11827_ (.A(net531),
    .B(_06762_),
    .C(_06764_),
    .X(net338));
 sky130_fd_sc_hd__or2_4 _11828_ (.A(_06321_),
    .B(_06646_),
    .X(_06765_));
 sky130_fd_sc_hd__nor2_2 _11829_ (.A(net668),
    .B(_06743_),
    .Y(_06766_));
 sky130_fd_sc_hd__a211oi_4 _11830_ (.A1(net668),
    .A2(_06765_),
    .B1(_06766_),
    .C1(net634),
    .Y(_06767_));
 sky130_fd_sc_hd__and2_1 _11831_ (.A(net528),
    .B(_06767_),
    .X(net339));
 sky130_fd_sc_hd__nor2_2 _11832_ (.A(_06245_),
    .B(_06646_),
    .Y(_06768_));
 sky130_fd_sc_hd__clkinv_2 _11833_ (.A(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__nand2_1 _11834_ (.A(net670),
    .B(_06744_),
    .Y(_06770_));
 sky130_fd_sc_hd__o211a_4 _11835_ (.A1(net670),
    .A2(_06768_),
    .B1(_06770_),
    .C1(net633),
    .X(_06771_));
 sky130_fd_sc_hd__and2_1 _11836_ (.A(net528),
    .B(_06771_),
    .X(net340));
 sky130_fd_sc_hd__or2_4 _11837_ (.A(_06167_),
    .B(net990),
    .X(_06772_));
 sky130_fd_sc_hd__a22o_1 _11838_ (.A1(net634),
    .A2(_06734_),
    .B1(_06747_),
    .B2(net670),
    .X(_06773_));
 sky130_fd_sc_hd__a21oi_4 _11839_ (.A1(net611),
    .A2(_06772_),
    .B1(_06773_),
    .Y(_06774_));
 sky130_fd_sc_hd__and2_1 _11840_ (.A(net528),
    .B(_06774_),
    .X(net341));
 sky130_fd_sc_hd__or2_2 _11841_ (.A(_06090_),
    .B(net990),
    .X(_06775_));
 sky130_fd_sc_hd__a22o_2 _11842_ (.A1(net634),
    .A2(_06736_),
    .B1(_06750_),
    .B2(net670),
    .X(_06776_));
 sky130_fd_sc_hd__a21oi_4 _11843_ (.A1(net610),
    .A2(_06775_),
    .B1(_06776_),
    .Y(_06777_));
 sky130_fd_sc_hd__and2_1 _11844_ (.A(net528),
    .B(_06777_),
    .X(net342));
 sky130_fd_sc_hd__or2_2 _11845_ (.A(_06012_),
    .B(net991),
    .X(_06778_));
 sky130_fd_sc_hd__nand2_1 _11846_ (.A(_06638_),
    .B(_06737_),
    .Y(_06779_));
 sky130_fd_sc_hd__a22o_1 _11847_ (.A1(net671),
    .A2(_06753_),
    .B1(_06779_),
    .B2(net635),
    .X(_06780_));
 sky130_fd_sc_hd__a21oi_4 _11848_ (.A1(net610),
    .A2(_06778_),
    .B1(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__and2_1 _11849_ (.A(net529),
    .B(_06781_),
    .X(net343));
 sky130_fd_sc_hd__or2_4 _11850_ (.A(_05936_),
    .B(net990),
    .X(_06782_));
 sky130_fd_sc_hd__o211a_1 _11851_ (.A1(net634),
    .A2(_06756_),
    .B1(_06739_),
    .C1(_06643_),
    .X(_06783_));
 sky130_fd_sc_hd__a21oi_4 _11852_ (.A1(net610),
    .A2(_06782_),
    .B1(_06783_),
    .Y(_06784_));
 sky130_fd_sc_hd__and2_1 _11853_ (.A(net529),
    .B(_06784_),
    .X(net344));
 sky130_fd_sc_hd__or2_2 _11854_ (.A(_05860_),
    .B(net990),
    .X(_06785_));
 sky130_fd_sc_hd__o211a_1 _11855_ (.A1(net634),
    .A2(_06758_),
    .B1(_06741_),
    .C1(_06643_),
    .X(_06786_));
 sky130_fd_sc_hd__a21oi_4 _11856_ (.A1(net610),
    .A2(_06785_),
    .B1(_06786_),
    .Y(_06787_));
 sky130_fd_sc_hd__and2_1 _11857_ (.A(net529),
    .B(_06787_),
    .X(net346));
 sky130_fd_sc_hd__or2_1 _11858_ (.A(net669),
    .B(_06761_),
    .X(_06788_));
 sky130_fd_sc_hd__nand2_8 _11859_ (.A(net669),
    .B(net634),
    .Y(_06789_));
 sky130_fd_sc_hd__or2_2 _11860_ (.A(_05780_),
    .B(net990),
    .X(_06790_));
 sky130_fd_sc_hd__a21oi_1 _11861_ (.A1(net669),
    .A2(_06790_),
    .B1(net635),
    .Y(_06791_));
 sky130_fd_sc_hd__a31o_1 _11862_ (.A1(_06638_),
    .A2(net635),
    .A3(_06742_),
    .B1(_06791_),
    .X(_06792_));
 sky130_fd_sc_hd__and3_4 _11863_ (.A(net531),
    .B(_06788_),
    .C(_06792_),
    .X(net347));
 sky130_fd_sc_hd__or2_2 _11864_ (.A(_05702_),
    .B(net990),
    .X(_06793_));
 sky130_fd_sc_hd__nand2_1 _11865_ (.A(net668),
    .B(_06743_),
    .Y(_06794_));
 sky130_fd_sc_hd__a22o_1 _11866_ (.A1(net670),
    .A2(_06765_),
    .B1(_06794_),
    .B2(net634),
    .X(_06795_));
 sky130_fd_sc_hd__a21oi_4 _11867_ (.A1(net610),
    .A2(_06793_),
    .B1(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__and2_1 _11868_ (.A(net529),
    .B(_06796_),
    .X(net348));
 sky130_fd_sc_hd__nand2_2 _11869_ (.A(_05626_),
    .B(_06634_),
    .Y(_06797_));
 sky130_fd_sc_hd__o21a_1 _11870_ (.A1(net670),
    .A2(_06744_),
    .B1(net634),
    .X(_06798_));
 sky130_fd_sc_hd__a221oi_4 _11871_ (.A1(net670),
    .A2(_06769_),
    .B1(_06797_),
    .B2(net610),
    .C1(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__and2_1 _11872_ (.A(net529),
    .B(_06799_),
    .X(net349));
 sky130_fd_sc_hd__o21ai_2 _11873_ (.A1(_05551_),
    .A2(net990),
    .B1(net612),
    .Y(_06800_));
 sky130_fd_sc_hd__nand2_8 _11874_ (.A(_04972_),
    .B(net670),
    .Y(_06801_));
 sky130_fd_sc_hd__nand2_8 _11875_ (.A(_06789_),
    .B(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__o22a_1 _11876_ (.A1(_06747_),
    .A2(_06789_),
    .B1(_06801_),
    .B2(_06772_),
    .X(_06803_));
 sky130_fd_sc_hd__o21ai_2 _11877_ (.A1(_06746_),
    .A2(_06802_),
    .B1(_06803_),
    .Y(_06804_));
 sky130_fd_sc_hd__and3_4 _11878_ (.A(net531),
    .B(_06800_),
    .C(_06804_),
    .X(net350));
 sky130_fd_sc_hd__o21ai_2 _11879_ (.A1(_05476_),
    .A2(net990),
    .B1(net612),
    .Y(_06805_));
 sky130_fd_sc_hd__o22a_1 _11880_ (.A1(_06750_),
    .A2(_06789_),
    .B1(_06801_),
    .B2(_06775_),
    .X(_06806_));
 sky130_fd_sc_hd__o21ai_2 _11881_ (.A1(_06749_),
    .A2(_06802_),
    .B1(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__and3_4 _11882_ (.A(net531),
    .B(_06805_),
    .C(_06807_),
    .X(net351));
 sky130_fd_sc_hd__o21ai_2 _11883_ (.A1(_05402_),
    .A2(net990),
    .B1(net611),
    .Y(_06808_));
 sky130_fd_sc_hd__o22a_1 _11884_ (.A1(_06753_),
    .A2(_06789_),
    .B1(_06801_),
    .B2(_06778_),
    .X(_06809_));
 sky130_fd_sc_hd__o21ai_2 _11885_ (.A1(_06752_),
    .A2(_06802_),
    .B1(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__and3_4 _11886_ (.A(net531),
    .B(_06808_),
    .C(_06810_),
    .X(net352));
 sky130_fd_sc_hd__o21ai_2 _11887_ (.A1(_05329_),
    .A2(net991),
    .B1(net611),
    .Y(_06811_));
 sky130_fd_sc_hd__o22a_1 _11888_ (.A1(_06756_),
    .A2(_06789_),
    .B1(_06801_),
    .B2(_06782_),
    .X(_06812_));
 sky130_fd_sc_hd__o21ai_4 _11889_ (.A1(_06755_),
    .A2(_06802_),
    .B1(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__and3_4 _11890_ (.A(net531),
    .B(_06811_),
    .C(_06813_),
    .X(net353));
 sky130_fd_sc_hd__o21ai_2 _11891_ (.A1(_05258_),
    .A2(net990),
    .B1(net610),
    .Y(_06814_));
 sky130_fd_sc_hd__o22a_1 _11892_ (.A1(_06758_),
    .A2(_06789_),
    .B1(_06801_),
    .B2(_06785_),
    .X(_06815_));
 sky130_fd_sc_hd__o21ai_2 _11893_ (.A1(_06759_),
    .A2(_06802_),
    .B1(_06815_),
    .Y(_06816_));
 sky130_fd_sc_hd__and3_4 _11894_ (.A(net531),
    .B(_06814_),
    .C(_06816_),
    .X(net354));
 sky130_fd_sc_hd__o21ai_2 _11895_ (.A1(_05183_),
    .A2(net991),
    .B1(net610),
    .Y(_06817_));
 sky130_fd_sc_hd__or2_1 _11896_ (.A(_06790_),
    .B(_06801_),
    .X(_06818_));
 sky130_fd_sc_hd__o31a_1 _11897_ (.A1(_06398_),
    .A2(_06646_),
    .A3(_06789_),
    .B1(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__o21ai_2 _11898_ (.A1(_06763_),
    .A2(_06802_),
    .B1(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__and3_4 _11899_ (.A(net531),
    .B(_06817_),
    .C(_06820_),
    .X(net355));
 sky130_fd_sc_hd__o21a_2 _11900_ (.A1(_05108_),
    .A2(net991),
    .B1(net610),
    .X(_06821_));
 sky130_fd_sc_hd__or2_1 _11901_ (.A(_06793_),
    .B(_06801_),
    .X(_06822_));
 sky130_fd_sc_hd__o221a_4 _11902_ (.A1(_06765_),
    .A2(_06789_),
    .B1(_06802_),
    .B2(_06766_),
    .C1(_06822_),
    .X(_06823_));
 sky130_fd_sc_hd__nor2_8 _11903_ (.A(_06821_),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__and2_1 _11904_ (.A(net529),
    .B(_06824_),
    .X(net357));
 sky130_fd_sc_hd__a21oi_4 _11905_ (.A1(_06579_),
    .A2(_06634_),
    .B1(_06643_),
    .Y(_06825_));
 sky130_fd_sc_hd__a21o_1 _11906_ (.A1(net670),
    .A2(_06744_),
    .B1(_06802_),
    .X(_06826_));
 sky130_fd_sc_hd__o221a_4 _11907_ (.A1(_06769_),
    .A2(_06789_),
    .B1(_06797_),
    .B2(_06801_),
    .C1(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__nor2_8 _11908_ (.A(_06825_),
    .B(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__and2_1 _11909_ (.A(net529),
    .B(_06828_),
    .X(net358));
 sky130_fd_sc_hd__a22o_4 _11910_ (.A1(\core.fetchProgramCounter[2] ),
    .A2(net1601),
    .B1(net532),
    .B2(_06713_),
    .X(net294));
 sky130_fd_sc_hd__a22o_4 _11911_ (.A1(\core.fetchProgramCounter[3] ),
    .A2(net1601),
    .B1(net532),
    .B2(_06715_),
    .X(net295));
 sky130_fd_sc_hd__a22o_4 _11912_ (.A1(\core.fetchProgramCounter[4] ),
    .A2(net1601),
    .B1(net532),
    .B2(_06716_),
    .X(net296));
 sky130_fd_sc_hd__a22o_4 _11913_ (.A1(\core.fetchProgramCounter[5] ),
    .A2(net1602),
    .B1(net532),
    .B2(_06718_),
    .X(net297));
 sky130_fd_sc_hd__a22o_4 _11914_ (.A1(\core.fetchProgramCounter[6] ),
    .A2(net1602),
    .B1(net532),
    .B2(_06720_),
    .X(net298));
 sky130_fd_sc_hd__a22o_4 _11915_ (.A1(\core.fetchProgramCounter[7] ),
    .A2(net1602),
    .B1(net532),
    .B2(_06722_),
    .X(net299));
 sky130_fd_sc_hd__a22o_4 _11916_ (.A1(\core.fetchProgramCounter[8] ),
    .A2(net1602),
    .B1(net532),
    .B2(_06723_),
    .X(net300));
 sky130_fd_sc_hd__a22o_4 _11917_ (.A1(\core.fetchProgramCounter[9] ),
    .A2(net1602),
    .B1(net532),
    .B2(_06725_),
    .X(net301));
 sky130_fd_sc_hd__a22o_4 _11918_ (.A1(\core.fetchProgramCounter[10] ),
    .A2(net1602),
    .B1(_06652_),
    .B2(_06726_),
    .X(net302));
 sky130_fd_sc_hd__and3b_1 _11919_ (.A_N(net505),
    .B(net1236),
    .C(_06702_),
    .X(_06829_));
 sky130_fd_sc_hd__a32o_4 _11920_ (.A1(net612),
    .A2(net501),
    .A3(_06733_),
    .B1(net495),
    .B2(net215),
    .X(net376));
 sky130_fd_sc_hd__a32o_4 _11921_ (.A1(net612),
    .A2(net501),
    .A3(_06735_),
    .B1(net495),
    .B2(net226),
    .X(net387));
 sky130_fd_sc_hd__a32o_4 _11922_ (.A1(net612),
    .A2(net501),
    .A3(_06737_),
    .B1(net495),
    .B2(net237),
    .X(net398));
 sky130_fd_sc_hd__a32o_4 _11923_ (.A1(net612),
    .A2(net501),
    .A3(net989),
    .B1(net495),
    .B2(net240),
    .X(net401));
 sky130_fd_sc_hd__a32o_4 _11924_ (.A1(net612),
    .A2(net501),
    .A3(_06740_),
    .B1(net495),
    .B2(net241),
    .X(net402));
 sky130_fd_sc_hd__a32o_4 _11925_ (.A1(net612),
    .A2(net501),
    .A3(_06742_),
    .B1(net495),
    .B2(net242),
    .X(net403));
 sky130_fd_sc_hd__a32o_4 _11926_ (.A1(net612),
    .A2(net501),
    .A3(_06743_),
    .B1(net495),
    .B2(net243),
    .X(net404));
 sky130_fd_sc_hd__a22o_4 _11927_ (.A1(net503),
    .A2(_06745_),
    .B1(net495),
    .B2(net244),
    .X(net405));
 sky130_fd_sc_hd__a32o_4 _11928_ (.A1(net633),
    .A2(net502),
    .A3(_06748_),
    .B1(net496),
    .B2(net245),
    .X(net406));
 sky130_fd_sc_hd__a32o_4 _11929_ (.A1(net633),
    .A2(net502),
    .A3(_06751_),
    .B1(net496),
    .B2(net246),
    .X(net407));
 sky130_fd_sc_hd__a32o_4 _11930_ (.A1(net633),
    .A2(net502),
    .A3(_06754_),
    .B1(net496),
    .B2(net216),
    .X(net377));
 sky130_fd_sc_hd__a32o_4 _11931_ (.A1(net633),
    .A2(net502),
    .A3(_06757_),
    .B1(net496),
    .B2(net217),
    .X(net378));
 sky130_fd_sc_hd__a22o_4 _11932_ (.A1(net501),
    .A2(_06760_),
    .B1(net495),
    .B2(net218),
    .X(net379));
 sky130_fd_sc_hd__a32o_4 _11933_ (.A1(net504),
    .A2(_06762_),
    .A3(_06764_),
    .B1(net498),
    .B2(net219),
    .X(net380));
 sky130_fd_sc_hd__a22o_2 _11934_ (.A1(net501),
    .A2(_06767_),
    .B1(net499),
    .B2(net220),
    .X(net381));
 sky130_fd_sc_hd__a22o_4 _11935_ (.A1(net503),
    .A2(_06771_),
    .B1(net495),
    .B2(net221),
    .X(net382));
 sky130_fd_sc_hd__a22o_4 _11936_ (.A1(net504),
    .A2(_06774_),
    .B1(net498),
    .B2(net222),
    .X(net383));
 sky130_fd_sc_hd__a22o_4 _11937_ (.A1(net503),
    .A2(_06777_),
    .B1(net497),
    .B2(net223),
    .X(net384));
 sky130_fd_sc_hd__a22o_4 _11938_ (.A1(net505),
    .A2(_06781_),
    .B1(net498),
    .B2(net224),
    .X(net385));
 sky130_fd_sc_hd__a22o_2 _11939_ (.A1(net501),
    .A2(_06784_),
    .B1(net497),
    .B2(net225),
    .X(net386));
 sky130_fd_sc_hd__a22o_2 _11940_ (.A1(net502),
    .A2(_06787_),
    .B1(net497),
    .B2(net227),
    .X(net388));
 sky130_fd_sc_hd__a32o_4 _11941_ (.A1(net505),
    .A2(_06788_),
    .A3(_06792_),
    .B1(net498),
    .B2(net228),
    .X(net389));
 sky130_fd_sc_hd__a22o_2 _11942_ (.A1(net502),
    .A2(_06796_),
    .B1(net496),
    .B2(net229),
    .X(net390));
 sky130_fd_sc_hd__a22o_2 _11943_ (.A1(net502),
    .A2(_06799_),
    .B1(net496),
    .B2(net230),
    .X(net391));
 sky130_fd_sc_hd__a32o_4 _11944_ (.A1(net502),
    .A2(_06800_),
    .A3(_06804_),
    .B1(net496),
    .B2(net231),
    .X(net392));
 sky130_fd_sc_hd__a32o_4 _11945_ (.A1(net503),
    .A2(_06805_),
    .A3(_06807_),
    .B1(net497),
    .B2(net232),
    .X(net393));
 sky130_fd_sc_hd__a32o_4 _11946_ (.A1(net504),
    .A2(_06808_),
    .A3(_06810_),
    .B1(net498),
    .B2(net233),
    .X(net394));
 sky130_fd_sc_hd__a32o_4 _11947_ (.A1(net505),
    .A2(_06811_),
    .A3(_06813_),
    .B1(net498),
    .B2(net234),
    .X(net395));
 sky130_fd_sc_hd__a32o_4 _11948_ (.A1(net504),
    .A2(_06814_),
    .A3(_06816_),
    .B1(net498),
    .B2(net235),
    .X(net396));
 sky130_fd_sc_hd__a32o_4 _11949_ (.A1(net505),
    .A2(_06817_),
    .A3(_06820_),
    .B1(net499),
    .B2(net236),
    .X(net397));
 sky130_fd_sc_hd__a22o_2 _11950_ (.A1(net504),
    .A2(_06824_),
    .B1(net498),
    .B2(net238),
    .X(net399));
 sky130_fd_sc_hd__a22o_2 _11951_ (.A1(net504),
    .A2(_06828_),
    .B1(net498),
    .B2(net239),
    .X(net400));
 sky130_fd_sc_hd__a31o_1 _11952_ (.A1(_06633_),
    .A2(net610),
    .A3(_06649_),
    .B1(net1601),
    .X(_06830_));
 sky130_fd_sc_hd__a22o_4 _11953_ (.A1(\wbSRAMInterface.currentByteSelect[0] ),
    .A2(net498),
    .B1(_06830_),
    .B2(net504),
    .X(net484));
 sky130_fd_sc_hd__a21o_1 _11954_ (.A1(_06633_),
    .A2(_06728_),
    .B1(net1601),
    .X(_06831_));
 sky130_fd_sc_hd__a22o_4 _11955_ (.A1(\wbSRAMInterface.currentByteSelect[1] ),
    .A2(net496),
    .B1(_06831_),
    .B2(net503),
    .X(net485));
 sky130_fd_sc_hd__a21o_1 _11956_ (.A1(_06633_),
    .A2(_06730_),
    .B1(net1601),
    .X(_06832_));
 sky130_fd_sc_hd__a22o_4 _11957_ (.A1(\wbSRAMInterface.currentByteSelect[2] ),
    .A2(net496),
    .B1(_06832_),
    .B2(net503),
    .X(net486));
 sky130_fd_sc_hd__a21o_1 _11958_ (.A1(_06633_),
    .A2(_06732_),
    .B1(net1601),
    .X(_06833_));
 sky130_fd_sc_hd__a22o_4 _11959_ (.A1(\wbSRAMInterface.currentByteSelect[3] ),
    .A2(net496),
    .B1(_06833_),
    .B2(net503),
    .X(net487));
 sky130_fd_sc_hd__a22o_4 _11960_ (.A1(\wbSRAMInterface.currentAddress[2] ),
    .A2(_06705_),
    .B1(net294),
    .B2(_06692_),
    .X(net285));
 sky130_fd_sc_hd__a22o_4 _11961_ (.A1(\wbSRAMInterface.currentAddress[3] ),
    .A2(_06705_),
    .B1(net295),
    .B2(net500),
    .X(net286));
 sky130_fd_sc_hd__a22o_4 _11962_ (.A1(\wbSRAMInterface.currentAddress[4] ),
    .A2(_06705_),
    .B1(net296),
    .B2(net500),
    .X(net287));
 sky130_fd_sc_hd__a22o_4 _11963_ (.A1(\wbSRAMInterface.currentAddress[5] ),
    .A2(_06705_),
    .B1(net297),
    .B2(_06692_),
    .X(net288));
 sky130_fd_sc_hd__a22o_4 _11964_ (.A1(\wbSRAMInterface.currentAddress[6] ),
    .A2(_06705_),
    .B1(net298),
    .B2(net500),
    .X(net289));
 sky130_fd_sc_hd__a22o_4 _11965_ (.A1(\wbSRAMInterface.currentAddress[7] ),
    .A2(_06705_),
    .B1(net299),
    .B2(net500),
    .X(net290));
 sky130_fd_sc_hd__a22o_4 _11966_ (.A1(\wbSRAMInterface.currentAddress[8] ),
    .A2(_06705_),
    .B1(net300),
    .B2(net500),
    .X(net291));
 sky130_fd_sc_hd__a22o_4 _11967_ (.A1(\wbSRAMInterface.currentAddress[9] ),
    .A2(_06705_),
    .B1(net301),
    .B2(net500),
    .X(net292));
 sky130_fd_sc_hd__a22o_4 _11968_ (.A1(\wbSRAMInterface.currentAddress[10] ),
    .A2(_06705_),
    .B1(net302),
    .B2(net500),
    .X(net293));
 sky130_fd_sc_hd__nand2_4 _11969_ (.A(\jtag.state[1] ),
    .B(net1721),
    .Y(_06834_));
 sky130_fd_sc_hd__and3_4 _11970_ (.A(\jtag.state[3] ),
    .B(_03818_),
    .C(net1720),
    .X(_06835_));
 sky130_fd_sc_hd__nand2_1 _11971_ (.A(net446),
    .B(net445),
    .Y(_06836_));
 sky130_fd_sc_hd__or4_4 _11972_ (.A(net449),
    .B(net448),
    .C(net447),
    .D(_06836_),
    .X(_06837_));
 sky130_fd_sc_hd__or4b_1 _11973_ (.A(net449),
    .B(net446),
    .C(net445),
    .D_N(net447),
    .X(_06838_));
 sky130_fd_sc_hd__o21a_2 _11974_ (.A1(net448),
    .A2(_06838_),
    .B1(_06837_),
    .X(_06839_));
 sky130_fd_sc_hd__and3_1 _11975_ (.A(net447),
    .B(net446),
    .C(net445),
    .X(_06840_));
 sky130_fd_sc_hd__and3_1 _11976_ (.A(net449),
    .B(net448),
    .C(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__or3b_1 _11977_ (.A(_06839_),
    .B(_06841_),
    .C_N(\jtag.dataIDRegister.data[31] ),
    .X(_06842_));
 sky130_fd_sc_hd__or3b_2 _11978_ (.A(net448),
    .B(net447),
    .C_N(net445),
    .X(_06843_));
 sky130_fd_sc_hd__nor3_4 _11979_ (.A(net449),
    .B(net446),
    .C(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__a21bo_1 _11980_ (.A1(\jtag.dataBypassRegister.data ),
    .A2(_06841_),
    .B1_N(_06842_),
    .X(_06845_));
 sky130_fd_sc_hd__or2_2 _11981_ (.A(\jtag.state[3] ),
    .B(_03818_),
    .X(_06846_));
 sky130_fd_sc_hd__nor3_4 _11982_ (.A(net1720),
    .B(net1721),
    .C(_06846_),
    .Y(_06847_));
 sky130_fd_sc_hd__mux2_1 _11983_ (.A0(_06845_),
    .A1(\jtag.dataBSRRegister.data[31] ),
    .S(_06844_),
    .X(_06848_));
 sky130_fd_sc_hd__a32o_4 _11984_ (.A1(\jtag.state[0] ),
    .A2(\jtag.instructionRegister.data[4] ),
    .A3(_06835_),
    .B1(_06847_),
    .B2(_06848_),
    .X(net408));
 sky130_fd_sc_hd__or4b_4 _11985_ (.A(_03828_),
    .B(net1906),
    .C(_03912_),
    .D_N(_03936_),
    .X(_06849_));
 sky130_fd_sc_hd__or2_4 _11986_ (.A(_03911_),
    .B(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__nor2_8 _11987_ (.A(_03910_),
    .B(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__or2_4 _11988_ (.A(_03910_),
    .B(_06850_),
    .X(_06852_));
 sky130_fd_sc_hd__or3_4 _11989_ (.A(\core.csr.currentInstruction[10] ),
    .B(net1801),
    .C(_03905_),
    .X(_06853_));
 sky130_fd_sc_hd__nor2_8 _11990_ (.A(_06852_),
    .B(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__mux2_1 _11991_ (.A0(\core.registers[19][0] ),
    .A1(net1078),
    .S(net827),
    .X(_00000_));
 sky130_fd_sc_hd__mux2_1 _11992_ (.A0(\core.registers[19][1] ),
    .A1(net1082),
    .S(net829),
    .X(_00001_));
 sky130_fd_sc_hd__mux2_1 _11993_ (.A0(\core.registers[19][2] ),
    .A1(net1085),
    .S(net827),
    .X(_00002_));
 sky130_fd_sc_hd__mux2_1 _11994_ (.A0(\core.registers[19][3] ),
    .A1(net1090),
    .S(net826),
    .X(_00003_));
 sky130_fd_sc_hd__mux2_1 _11995_ (.A0(\core.registers[19][4] ),
    .A1(net1028),
    .S(net829),
    .X(_00004_));
 sky130_fd_sc_hd__mux2_1 _11996_ (.A0(\core.registers[19][5] ),
    .A1(net1033),
    .S(net829),
    .X(_00005_));
 sky130_fd_sc_hd__mux2_1 _11997_ (.A0(\core.registers[19][6] ),
    .A1(net1037),
    .S(net829),
    .X(_00006_));
 sky130_fd_sc_hd__mux2_1 _11998_ (.A0(\core.registers[19][7] ),
    .A1(net1138),
    .S(net829),
    .X(_00007_));
 sky130_fd_sc_hd__mux2_1 _11999_ (.A0(\core.registers[19][8] ),
    .A1(net898),
    .S(net828),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _12000_ (.A0(\core.registers[19][9] ),
    .A1(net900),
    .S(net828),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _12001_ (.A0(\core.registers[19][10] ),
    .A1(net760),
    .S(net828),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _12002_ (.A0(\core.registers[19][11] ),
    .A1(net761),
    .S(net828),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _12003_ (.A0(\core.registers[19][12] ),
    .A1(net729),
    .S(net829),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _12004_ (.A0(\core.registers[19][13] ),
    .A1(net733),
    .S(net828),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _12005_ (.A0(\core.registers[19][14] ),
    .A1(net738),
    .S(net826),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _12006_ (.A0(\core.registers[19][15] ),
    .A1(net742),
    .S(net827),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _12007_ (.A0(\core.registers[19][16] ),
    .A1(net830),
    .S(net827),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _12008_ (.A0(\core.registers[19][17] ),
    .A1(net834),
    .S(net826),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _12009_ (.A0(\core.registers[19][18] ),
    .A1(net838),
    .S(net828),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _12010_ (.A0(\core.registers[19][19] ),
    .A1(net842),
    .S(net826),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _12011_ (.A0(\core.registers[19][20] ),
    .A1(net848),
    .S(net826),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _12012_ (.A0(\core.registers[19][21] ),
    .A1(net852),
    .S(net826),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _12013_ (.A0(\core.registers[19][22] ),
    .A1(net857),
    .S(net827),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _12014_ (.A0(\core.registers[19][23] ),
    .A1(net862),
    .S(net826),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _12015_ (.A0(\core.registers[19][24] ),
    .A1(net994),
    .S(net826),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _12016_ (.A0(\core.registers[19][25] ),
    .A1(net998),
    .S(net826),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _12017_ (.A0(\core.registers[19][26] ),
    .A1(net1002),
    .S(net828),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _12018_ (.A0(\core.registers[19][27] ),
    .A1(net866),
    .S(net828),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _12019_ (.A0(\core.registers[19][28] ),
    .A1(net871),
    .S(net829),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _12020_ (.A0(\core.registers[19][29] ),
    .A1(net874),
    .S(net828),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _12021_ (.A0(\core.registers[19][30] ),
    .A1(net878),
    .S(net828),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _12022_ (.A0(\core.registers[19][31] ),
    .A1(net1023),
    .S(net826),
    .X(_00031_));
 sky130_fd_sc_hd__nor2_1 _12023_ (.A(net1633),
    .B(net597),
    .Y(_06855_));
 sky130_fd_sc_hd__nand2_2 _12024_ (.A(net1632),
    .B(net602),
    .Y(_06856_));
 sky130_fd_sc_hd__or2_1 _12025_ (.A(\core.csr.currentInstruction[0] ),
    .B(net588),
    .X(_06857_));
 sky130_fd_sc_hd__o211a_1 _12026_ (.A1(\core.pipe0_currentInstruction[0] ),
    .A2(net584),
    .B1(_06857_),
    .C1(net1822),
    .X(_00032_));
 sky130_fd_sc_hd__or2_1 _12027_ (.A(\core.csr.currentInstruction[1] ),
    .B(net588),
    .X(_06858_));
 sky130_fd_sc_hd__o211a_1 _12028_ (.A1(\core.pipe0_currentInstruction[1] ),
    .A2(net585),
    .B1(_06858_),
    .C1(net1835),
    .X(_00033_));
 sky130_fd_sc_hd__nand2_1 _12029_ (.A(_03848_),
    .B(net585),
    .Y(_06859_));
 sky130_fd_sc_hd__o211a_1 _12030_ (.A1(\core.pipe0_currentInstruction[2] ),
    .A2(net585),
    .B1(_06859_),
    .C1(net1834),
    .X(_00034_));
 sky130_fd_sc_hd__or2_1 _12031_ (.A(\core.csr.currentInstruction[3] ),
    .B(net591),
    .X(_06860_));
 sky130_fd_sc_hd__o211a_1 _12032_ (.A1(\core.pipe0_currentInstruction[3] ),
    .A2(net585),
    .B1(_06860_),
    .C1(net1835),
    .X(_00035_));
 sky130_fd_sc_hd__or2_1 _12033_ (.A(\core.csr.currentInstruction[4] ),
    .B(net588),
    .X(_06861_));
 sky130_fd_sc_hd__o211a_1 _12034_ (.A1(\core.pipe0_currentInstruction[4] ),
    .A2(net584),
    .B1(_06861_),
    .C1(net1834),
    .X(_00036_));
 sky130_fd_sc_hd__nand2_1 _12035_ (.A(_03847_),
    .B(net585),
    .Y(_06862_));
 sky130_fd_sc_hd__o211a_1 _12036_ (.A1(\core.pipe0_currentInstruction[5] ),
    .A2(net584),
    .B1(_06862_),
    .C1(net1834),
    .X(_00037_));
 sky130_fd_sc_hd__or2_1 _12037_ (.A(\core.csr.currentInstruction[6] ),
    .B(net588),
    .X(_06863_));
 sky130_fd_sc_hd__o211a_1 _12038_ (.A1(\core.pipe0_currentInstruction[6] ),
    .A2(net585),
    .B1(_06863_),
    .C1(net1834),
    .X(_00038_));
 sky130_fd_sc_hd__or2_1 _12039_ (.A(\core.csr.currentInstruction[7] ),
    .B(net588),
    .X(_06864_));
 sky130_fd_sc_hd__o211a_1 _12040_ (.A1(\core.pipe0_currentInstruction[7] ),
    .A2(net584),
    .B1(_06864_),
    .C1(net1821),
    .X(_00039_));
 sky130_fd_sc_hd__or2_1 _12041_ (.A(\core.csr.currentInstruction[8] ),
    .B(net588),
    .X(_06865_));
 sky130_fd_sc_hd__o211a_1 _12042_ (.A1(\core.pipe0_currentInstruction[8] ),
    .A2(net584),
    .B1(_06865_),
    .C1(net1821),
    .X(_00040_));
 sky130_fd_sc_hd__or2_1 _12043_ (.A(net1801),
    .B(net588),
    .X(_06866_));
 sky130_fd_sc_hd__o211a_1 _12044_ (.A1(\core.pipe0_currentInstruction[9] ),
    .A2(net584),
    .B1(_06866_),
    .C1(net1821),
    .X(_00041_));
 sky130_fd_sc_hd__or2_1 _12045_ (.A(\core.csr.currentInstruction[10] ),
    .B(net588),
    .X(_06867_));
 sky130_fd_sc_hd__o211a_1 _12046_ (.A1(\core.pipe0_currentInstruction[10] ),
    .A2(net584),
    .B1(_06867_),
    .C1(net1821),
    .X(_00042_));
 sky130_fd_sc_hd__or2_1 _12047_ (.A(\core.csr.currentInstruction[11] ),
    .B(net588),
    .X(_06868_));
 sky130_fd_sc_hd__o211a_1 _12048_ (.A1(\core.pipe0_currentInstruction[11] ),
    .A2(net584),
    .B1(_06868_),
    .C1(net1821),
    .X(_00043_));
 sky130_fd_sc_hd__or2_1 _12049_ (.A(\core.csr.currentInstruction[12] ),
    .B(net591),
    .X(_06869_));
 sky130_fd_sc_hd__o211a_1 _12050_ (.A1(\core.pipe0_currentInstruction[12] ),
    .A2(net584),
    .B1(_06869_),
    .C1(net1822),
    .X(_00044_));
 sky130_fd_sc_hd__or2_1 _12051_ (.A(net1800),
    .B(net588),
    .X(_06870_));
 sky130_fd_sc_hd__o211a_1 _12052_ (.A1(\core.pipe0_currentInstruction[13] ),
    .A2(net584),
    .B1(_06870_),
    .C1(net1822),
    .X(_00045_));
 sky130_fd_sc_hd__or2_1 _12053_ (.A(net1799),
    .B(net591),
    .X(_06871_));
 sky130_fd_sc_hd__o211a_1 _12054_ (.A1(\core.pipe0_currentInstruction[14] ),
    .A2(net585),
    .B1(_06871_),
    .C1(net1835),
    .X(_00046_));
 sky130_fd_sc_hd__or2_1 _12055_ (.A(\core.csr.currentInstruction[15] ),
    .B(net589),
    .X(_06872_));
 sky130_fd_sc_hd__o211a_1 _12056_ (.A1(net1793),
    .A2(net586),
    .B1(_06872_),
    .C1(net1823),
    .X(_00047_));
 sky130_fd_sc_hd__or2_1 _12057_ (.A(\core.csr.currentInstruction[16] ),
    .B(net589),
    .X(_06873_));
 sky130_fd_sc_hd__o211a_1 _12058_ (.A1(net1792),
    .A2(net586),
    .B1(_06873_),
    .C1(net1823),
    .X(_00048_));
 sky130_fd_sc_hd__or2_1 _12059_ (.A(\core.csr.currentInstruction[17] ),
    .B(net591),
    .X(_06874_));
 sky130_fd_sc_hd__o211a_1 _12060_ (.A1(net1784),
    .A2(net586),
    .B1(_06874_),
    .C1(net1823),
    .X(_00049_));
 sky130_fd_sc_hd__or2_1 _12061_ (.A(\core.csr.currentInstruction[18] ),
    .B(net589),
    .X(_06875_));
 sky130_fd_sc_hd__o211a_1 _12062_ (.A1(\core.pipe0_currentInstruction[18] ),
    .A2(net586),
    .B1(_06875_),
    .C1(net1823),
    .X(_00050_));
 sky130_fd_sc_hd__or2_1 _12063_ (.A(\core.csr.currentInstruction[19] ),
    .B(net589),
    .X(_06876_));
 sky130_fd_sc_hd__o211a_1 _12064_ (.A1(net1783),
    .A2(net586),
    .B1(_06876_),
    .C1(net1824),
    .X(_00051_));
 sky130_fd_sc_hd__or2_1 _12065_ (.A(\core.csr.currentInstruction[20] ),
    .B(net589),
    .X(_06877_));
 sky130_fd_sc_hd__o211a_1 _12066_ (.A1(net1777),
    .A2(net587),
    .B1(_06877_),
    .C1(net1844),
    .X(_00052_));
 sky130_fd_sc_hd__or2_1 _12067_ (.A(\core.csr.currentInstruction[21] ),
    .B(net590),
    .X(_06878_));
 sky130_fd_sc_hd__o211a_1 _12068_ (.A1(net1775),
    .A2(net587),
    .B1(_06878_),
    .C1(net1844),
    .X(_00053_));
 sky130_fd_sc_hd__or2_1 _12069_ (.A(\core.csr.currentInstruction[22] ),
    .B(net590),
    .X(_06879_));
 sky130_fd_sc_hd__o211a_1 _12070_ (.A1(net1767),
    .A2(net587),
    .B1(_06879_),
    .C1(net1829),
    .X(_00054_));
 sky130_fd_sc_hd__or2_1 _12071_ (.A(\core.csr.currentInstruction[23] ),
    .B(net589),
    .X(_06880_));
 sky130_fd_sc_hd__o211a_1 _12072_ (.A1(net1762),
    .A2(net586),
    .B1(_06880_),
    .C1(net1829),
    .X(_00055_));
 sky130_fd_sc_hd__or2_1 _12073_ (.A(\core.csr.currentInstruction[24] ),
    .B(net591),
    .X(_06881_));
 sky130_fd_sc_hd__o211a_1 _12074_ (.A1(net1755),
    .A2(net586),
    .B1(_06881_),
    .C1(net1823),
    .X(_00056_));
 sky130_fd_sc_hd__or2_1 _12075_ (.A(\core.csr.currentInstruction[25] ),
    .B(net589),
    .X(_06882_));
 sky130_fd_sc_hd__o211a_1 _12076_ (.A1(\core.pipe0_currentInstruction[25] ),
    .A2(net586),
    .B1(_06882_),
    .C1(net1829),
    .X(_00057_));
 sky130_fd_sc_hd__or2_1 _12077_ (.A(\core.csr.currentInstruction[26] ),
    .B(net589),
    .X(_06883_));
 sky130_fd_sc_hd__o211a_1 _12078_ (.A1(\core.pipe0_currentInstruction[26] ),
    .A2(net586),
    .B1(_06883_),
    .C1(net1829),
    .X(_00058_));
 sky130_fd_sc_hd__or2_1 _12079_ (.A(\core.csr.currentInstruction[27] ),
    .B(net589),
    .X(_06884_));
 sky130_fd_sc_hd__o211a_1 _12080_ (.A1(\core.pipe0_currentInstruction[27] ),
    .A2(net587),
    .B1(_06884_),
    .C1(net1829),
    .X(_00059_));
 sky130_fd_sc_hd__or2_1 _12081_ (.A(\core.csr.currentInstruction[28] ),
    .B(net590),
    .X(_06885_));
 sky130_fd_sc_hd__o211a_1 _12082_ (.A1(\core.pipe0_currentInstruction[28] ),
    .A2(net587),
    .B1(_06885_),
    .C1(net1844),
    .X(_00060_));
 sky130_fd_sc_hd__or2_1 _12083_ (.A(\core.csr.currentInstruction[29] ),
    .B(net590),
    .X(_06886_));
 sky130_fd_sc_hd__o211a_1 _12084_ (.A1(\core.pipe0_currentInstruction[29] ),
    .A2(net587),
    .B1(_06886_),
    .C1(net1844),
    .X(_00061_));
 sky130_fd_sc_hd__or2_1 _12085_ (.A(\core.csr.currentInstruction[30] ),
    .B(net589),
    .X(_06887_));
 sky130_fd_sc_hd__o211a_1 _12086_ (.A1(net1752),
    .A2(net586),
    .B1(_06887_),
    .C1(net1829),
    .X(_00062_));
 sky130_fd_sc_hd__or2_1 _12087_ (.A(\core.csr.currentInstruction[31] ),
    .B(net590),
    .X(_06888_));
 sky130_fd_sc_hd__o211a_1 _12088_ (.A1(\core.pipe0_currentInstruction[31] ),
    .A2(net587),
    .B1(_06888_),
    .C1(net1844),
    .X(_00063_));
 sky130_fd_sc_hd__nand2_1 _12089_ (.A(_03808_),
    .B(net596),
    .Y(_06889_));
 sky130_fd_sc_hd__a21o_1 _12090_ (.A1(net585),
    .A2(_06889_),
    .B1(net1906),
    .X(_00064_));
 sky130_fd_sc_hd__nor2_1 _12091_ (.A(net1889),
    .B(\core.csr.cycleTimer.currentValue[0] ),
    .Y(_00065_));
 sky130_fd_sc_hd__a21oi_1 _12092_ (.A1(\core.csr.cycleTimer.currentValue[0] ),
    .A2(\core.csr.cycleTimer.currentValue[1] ),
    .B1(net1889),
    .Y(_06890_));
 sky130_fd_sc_hd__o21a_1 _12093_ (.A1(\core.csr.cycleTimer.currentValue[0] ),
    .A2(\core.csr.cycleTimer.currentValue[1] ),
    .B1(_06890_),
    .X(_00066_));
 sky130_fd_sc_hd__a21oi_1 _12094_ (.A1(\core.csr.cycleTimer.currentValue[0] ),
    .A2(\core.csr.cycleTimer.currentValue[1] ),
    .B1(\core.csr.cycleTimer.currentValue[2] ),
    .Y(_06891_));
 sky130_fd_sc_hd__and3_2 _12095_ (.A(\core.csr.cycleTimer.currentValue[0] ),
    .B(\core.csr.cycleTimer.currentValue[1] ),
    .C(\core.csr.cycleTimer.currentValue[2] ),
    .X(_06892_));
 sky130_fd_sc_hd__nor3_1 _12096_ (.A(net1889),
    .B(_06891_),
    .C(_06892_),
    .Y(_00067_));
 sky130_fd_sc_hd__and2_1 _12097_ (.A(\core.csr.cycleTimer.currentValue[3] ),
    .B(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__nor2_1 _12098_ (.A(net1889),
    .B(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__o21a_1 _12099_ (.A1(\core.csr.cycleTimer.currentValue[3] ),
    .A2(_06892_),
    .B1(_06894_),
    .X(_00068_));
 sky130_fd_sc_hd__and3_2 _12100_ (.A(\core.csr.cycleTimer.currentValue[3] ),
    .B(\core.csr.cycleTimer.currentValue[4] ),
    .C(_06892_),
    .X(_06895_));
 sky130_fd_sc_hd__nor2_1 _12101_ (.A(net1889),
    .B(_06895_),
    .Y(_06896_));
 sky130_fd_sc_hd__o21a_1 _12102_ (.A1(\core.csr.cycleTimer.currentValue[4] ),
    .A2(_06893_),
    .B1(_06896_),
    .X(_00069_));
 sky130_fd_sc_hd__and2_1 _12103_ (.A(\core.csr.cycleTimer.currentValue[5] ),
    .B(_06895_),
    .X(_06897_));
 sky130_fd_sc_hd__nor2_1 _12104_ (.A(net1889),
    .B(_06897_),
    .Y(_06898_));
 sky130_fd_sc_hd__o21a_1 _12105_ (.A1(\core.csr.cycleTimer.currentValue[5] ),
    .A2(_06895_),
    .B1(_06898_),
    .X(_00070_));
 sky130_fd_sc_hd__and3_2 _12106_ (.A(\core.csr.cycleTimer.currentValue[5] ),
    .B(\core.csr.cycleTimer.currentValue[6] ),
    .C(_06895_),
    .X(_06899_));
 sky130_fd_sc_hd__nor2_1 _12107_ (.A(net1889),
    .B(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__o21a_1 _12108_ (.A1(\core.csr.cycleTimer.currentValue[6] ),
    .A2(_06897_),
    .B1(_06900_),
    .X(_00071_));
 sky130_fd_sc_hd__a21oi_1 _12109_ (.A1(\core.csr.cycleTimer.currentValue[7] ),
    .A2(_06899_),
    .B1(net1887),
    .Y(_06901_));
 sky130_fd_sc_hd__o21a_1 _12110_ (.A1(\core.csr.cycleTimer.currentValue[7] ),
    .A2(_06899_),
    .B1(_06901_),
    .X(_00072_));
 sky130_fd_sc_hd__a21oi_1 _12111_ (.A1(\core.csr.cycleTimer.currentValue[7] ),
    .A2(_06899_),
    .B1(\core.csr.cycleTimer.currentValue[8] ),
    .Y(_06902_));
 sky130_fd_sc_hd__and3_1 _12112_ (.A(\core.csr.cycleTimer.currentValue[7] ),
    .B(\core.csr.cycleTimer.currentValue[8] ),
    .C(_06899_),
    .X(_06903_));
 sky130_fd_sc_hd__nor3_1 _12113_ (.A(net1892),
    .B(_06902_),
    .C(_06903_),
    .Y(_00073_));
 sky130_fd_sc_hd__and2_2 _12114_ (.A(\core.csr.cycleTimer.currentValue[9] ),
    .B(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__nor2_1 _12115_ (.A(net1892),
    .B(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__o21a_1 _12116_ (.A1(\core.csr.cycleTimer.currentValue[9] ),
    .A2(_06903_),
    .B1(_06905_),
    .X(_00074_));
 sky130_fd_sc_hd__a21oi_1 _12117_ (.A1(\core.csr.cycleTimer.currentValue[10] ),
    .A2(_06904_),
    .B1(net1893),
    .Y(_06906_));
 sky130_fd_sc_hd__o21a_1 _12118_ (.A1(\core.csr.cycleTimer.currentValue[10] ),
    .A2(_06904_),
    .B1(_06906_),
    .X(_00075_));
 sky130_fd_sc_hd__a21oi_1 _12119_ (.A1(\core.csr.cycleTimer.currentValue[10] ),
    .A2(_06904_),
    .B1(\core.csr.cycleTimer.currentValue[11] ),
    .Y(_06907_));
 sky130_fd_sc_hd__and3_1 _12120_ (.A(\core.csr.cycleTimer.currentValue[10] ),
    .B(\core.csr.cycleTimer.currentValue[11] ),
    .C(_06904_),
    .X(_06908_));
 sky130_fd_sc_hd__nor3_1 _12121_ (.A(net1893),
    .B(_06907_),
    .C(_06908_),
    .Y(_00076_));
 sky130_fd_sc_hd__and2_2 _12122_ (.A(\core.csr.cycleTimer.currentValue[12] ),
    .B(_06908_),
    .X(_06909_));
 sky130_fd_sc_hd__nor2_1 _12123_ (.A(net1885),
    .B(_06909_),
    .Y(_06910_));
 sky130_fd_sc_hd__o21a_1 _12124_ (.A1(\core.csr.cycleTimer.currentValue[12] ),
    .A2(_06908_),
    .B1(_06910_),
    .X(_00077_));
 sky130_fd_sc_hd__a21oi_1 _12125_ (.A1(\core.csr.cycleTimer.currentValue[13] ),
    .A2(_06909_),
    .B1(net1885),
    .Y(_06911_));
 sky130_fd_sc_hd__o21a_1 _12126_ (.A1(\core.csr.cycleTimer.currentValue[13] ),
    .A2(_06909_),
    .B1(_06911_),
    .X(_00078_));
 sky130_fd_sc_hd__a21oi_1 _12127_ (.A1(\core.csr.cycleTimer.currentValue[13] ),
    .A2(_06909_),
    .B1(\core.csr.cycleTimer.currentValue[14] ),
    .Y(_06912_));
 sky130_fd_sc_hd__and3_1 _12128_ (.A(\core.csr.cycleTimer.currentValue[13] ),
    .B(\core.csr.cycleTimer.currentValue[14] ),
    .C(_06909_),
    .X(_06913_));
 sky130_fd_sc_hd__nor3_1 _12129_ (.A(net1885),
    .B(_06912_),
    .C(_06913_),
    .Y(_00079_));
 sky130_fd_sc_hd__and2_2 _12130_ (.A(\core.csr.cycleTimer.currentValue[15] ),
    .B(_06913_),
    .X(_06914_));
 sky130_fd_sc_hd__nor2_1 _12131_ (.A(net1885),
    .B(_06914_),
    .Y(_06915_));
 sky130_fd_sc_hd__o21a_1 _12132_ (.A1(\core.csr.cycleTimer.currentValue[15] ),
    .A2(_06913_),
    .B1(_06915_),
    .X(_00080_));
 sky130_fd_sc_hd__a21oi_1 _12133_ (.A1(\core.csr.cycleTimer.currentValue[16] ),
    .A2(_06914_),
    .B1(net1885),
    .Y(_06916_));
 sky130_fd_sc_hd__o21a_1 _12134_ (.A1(\core.csr.cycleTimer.currentValue[16] ),
    .A2(_06914_),
    .B1(_06916_),
    .X(_00081_));
 sky130_fd_sc_hd__a21oi_1 _12135_ (.A1(\core.csr.cycleTimer.currentValue[16] ),
    .A2(_06914_),
    .B1(\core.csr.cycleTimer.currentValue[17] ),
    .Y(_06917_));
 sky130_fd_sc_hd__and3_1 _12136_ (.A(\core.csr.cycleTimer.currentValue[16] ),
    .B(\core.csr.cycleTimer.currentValue[17] ),
    .C(_06914_),
    .X(_06918_));
 sky130_fd_sc_hd__nor3_1 _12137_ (.A(net1885),
    .B(_06917_),
    .C(_06918_),
    .Y(_00082_));
 sky130_fd_sc_hd__and2_2 _12138_ (.A(\core.csr.cycleTimer.currentValue[18] ),
    .B(_06918_),
    .X(_06919_));
 sky130_fd_sc_hd__nor2_1 _12139_ (.A(net1885),
    .B(_06919_),
    .Y(_06920_));
 sky130_fd_sc_hd__o21a_1 _12140_ (.A1(\core.csr.cycleTimer.currentValue[18] ),
    .A2(_06918_),
    .B1(_06920_),
    .X(_00083_));
 sky130_fd_sc_hd__a21oi_1 _12141_ (.A1(\core.csr.cycleTimer.currentValue[19] ),
    .A2(_06919_),
    .B1(net1881),
    .Y(_06921_));
 sky130_fd_sc_hd__o21a_1 _12142_ (.A1(\core.csr.cycleTimer.currentValue[19] ),
    .A2(_06919_),
    .B1(_06921_),
    .X(_00084_));
 sky130_fd_sc_hd__a21oi_1 _12143_ (.A1(\core.csr.cycleTimer.currentValue[19] ),
    .A2(_06919_),
    .B1(\core.csr.cycleTimer.currentValue[20] ),
    .Y(_06922_));
 sky130_fd_sc_hd__and3_1 _12144_ (.A(\core.csr.cycleTimer.currentValue[19] ),
    .B(\core.csr.cycleTimer.currentValue[20] ),
    .C(_06919_),
    .X(_06923_));
 sky130_fd_sc_hd__nor3_1 _12145_ (.A(net1881),
    .B(_06922_),
    .C(_06923_),
    .Y(_00085_));
 sky130_fd_sc_hd__and2_2 _12146_ (.A(\core.csr.cycleTimer.currentValue[21] ),
    .B(_06923_),
    .X(_06924_));
 sky130_fd_sc_hd__nor2_1 _12147_ (.A(net1880),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__o21a_1 _12148_ (.A1(\core.csr.cycleTimer.currentValue[21] ),
    .A2(_06923_),
    .B1(_06925_),
    .X(_00086_));
 sky130_fd_sc_hd__a21oi_1 _12149_ (.A1(\core.csr.cycleTimer.currentValue[22] ),
    .A2(_06924_),
    .B1(net1880),
    .Y(_06926_));
 sky130_fd_sc_hd__o21a_1 _12150_ (.A1(\core.csr.cycleTimer.currentValue[22] ),
    .A2(_06924_),
    .B1(_06926_),
    .X(_00087_));
 sky130_fd_sc_hd__a21oi_1 _12151_ (.A1(\core.csr.cycleTimer.currentValue[22] ),
    .A2(_06924_),
    .B1(\core.csr.cycleTimer.currentValue[23] ),
    .Y(_06927_));
 sky130_fd_sc_hd__and3_2 _12152_ (.A(\core.csr.cycleTimer.currentValue[22] ),
    .B(\core.csr.cycleTimer.currentValue[23] ),
    .C(_06924_),
    .X(_06928_));
 sky130_fd_sc_hd__nor3_1 _12153_ (.A(net1880),
    .B(_06927_),
    .C(_06928_),
    .Y(_00088_));
 sky130_fd_sc_hd__and2_2 _12154_ (.A(\core.csr.cycleTimer.currentValue[24] ),
    .B(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__nor2_1 _12155_ (.A(net1882),
    .B(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__o21a_1 _12156_ (.A1(\core.csr.cycleTimer.currentValue[24] ),
    .A2(_06928_),
    .B1(_06930_),
    .X(_00089_));
 sky130_fd_sc_hd__a21oi_1 _12157_ (.A1(\core.csr.cycleTimer.currentValue[25] ),
    .A2(_06929_),
    .B1(net1883),
    .Y(_06931_));
 sky130_fd_sc_hd__o21a_1 _12158_ (.A1(\core.csr.cycleTimer.currentValue[25] ),
    .A2(_06929_),
    .B1(_06931_),
    .X(_00090_));
 sky130_fd_sc_hd__a21oi_1 _12159_ (.A1(\core.csr.cycleTimer.currentValue[25] ),
    .A2(_06929_),
    .B1(\core.csr.cycleTimer.currentValue[26] ),
    .Y(_06932_));
 sky130_fd_sc_hd__and3_1 _12160_ (.A(\core.csr.cycleTimer.currentValue[25] ),
    .B(\core.csr.cycleTimer.currentValue[26] ),
    .C(_06929_),
    .X(_06933_));
 sky130_fd_sc_hd__nor3_1 _12161_ (.A(net1883),
    .B(_06932_),
    .C(_06933_),
    .Y(_00091_));
 sky130_fd_sc_hd__and2_2 _12162_ (.A(\core.csr.cycleTimer.currentValue[27] ),
    .B(_06933_),
    .X(_06934_));
 sky130_fd_sc_hd__nor2_1 _12163_ (.A(net1883),
    .B(_06934_),
    .Y(_06935_));
 sky130_fd_sc_hd__o21a_1 _12164_ (.A1(\core.csr.cycleTimer.currentValue[27] ),
    .A2(_06933_),
    .B1(_06935_),
    .X(_00092_));
 sky130_fd_sc_hd__a21oi_1 _12165_ (.A1(\core.csr.cycleTimer.currentValue[28] ),
    .A2(_06934_),
    .B1(net1894),
    .Y(_06936_));
 sky130_fd_sc_hd__o21a_1 _12166_ (.A1(\core.csr.cycleTimer.currentValue[28] ),
    .A2(_06934_),
    .B1(_06936_),
    .X(_00093_));
 sky130_fd_sc_hd__a21oi_1 _12167_ (.A1(\core.csr.cycleTimer.currentValue[28] ),
    .A2(_06934_),
    .B1(\core.csr.cycleTimer.currentValue[29] ),
    .Y(_06937_));
 sky130_fd_sc_hd__and3_1 _12168_ (.A(\core.csr.cycleTimer.currentValue[28] ),
    .B(\core.csr.cycleTimer.currentValue[29] ),
    .C(_06934_),
    .X(_06938_));
 sky130_fd_sc_hd__nor3_1 _12169_ (.A(net1893),
    .B(_06937_),
    .C(_06938_),
    .Y(_00094_));
 sky130_fd_sc_hd__and2_2 _12170_ (.A(\core.csr.cycleTimer.currentValue[30] ),
    .B(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__nor2_1 _12171_ (.A(net1893),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__o21a_1 _12172_ (.A1(\core.csr.cycleTimer.currentValue[30] ),
    .A2(_06938_),
    .B1(_06940_),
    .X(_00095_));
 sky130_fd_sc_hd__a21oi_1 _12173_ (.A1(\core.csr.cycleTimer.currentValue[31] ),
    .A2(_06939_),
    .B1(net1892),
    .Y(_06941_));
 sky130_fd_sc_hd__o21a_1 _12174_ (.A1(\core.csr.cycleTimer.currentValue[31] ),
    .A2(_06939_),
    .B1(_06941_),
    .X(_00096_));
 sky130_fd_sc_hd__a21oi_1 _12175_ (.A1(\core.csr.cycleTimer.currentValue[31] ),
    .A2(_06939_),
    .B1(\core.csr.cycleTimer.currentValue[32] ),
    .Y(_06942_));
 sky130_fd_sc_hd__and3_1 _12176_ (.A(\core.csr.cycleTimer.currentValue[32] ),
    .B(\core.csr.cycleTimer.currentValue[31] ),
    .C(_06939_),
    .X(_06943_));
 sky130_fd_sc_hd__nor3_1 _12177_ (.A(net1892),
    .B(_06942_),
    .C(_06943_),
    .Y(_00097_));
 sky130_fd_sc_hd__and2_2 _12178_ (.A(\core.csr.cycleTimer.currentValue[33] ),
    .B(_06943_),
    .X(_06944_));
 sky130_fd_sc_hd__nor2_1 _12179_ (.A(net1890),
    .B(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__o21a_1 _12180_ (.A1(\core.csr.cycleTimer.currentValue[33] ),
    .A2(_06943_),
    .B1(_06945_),
    .X(_00098_));
 sky130_fd_sc_hd__a21oi_1 _12181_ (.A1(\core.csr.cycleTimer.currentValue[34] ),
    .A2(_06944_),
    .B1(net1890),
    .Y(_06946_));
 sky130_fd_sc_hd__o21a_1 _12182_ (.A1(\core.csr.cycleTimer.currentValue[34] ),
    .A2(_06944_),
    .B1(_06946_),
    .X(_00099_));
 sky130_fd_sc_hd__a21oi_1 _12183_ (.A1(\core.csr.cycleTimer.currentValue[34] ),
    .A2(_06944_),
    .B1(\core.csr.cycleTimer.currentValue[35] ),
    .Y(_06947_));
 sky130_fd_sc_hd__and3_1 _12184_ (.A(\core.csr.cycleTimer.currentValue[34] ),
    .B(\core.csr.cycleTimer.currentValue[35] ),
    .C(_06944_),
    .X(_06948_));
 sky130_fd_sc_hd__nor3_1 _12185_ (.A(net1890),
    .B(_06947_),
    .C(_06948_),
    .Y(_00100_));
 sky130_fd_sc_hd__and2_2 _12186_ (.A(\core.csr.cycleTimer.currentValue[36] ),
    .B(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__nor2_1 _12187_ (.A(net1890),
    .B(_06949_),
    .Y(_06950_));
 sky130_fd_sc_hd__o21a_1 _12188_ (.A1(\core.csr.cycleTimer.currentValue[36] ),
    .A2(_06948_),
    .B1(_06950_),
    .X(_00101_));
 sky130_fd_sc_hd__a21oi_1 _12189_ (.A1(\core.csr.cycleTimer.currentValue[37] ),
    .A2(_06949_),
    .B1(net1899),
    .Y(_06951_));
 sky130_fd_sc_hd__o21a_1 _12190_ (.A1(\core.csr.cycleTimer.currentValue[37] ),
    .A2(_06949_),
    .B1(_06951_),
    .X(_00102_));
 sky130_fd_sc_hd__a21oi_1 _12191_ (.A1(\core.csr.cycleTimer.currentValue[37] ),
    .A2(_06949_),
    .B1(\core.csr.cycleTimer.currentValue[38] ),
    .Y(_06952_));
 sky130_fd_sc_hd__and3_1 _12192_ (.A(\core.csr.cycleTimer.currentValue[37] ),
    .B(\core.csr.cycleTimer.currentValue[38] ),
    .C(_06949_),
    .X(_06953_));
 sky130_fd_sc_hd__nor3_1 _12193_ (.A(net1898),
    .B(_06952_),
    .C(_06953_),
    .Y(_00103_));
 sky130_fd_sc_hd__and2_2 _12194_ (.A(\core.csr.cycleTimer.currentValue[39] ),
    .B(_06953_),
    .X(_06954_));
 sky130_fd_sc_hd__nor2_1 _12195_ (.A(net1898),
    .B(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__o21a_1 _12196_ (.A1(\core.csr.cycleTimer.currentValue[39] ),
    .A2(_06953_),
    .B1(_06955_),
    .X(_00104_));
 sky130_fd_sc_hd__a21oi_1 _12197_ (.A1(\core.csr.cycleTimer.currentValue[40] ),
    .A2(_06954_),
    .B1(net1892),
    .Y(_06956_));
 sky130_fd_sc_hd__o21a_1 _12198_ (.A1(\core.csr.cycleTimer.currentValue[40] ),
    .A2(_06954_),
    .B1(_06956_),
    .X(_00105_));
 sky130_fd_sc_hd__a21oi_1 _12199_ (.A1(\core.csr.cycleTimer.currentValue[40] ),
    .A2(_06954_),
    .B1(\core.csr.cycleTimer.currentValue[41] ),
    .Y(_06957_));
 sky130_fd_sc_hd__and3_1 _12200_ (.A(\core.csr.cycleTimer.currentValue[40] ),
    .B(\core.csr.cycleTimer.currentValue[41] ),
    .C(_06954_),
    .X(_06958_));
 sky130_fd_sc_hd__nor3_1 _12201_ (.A(net1892),
    .B(_06957_),
    .C(_06958_),
    .Y(_00106_));
 sky130_fd_sc_hd__and2_2 _12202_ (.A(\core.csr.cycleTimer.currentValue[42] ),
    .B(_06958_),
    .X(_06959_));
 sky130_fd_sc_hd__nor2_1 _12203_ (.A(net1892),
    .B(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__o21a_1 _12204_ (.A1(\core.csr.cycleTimer.currentValue[42] ),
    .A2(_06958_),
    .B1(_06960_),
    .X(_00107_));
 sky130_fd_sc_hd__a21oi_1 _12205_ (.A1(\core.csr.cycleTimer.currentValue[43] ),
    .A2(_06959_),
    .B1(net1893),
    .Y(_06961_));
 sky130_fd_sc_hd__o21a_1 _12206_ (.A1(\core.csr.cycleTimer.currentValue[43] ),
    .A2(_06959_),
    .B1(_06961_),
    .X(_00108_));
 sky130_fd_sc_hd__a21oi_1 _12207_ (.A1(\core.csr.cycleTimer.currentValue[43] ),
    .A2(_06959_),
    .B1(\core.csr.cycleTimer.currentValue[44] ),
    .Y(_06962_));
 sky130_fd_sc_hd__and3_1 _12208_ (.A(\core.csr.cycleTimer.currentValue[43] ),
    .B(\core.csr.cycleTimer.currentValue[44] ),
    .C(_06959_),
    .X(_06963_));
 sky130_fd_sc_hd__nor3_1 _12209_ (.A(net1893),
    .B(_06962_),
    .C(_06963_),
    .Y(_00109_));
 sky130_fd_sc_hd__and2_2 _12210_ (.A(\core.csr.cycleTimer.currentValue[45] ),
    .B(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__nor2_1 _12211_ (.A(net1893),
    .B(_06964_),
    .Y(_06965_));
 sky130_fd_sc_hd__o21a_1 _12212_ (.A1(\core.csr.cycleTimer.currentValue[45] ),
    .A2(_06963_),
    .B1(_06965_),
    .X(_00110_));
 sky130_fd_sc_hd__a21oi_1 _12213_ (.A1(\core.csr.cycleTimer.currentValue[46] ),
    .A2(_06964_),
    .B1(net1885),
    .Y(_06966_));
 sky130_fd_sc_hd__o21a_1 _12214_ (.A1(\core.csr.cycleTimer.currentValue[46] ),
    .A2(_06964_),
    .B1(_06966_),
    .X(_00111_));
 sky130_fd_sc_hd__a21oi_1 _12215_ (.A1(\core.csr.cycleTimer.currentValue[46] ),
    .A2(_06964_),
    .B1(\core.csr.cycleTimer.currentValue[47] ),
    .Y(_06967_));
 sky130_fd_sc_hd__and3_1 _12216_ (.A(\core.csr.cycleTimer.currentValue[46] ),
    .B(\core.csr.cycleTimer.currentValue[47] ),
    .C(_06964_),
    .X(_06968_));
 sky130_fd_sc_hd__nor3_1 _12217_ (.A(net1885),
    .B(_06967_),
    .C(_06968_),
    .Y(_00112_));
 sky130_fd_sc_hd__and2_2 _12218_ (.A(\core.csr.cycleTimer.currentValue[48] ),
    .B(_06968_),
    .X(_06969_));
 sky130_fd_sc_hd__nor2_1 _12219_ (.A(net1885),
    .B(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__o21a_1 _12220_ (.A1(\core.csr.cycleTimer.currentValue[48] ),
    .A2(_06968_),
    .B1(_06970_),
    .X(_00113_));
 sky130_fd_sc_hd__a21oi_1 _12221_ (.A1(\core.csr.cycleTimer.currentValue[49] ),
    .A2(_06969_),
    .B1(net1882),
    .Y(_06971_));
 sky130_fd_sc_hd__o21a_1 _12222_ (.A1(\core.csr.cycleTimer.currentValue[49] ),
    .A2(_06969_),
    .B1(_06971_),
    .X(_00114_));
 sky130_fd_sc_hd__a21oi_1 _12223_ (.A1(\core.csr.cycleTimer.currentValue[49] ),
    .A2(_06969_),
    .B1(\core.csr.cycleTimer.currentValue[50] ),
    .Y(_06972_));
 sky130_fd_sc_hd__and3_1 _12224_ (.A(\core.csr.cycleTimer.currentValue[49] ),
    .B(\core.csr.cycleTimer.currentValue[50] ),
    .C(_06969_),
    .X(_06973_));
 sky130_fd_sc_hd__nor3_1 _12225_ (.A(net1882),
    .B(_06972_),
    .C(_06973_),
    .Y(_00115_));
 sky130_fd_sc_hd__and2_2 _12226_ (.A(\core.csr.cycleTimer.currentValue[51] ),
    .B(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__nor2_1 _12227_ (.A(net1882),
    .B(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__o21a_1 _12228_ (.A1(\core.csr.cycleTimer.currentValue[51] ),
    .A2(_06973_),
    .B1(_06975_),
    .X(_00116_));
 sky130_fd_sc_hd__a21oi_1 _12229_ (.A1(\core.csr.cycleTimer.currentValue[52] ),
    .A2(_06974_),
    .B1(net1882),
    .Y(_06976_));
 sky130_fd_sc_hd__o21a_1 _12230_ (.A1(\core.csr.cycleTimer.currentValue[52] ),
    .A2(_06974_),
    .B1(_06976_),
    .X(_00117_));
 sky130_fd_sc_hd__a21oi_1 _12231_ (.A1(\core.csr.cycleTimer.currentValue[52] ),
    .A2(_06974_),
    .B1(\core.csr.cycleTimer.currentValue[53] ),
    .Y(_06977_));
 sky130_fd_sc_hd__and3_1 _12232_ (.A(\core.csr.cycleTimer.currentValue[52] ),
    .B(\core.csr.cycleTimer.currentValue[53] ),
    .C(_06974_),
    .X(_06978_));
 sky130_fd_sc_hd__nor3_1 _12233_ (.A(net1882),
    .B(_06977_),
    .C(_06978_),
    .Y(_00118_));
 sky130_fd_sc_hd__and2_2 _12234_ (.A(\core.csr.cycleTimer.currentValue[54] ),
    .B(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__nor2_1 _12235_ (.A(net1882),
    .B(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__o21a_1 _12236_ (.A1(\core.csr.cycleTimer.currentValue[54] ),
    .A2(_06978_),
    .B1(_06980_),
    .X(_00119_));
 sky130_fd_sc_hd__a21oi_1 _12237_ (.A1(\core.csr.cycleTimer.currentValue[55] ),
    .A2(_06979_),
    .B1(net1882),
    .Y(_06981_));
 sky130_fd_sc_hd__o21a_1 _12238_ (.A1(\core.csr.cycleTimer.currentValue[55] ),
    .A2(_06979_),
    .B1(_06981_),
    .X(_00120_));
 sky130_fd_sc_hd__a21oi_1 _12239_ (.A1(\core.csr.cycleTimer.currentValue[55] ),
    .A2(_06979_),
    .B1(\core.csr.cycleTimer.currentValue[56] ),
    .Y(_06982_));
 sky130_fd_sc_hd__and3_1 _12240_ (.A(\core.csr.cycleTimer.currentValue[55] ),
    .B(\core.csr.cycleTimer.currentValue[56] ),
    .C(_06979_),
    .X(_06983_));
 sky130_fd_sc_hd__nor3_1 _12241_ (.A(net1882),
    .B(_06982_),
    .C(_06983_),
    .Y(_00121_));
 sky130_fd_sc_hd__and2_2 _12242_ (.A(\core.csr.cycleTimer.currentValue[57] ),
    .B(_06983_),
    .X(_06984_));
 sky130_fd_sc_hd__nor2_1 _12243_ (.A(net1883),
    .B(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__o21a_1 _12244_ (.A1(\core.csr.cycleTimer.currentValue[57] ),
    .A2(_06983_),
    .B1(_06985_),
    .X(_00122_));
 sky130_fd_sc_hd__a21oi_1 _12245_ (.A1(\core.csr.cycleTimer.currentValue[58] ),
    .A2(_06984_),
    .B1(net1883),
    .Y(_06986_));
 sky130_fd_sc_hd__o21a_1 _12246_ (.A1(\core.csr.cycleTimer.currentValue[58] ),
    .A2(_06984_),
    .B1(_06986_),
    .X(_00123_));
 sky130_fd_sc_hd__a21oi_1 _12247_ (.A1(\core.csr.cycleTimer.currentValue[58] ),
    .A2(_06984_),
    .B1(\core.csr.cycleTimer.currentValue[59] ),
    .Y(_06987_));
 sky130_fd_sc_hd__and3_2 _12248_ (.A(\core.csr.cycleTimer.currentValue[58] ),
    .B(\core.csr.cycleTimer.currentValue[59] ),
    .C(_06984_),
    .X(_06988_));
 sky130_fd_sc_hd__nor3_1 _12249_ (.A(net1884),
    .B(_06987_),
    .C(_06988_),
    .Y(_00124_));
 sky130_fd_sc_hd__and2_1 _12250_ (.A(\core.csr.cycleTimer.currentValue[60] ),
    .B(_06988_),
    .X(_06989_));
 sky130_fd_sc_hd__nor2_1 _12251_ (.A(net1894),
    .B(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__o21a_1 _12252_ (.A1(\core.csr.cycleTimer.currentValue[60] ),
    .A2(_06988_),
    .B1(_06990_),
    .X(_00125_));
 sky130_fd_sc_hd__and3_1 _12253_ (.A(\core.csr.cycleTimer.currentValue[60] ),
    .B(\core.csr.cycleTimer.currentValue[61] ),
    .C(_06988_),
    .X(_06991_));
 sky130_fd_sc_hd__nor2_1 _12254_ (.A(net1894),
    .B(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__o21a_1 _12255_ (.A1(\core.csr.cycleTimer.currentValue[61] ),
    .A2(_06989_),
    .B1(_06992_),
    .X(_00126_));
 sky130_fd_sc_hd__and2_1 _12256_ (.A(\core.csr.cycleTimer.currentValue[62] ),
    .B(_06991_),
    .X(_06993_));
 sky130_fd_sc_hd__nor2_1 _12257_ (.A(net1893),
    .B(_06993_),
    .Y(_06994_));
 sky130_fd_sc_hd__o21a_1 _12258_ (.A1(\core.csr.cycleTimer.currentValue[62] ),
    .A2(_06991_),
    .B1(_06994_),
    .X(_00127_));
 sky130_fd_sc_hd__a21oi_1 _12259_ (.A1(\core.csr.cycleTimer.currentValue[63] ),
    .A2(_06993_),
    .B1(net1892),
    .Y(_06995_));
 sky130_fd_sc_hd__o21a_1 _12260_ (.A1(\core.csr.cycleTimer.currentValue[63] ),
    .A2(_06993_),
    .B1(_06995_),
    .X(_00128_));
 sky130_fd_sc_hd__nand2_2 _12261_ (.A(\core.pipe0_currentInstruction[6] ),
    .B(_04050_),
    .Y(_06996_));
 sky130_fd_sc_hd__or3b_4 _12262_ (.A(_03858_),
    .B(_06996_),
    .C_N(_04052_),
    .X(_06997_));
 sky130_fd_sc_hd__inv_2 _12263_ (.A(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__and3_2 _12264_ (.A(_04047_),
    .B(_04048_),
    .C(_04062_),
    .X(_06999_));
 sky130_fd_sc_hd__nand2_4 _12265_ (.A(_04062_),
    .B(_06644_),
    .Y(_07000_));
 sky130_fd_sc_hd__nand2_1 _12266_ (.A(\core.pipe0_currentInstruction[3] ),
    .B(\core.pipe0_currentInstruction[2] ),
    .Y(_07001_));
 sky130_fd_sc_hd__or2_4 _12267_ (.A(_03857_),
    .B(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__o31ai_2 _12268_ (.A1(_04066_),
    .A2(net1235),
    .A3(_07002_),
    .B1(_06997_),
    .Y(_07003_));
 sky130_fd_sc_hd__or4b_4 _12269_ (.A(net203),
    .B(net202),
    .C(net204),
    .D_N(net205),
    .X(_07004_));
 sky130_fd_sc_hd__nor2_2 _12270_ (.A(_06697_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__or2_1 _12271_ (.A(_06697_),
    .B(_07004_),
    .X(_07006_));
 sky130_fd_sc_hd__and3b_2 _12272_ (.A_N(\jtag.managementState[1] ),
    .B(_03816_),
    .C(\jtag.managementState[2] ),
    .X(_07007_));
 sky130_fd_sc_hd__or3b_4 _12273_ (.A(\jtag.managementState[1] ),
    .B(\jtag.managementState[0] ),
    .C_N(\jtag.managementState[2] ),
    .X(_07008_));
 sky130_fd_sc_hd__or2_4 _12274_ (.A(\jtag.managementState[2] ),
    .B(\jtag.managementState[1] ),
    .X(_07009_));
 sky130_fd_sc_hd__nor2_4 _12275_ (.A(_03816_),
    .B(net1610),
    .Y(_07010_));
 sky130_fd_sc_hd__or2_2 _12276_ (.A(net1305),
    .B(_07010_),
    .X(_07011_));
 sky130_fd_sc_hd__nor2_1 _12277_ (.A(_07006_),
    .B(net1273),
    .Y(_07012_));
 sky130_fd_sc_hd__a22oi_4 _12278_ (.A1(\jtag.managementAddress[10] ),
    .A2(net1272),
    .B1(net1231),
    .B2(\wbSRAMInterface.currentAddress[10] ),
    .Y(_07013_));
 sky130_fd_sc_hd__a22oi_4 _12279_ (.A1(\jtag.managementAddress[12] ),
    .A2(net1272),
    .B1(net1231),
    .B2(\wbSRAMInterface.currentAddress[12] ),
    .Y(_07014_));
 sky130_fd_sc_hd__a22oi_4 _12280_ (.A1(\jtag.managementAddress[11] ),
    .A2(net1272),
    .B1(net1232),
    .B2(\wbSRAMInterface.currentAddress[11] ),
    .Y(_07015_));
 sky130_fd_sc_hd__a22o_2 _12281_ (.A1(\jtag.managementAddress[13] ),
    .A2(net1272),
    .B1(net1231),
    .B2(\wbSRAMInterface.currentAddress[13] ),
    .X(_07016_));
 sky130_fd_sc_hd__a22o_1 _12282_ (.A1(\jtag.managementAddress[8] ),
    .A2(net1272),
    .B1(net1231),
    .B2(\wbSRAMInterface.currentAddress[8] ),
    .X(_07017_));
 sky130_fd_sc_hd__a22o_1 _12283_ (.A1(\jtag.managementAddress[9] ),
    .A2(net1272),
    .B1(net1231),
    .B2(\wbSRAMInterface.currentAddress[9] ),
    .X(_07018_));
 sky130_fd_sc_hd__and3_1 _12284_ (.A(_07013_),
    .B(_07014_),
    .C(_07015_),
    .X(_07019_));
 sky130_fd_sc_hd__or4b_4 _12285_ (.A(_07016_),
    .B(_07017_),
    .C(_07018_),
    .D_N(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__a22o_4 _12286_ (.A1(\jtag.managementAddress[14] ),
    .A2(net1272),
    .B1(net1231),
    .B2(\wbSRAMInterface.currentAddress[14] ),
    .X(_07021_));
 sky130_fd_sc_hd__a22o_1 _12287_ (.A1(\jtag.managementAddress[7] ),
    .A2(net1272),
    .B1(net1231),
    .B2(\wbSRAMInterface.currentAddress[7] ),
    .X(_07022_));
 sky130_fd_sc_hd__a22o_2 _12288_ (.A1(\jtag.managementAddress[15] ),
    .A2(net1272),
    .B1(net1231),
    .B2(\wbSRAMInterface.currentAddress[15] ),
    .X(_07023_));
 sky130_fd_sc_hd__a22o_4 _12289_ (.A1(\jtag.managementAddress[6] ),
    .A2(net1273),
    .B1(net1230),
    .B2(\wbSRAMInterface.currentAddress[6] ),
    .X(_07024_));
 sky130_fd_sc_hd__or2_2 _12290_ (.A(_07022_),
    .B(_07023_),
    .X(_07025_));
 sky130_fd_sc_hd__nor2_1 _12291_ (.A(_07024_),
    .B(_07025_),
    .Y(_07026_));
 sky130_fd_sc_hd__or3_2 _12292_ (.A(_07021_),
    .B(_07024_),
    .C(_07025_),
    .X(_07027_));
 sky130_fd_sc_hd__a22o_2 _12293_ (.A1(\jtag.managementAddress[5] ),
    .A2(net1273),
    .B1(net1230),
    .B2(\wbSRAMInterface.currentAddress[5] ),
    .X(_07028_));
 sky130_fd_sc_hd__a22o_2 _12294_ (.A1(\jtag.managementAddress[4] ),
    .A2(net1273),
    .B1(net1230),
    .B2(\wbSRAMInterface.currentAddress[4] ),
    .X(_07029_));
 sky130_fd_sc_hd__or2_1 _12295_ (.A(_07028_),
    .B(_07029_),
    .X(_07030_));
 sky130_fd_sc_hd__or2_2 _12296_ (.A(_07027_),
    .B(_07030_),
    .X(_07031_));
 sky130_fd_sc_hd__a22o_2 _12297_ (.A1(\jtag.managementAddress[3] ),
    .A2(net1273),
    .B1(net1232),
    .B2(\wbSRAMInterface.currentAddress[3] ),
    .X(_07032_));
 sky130_fd_sc_hd__a22o_4 _12298_ (.A1(\jtag.managementAddress[2] ),
    .A2(net1273),
    .B1(net1230),
    .B2(\wbSRAMInterface.currentAddress[2] ),
    .X(_07033_));
 sky130_fd_sc_hd__or3b_4 _12299_ (.A(\jtag.managementAddress[1] ),
    .B(\jtag.managementAddress[0] ),
    .C_N(net1273),
    .X(_07034_));
 sky130_fd_sc_hd__o31a_1 _12300_ (.A1(\wbSRAMInterface.currentAddress[0] ),
    .A2(\wbSRAMInterface.currentAddress[1] ),
    .A3(net1273),
    .B1(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__or3b_1 _12301_ (.A(_07033_),
    .B(_07035_),
    .C_N(_07032_),
    .X(_07036_));
 sky130_fd_sc_hd__o31a_4 _12302_ (.A1(_06703_),
    .A2(_07004_),
    .A3(_07010_),
    .B1(_07008_),
    .X(_07037_));
 sky130_fd_sc_hd__or3_4 _12303_ (.A(\jtag.managementAddress[19] ),
    .B(\jtag.managementAddress[18] ),
    .C(\jtag.managementAddress[17] ),
    .X(_07038_));
 sky130_fd_sc_hd__a22o_2 _12304_ (.A1(_06699_),
    .A2(net1231),
    .B1(_07038_),
    .B2(_07011_),
    .X(_07039_));
 sky130_fd_sc_hd__a22o_2 _12305_ (.A1(\jtag.managementAddress[16] ),
    .A2(net1272),
    .B1(net1231),
    .B2(\wbSRAMInterface.currentAddress[16] ),
    .X(_07040_));
 sky130_fd_sc_hd__or3b_4 _12306_ (.A(net1725),
    .B(_07039_),
    .C_N(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__inv_2 _12307_ (.A(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__or4_1 _12308_ (.A(_07020_),
    .B(_07036_),
    .C(_07037_),
    .D(_07041_),
    .X(_07043_));
 sky130_fd_sc_hd__and3b_1 _12309_ (.A_N(_07039_),
    .B(_07040_),
    .C(net1714),
    .X(_07044_));
 sky130_fd_sc_hd__o21ai_2 _12310_ (.A1(_07031_),
    .A2(_07043_),
    .B1(net1713),
    .Y(_07045_));
 sky130_fd_sc_hd__clkinv_2 _12311_ (.A(_07045_),
    .Y(_07046_));
 sky130_fd_sc_hd__or2_4 _12312_ (.A(_07003_),
    .B(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__nor2_4 _12313_ (.A(_06996_),
    .B(_07002_),
    .Y(_07048_));
 sky130_fd_sc_hd__or2_4 _12314_ (.A(_06996_),
    .B(_07002_),
    .X(_07049_));
 sky130_fd_sc_hd__or2_4 _12315_ (.A(_03877_),
    .B(_06996_),
    .X(_07050_));
 sky130_fd_sc_hd__nor2_4 _12316_ (.A(net1234),
    .B(_07050_),
    .Y(_07051_));
 sky130_fd_sc_hd__or2_1 _12317_ (.A(net1234),
    .B(_07050_),
    .X(_07052_));
 sky130_fd_sc_hd__nor2_2 _12318_ (.A(net1229),
    .B(net1185),
    .Y(_07053_));
 sky130_fd_sc_hd__nand2_1 _12319_ (.A(net1221),
    .B(net1179),
    .Y(_07054_));
 sky130_fd_sc_hd__or4b_1 _12320_ (.A(net1764),
    .B(net1780),
    .C(_03869_),
    .D_N(net1319),
    .X(_07055_));
 sky130_fd_sc_hd__or4bb_4 _12321_ (.A(\core.pipe0_currentInstruction[27] ),
    .B(_07055_),
    .C_N(\core.pipe0_currentInstruction[29] ),
    .D_N(\core.pipe0_currentInstruction[28] ),
    .X(_07056_));
 sky130_fd_sc_hd__nor2_8 _12322_ (.A(_03867_),
    .B(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__or2_4 _12323_ (.A(_03867_),
    .B(_07056_),
    .X(_07058_));
 sky130_fd_sc_hd__o2111ai_1 _12324_ (.A1(net1796),
    .A2(_03900_),
    .B1(_03915_),
    .C1(\core.csr.currentInstruction[3] ),
    .D1(_03899_),
    .Y(_07059_));
 sky130_fd_sc_hd__a21o_1 _12325_ (.A1(_03931_),
    .A2(_07059_),
    .B1(_03928_),
    .X(_07060_));
 sky130_fd_sc_hd__or4_4 _12326_ (.A(\core.csr.currentInstruction[10] ),
    .B(net1801),
    .C(\core.csr.currentInstruction[8] ),
    .D(\core.csr.currentInstruction[7] ),
    .X(_07061_));
 sky130_fd_sc_hd__or4b_1 _12327_ (.A(\core.csr.currentInstruction[20] ),
    .B(\core.csr.currentInstruction[19] ),
    .C(\core.csr.currentInstruction[18] ),
    .D_N(\core.csr.currentInstruction[21] ),
    .X(_07062_));
 sky130_fd_sc_hd__or4_1 _12328_ (.A(\core.csr.currentInstruction[25] ),
    .B(\core.csr.currentInstruction[24] ),
    .C(\core.csr.currentInstruction[23] ),
    .D(\core.csr.currentInstruction[22] ),
    .X(_07063_));
 sky130_fd_sc_hd__or4bb_1 _12329_ (.A(\core.csr.currentInstruction[31] ),
    .B(\core.csr.currentInstruction[30] ),
    .C_N(\core.csr.currentInstruction[29] ),
    .D_N(\core.csr.currentInstruction[28] ),
    .X(_07064_));
 sky130_fd_sc_hd__or4_1 _12330_ (.A(\core.csr.currentInstruction[27] ),
    .B(\core.csr.currentInstruction[26] ),
    .C(_07062_),
    .D(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__or4_1 _12331_ (.A(\core.csr.currentInstruction[17] ),
    .B(\core.csr.currentInstruction[16] ),
    .C(\core.csr.currentInstruction[15] ),
    .D(\core.csr.currentInstruction[14] ),
    .X(_07066_));
 sky130_fd_sc_hd__or4_1 _12332_ (.A(\core.csr.currentInstruction[13] ),
    .B(\core.csr.currentInstruction[12] ),
    .C(\core.csr.currentInstruction[11] ),
    .D(_07066_),
    .X(_07067_));
 sky130_fd_sc_hd__or4_4 _12333_ (.A(_07061_),
    .B(_07063_),
    .C(_07065_),
    .D(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__o21ai_1 _12334_ (.A1(_03917_),
    .A2(_07068_),
    .B1(_07060_),
    .Y(_07069_));
 sky130_fd_sc_hd__a41o_2 _12335_ (.A1(\core.csr.currentInstruction[6] ),
    .A2(_03893_),
    .A3(_03898_),
    .A4(_03930_),
    .B1(_07069_),
    .X(_07070_));
 sky130_fd_sc_hd__o41a_1 _12336_ (.A1(_07047_),
    .A2(net1133),
    .A3(net1131),
    .A4(_07070_),
    .B1(net602),
    .X(_07071_));
 sky130_fd_sc_hd__a211o_1 _12337_ (.A1(\core.pipe0_fetch.currentPipeStall ),
    .A2(net596),
    .B1(_07071_),
    .C1(net1879),
    .X(_00129_));
 sky130_fd_sc_hd__nor2_4 _12338_ (.A(\core.pipe0_fetch.currentPipeStall ),
    .B(net596),
    .Y(_07072_));
 sky130_fd_sc_hd__a2bb2o_2 _12339_ (.A1_N(\coreWBInterface.readDataBuffered[0] ),
    .A2_N(net1315),
    .B1(_04979_),
    .B2(net1746),
    .X(_07073_));
 sky130_fd_sc_hd__nand2_1 _12340_ (.A(net576),
    .B(_07073_),
    .Y(_07074_));
 sky130_fd_sc_hd__o211a_1 _12341_ (.A1(\core.pipe0_currentInstruction[0] ),
    .A2(net576),
    .B1(_07074_),
    .C1(net1834),
    .X(_00130_));
 sky130_fd_sc_hd__a2bb2o_1 _12342_ (.A1_N(\coreWBInterface.readDataBuffered[1] ),
    .A2_N(net1315),
    .B1(_04895_),
    .B2(net1746),
    .X(_07075_));
 sky130_fd_sc_hd__nand2_1 _12343_ (.A(net577),
    .B(_07075_),
    .Y(_07076_));
 sky130_fd_sc_hd__o211a_1 _12344_ (.A1(\core.pipe0_currentInstruction[1] ),
    .A2(net576),
    .B1(_07076_),
    .C1(net1835),
    .X(_00131_));
 sky130_fd_sc_hd__o32ai_4 _12345_ (.A1(net1635),
    .A2(net1619),
    .A3(_04810_),
    .B1(net1315),
    .B2(\coreWBInterface.readDataBuffered[2] ),
    .Y(_07077_));
 sky130_fd_sc_hd__nand2_1 _12346_ (.A(net577),
    .B(_07077_),
    .Y(_07078_));
 sky130_fd_sc_hd__o211a_1 _12347_ (.A1(\core.pipe0_currentInstruction[2] ),
    .A2(net577),
    .B1(_07078_),
    .C1(net1835),
    .X(_00132_));
 sky130_fd_sc_hd__o32ai_4 _12348_ (.A1(net1637),
    .A2(net1620),
    .A3(_04726_),
    .B1(net1318),
    .B2(\coreWBInterface.readDataBuffered[3] ),
    .Y(_07079_));
 sky130_fd_sc_hd__nand2_1 _12349_ (.A(net577),
    .B(_07079_),
    .Y(_07080_));
 sky130_fd_sc_hd__o211a_1 _12350_ (.A1(\core.pipe0_currentInstruction[3] ),
    .A2(net576),
    .B1(_07080_),
    .C1(net1835),
    .X(_00133_));
 sky130_fd_sc_hd__o32ai_4 _12351_ (.A1(net1635),
    .A2(net1619),
    .A3(_04637_),
    .B1(net1315),
    .B2(\coreWBInterface.readDataBuffered[4] ),
    .Y(_07081_));
 sky130_fd_sc_hd__nand2_1 _12352_ (.A(net578),
    .B(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__o211a_1 _12353_ (.A1(\core.pipe0_currentInstruction[4] ),
    .A2(net577),
    .B1(_07082_),
    .C1(net1834),
    .X(_00134_));
 sky130_fd_sc_hd__o32ai_2 _12354_ (.A1(net1635),
    .A2(net1619),
    .A3(_04551_),
    .B1(net1315),
    .B2(\coreWBInterface.readDataBuffered[5] ),
    .Y(_07083_));
 sky130_fd_sc_hd__nand2_1 _12355_ (.A(net578),
    .B(_07083_),
    .Y(_07084_));
 sky130_fd_sc_hd__o211a_1 _12356_ (.A1(\core.pipe0_currentInstruction[5] ),
    .A2(net578),
    .B1(_07084_),
    .C1(net1836),
    .X(_00135_));
 sky130_fd_sc_hd__o32ai_4 _12357_ (.A1(net1635),
    .A2(net1619),
    .A3(_04465_),
    .B1(net1315),
    .B2(\coreWBInterface.readDataBuffered[6] ),
    .Y(_07085_));
 sky130_fd_sc_hd__nand2_1 _12358_ (.A(net580),
    .B(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__o211a_1 _12359_ (.A1(\core.pipe0_currentInstruction[6] ),
    .A2(net580),
    .B1(_07086_),
    .C1(net1837),
    .X(_00136_));
 sky130_fd_sc_hd__or2_1 _12360_ (.A(\core.pipe0_currentInstruction[7] ),
    .B(net576),
    .X(_07087_));
 sky130_fd_sc_hd__o32a_1 _12361_ (.A1(net1637),
    .A2(net1619),
    .A3(_03999_),
    .B1(net1318),
    .B2(\coreWBInterface.readDataBuffered[7] ),
    .X(_07088_));
 sky130_fd_sc_hd__o311a_1 _12362_ (.A1(\core.pipe0_fetch.currentPipeStall ),
    .A2(net597),
    .A3(_07088_),
    .B1(_07087_),
    .C1(net1834),
    .X(_00137_));
 sky130_fd_sc_hd__o32ai_4 _12363_ (.A1(net1636),
    .A2(_03989_),
    .A3(_04317_),
    .B1(net1317),
    .B2(\coreWBInterface.readDataBuffered[8] ),
    .Y(_07089_));
 sky130_fd_sc_hd__nand2_1 _12364_ (.A(net579),
    .B(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__o211a_1 _12365_ (.A1(\core.pipe0_currentInstruction[8] ),
    .A2(net580),
    .B1(_07090_),
    .C1(net1836),
    .X(_00138_));
 sky130_fd_sc_hd__a2bb2o_2 _12366_ (.A1_N(\coreWBInterface.readDataBuffered[9] ),
    .A2_N(net1317),
    .B1(_04231_),
    .B2(net1746),
    .X(_07091_));
 sky130_fd_sc_hd__nand2_1 _12367_ (.A(net579),
    .B(_07091_),
    .Y(_07092_));
 sky130_fd_sc_hd__o211a_1 _12368_ (.A1(\core.pipe0_currentInstruction[9] ),
    .A2(net579),
    .B1(_07092_),
    .C1(net1836),
    .X(_00139_));
 sky130_fd_sc_hd__a2bb2o_2 _12369_ (.A1_N(\coreWBInterface.readDataBuffered[10] ),
    .A2_N(net1317),
    .B1(_04142_),
    .B2(net1746),
    .X(_07093_));
 sky130_fd_sc_hd__nand2_1 _12370_ (.A(net576),
    .B(_07093_),
    .Y(_07094_));
 sky130_fd_sc_hd__o211a_1 _12371_ (.A1(\core.pipe0_currentInstruction[10] ),
    .A2(net576),
    .B1(_07094_),
    .C1(net1834),
    .X(_00140_));
 sky130_fd_sc_hd__a2bb2o_1 _12372_ (.A1_N(\coreWBInterface.readDataBuffered[11] ),
    .A2_N(net1318),
    .B1(_04033_),
    .B2(\memoryController.last_instruction_enableLocalMemory ),
    .X(_07095_));
 sky130_fd_sc_hd__nand2_1 _12373_ (.A(net583),
    .B(_07095_),
    .Y(_07096_));
 sky130_fd_sc_hd__o211a_1 _12374_ (.A1(\core.pipe0_currentInstruction[11] ),
    .A2(net580),
    .B1(_07096_),
    .C1(net1843),
    .X(_00141_));
 sky130_fd_sc_hd__a2bb2o_2 _12375_ (.A1_N(\coreWBInterface.readDataBuffered[12] ),
    .A2_N(net1316),
    .B1(_04640_),
    .B2(net1746),
    .X(_07097_));
 sky130_fd_sc_hd__nand2_1 _12376_ (.A(net579),
    .B(_07097_),
    .Y(_07098_));
 sky130_fd_sc_hd__o211a_1 _12377_ (.A1(\core.pipe0_currentInstruction[12] ),
    .A2(net579),
    .B1(_07098_),
    .C1(net1836),
    .X(_00142_));
 sky130_fd_sc_hd__a2bb2o_2 _12378_ (.A1_N(\coreWBInterface.readDataBuffered[13] ),
    .A2_N(net1316),
    .B1(_04554_),
    .B2(net1746),
    .X(_07099_));
 sky130_fd_sc_hd__nand2_1 _12379_ (.A(net578),
    .B(_07099_),
    .Y(_07100_));
 sky130_fd_sc_hd__o211a_1 _12380_ (.A1(\core.pipe0_currentInstruction[13] ),
    .A2(net576),
    .B1(_07100_),
    .C1(net1834),
    .X(_00143_));
 sky130_fd_sc_hd__a2bb2o_2 _12381_ (.A1_N(\coreWBInterface.readDataBuffered[14] ),
    .A2_N(net1316),
    .B1(_04468_),
    .B2(net1746),
    .X(_07101_));
 sky130_fd_sc_hd__nand2_1 _12382_ (.A(net576),
    .B(_07101_),
    .Y(_07102_));
 sky130_fd_sc_hd__o211a_1 _12383_ (.A1(\core.pipe0_currentInstruction[14] ),
    .A2(net576),
    .B1(_07102_),
    .C1(net1834),
    .X(_00144_));
 sky130_fd_sc_hd__o32a_1 _12384_ (.A1(net1635),
    .A2(_03989_),
    .A3(_03990_),
    .B1(net1315),
    .B2(\coreWBInterface.readDataBuffered[15] ),
    .X(_07103_));
 sky130_fd_sc_hd__or3_1 _12385_ (.A(\core.pipe0_fetch.currentPipeStall ),
    .B(net597),
    .C(_07103_),
    .X(_07104_));
 sky130_fd_sc_hd__o211a_1 _12386_ (.A1(\core.pipe0_currentInstruction[15] ),
    .A2(net579),
    .B1(_07104_),
    .C1(net1836),
    .X(_00145_));
 sky130_fd_sc_hd__o32ai_2 _12387_ (.A1(net1637),
    .A2(net1622),
    .A3(_04311_),
    .B1(net1317),
    .B2(\coreWBInterface.readDataBuffered[16] ),
    .Y(_07105_));
 sky130_fd_sc_hd__nand2_1 _12388_ (.A(net581),
    .B(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__o211a_1 _12389_ (.A1(net1792),
    .A2(net581),
    .B1(_07106_),
    .C1(net1858),
    .X(_00146_));
 sky130_fd_sc_hd__a2bb2o_1 _12390_ (.A1_N(\coreWBInterface.readDataBuffered[17] ),
    .A2_N(net1316),
    .B1(_04224_),
    .B2(net1746),
    .X(_07107_));
 sky130_fd_sc_hd__nand2_1 _12391_ (.A(net581),
    .B(_07107_),
    .Y(_07108_));
 sky130_fd_sc_hd__o211a_1 _12392_ (.A1(net1786),
    .A2(net581),
    .B1(_07108_),
    .C1(net1858),
    .X(_00147_));
 sky130_fd_sc_hd__o32ai_4 _12393_ (.A1(net1636),
    .A2(net1621),
    .A3(_04137_),
    .B1(net1317),
    .B2(\coreWBInterface.readDataBuffered[18] ),
    .Y(_07109_));
 sky130_fd_sc_hd__nand2_1 _12394_ (.A(net579),
    .B(_07109_),
    .Y(_07110_));
 sky130_fd_sc_hd__o211a_1 _12395_ (.A1(\core.pipe0_currentInstruction[18] ),
    .A2(net579),
    .B1(_07110_),
    .C1(net1836),
    .X(_00148_));
 sky130_fd_sc_hd__o32ai_2 _12396_ (.A1(net1636),
    .A2(net1622),
    .A3(_04023_),
    .B1(net1317),
    .B2(\coreWBInterface.readDataBuffered[19] ),
    .Y(_07111_));
 sky130_fd_sc_hd__nand2_1 _12397_ (.A(net583),
    .B(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__o211a_1 _12398_ (.A1(net1783),
    .A2(net583),
    .B1(_07112_),
    .C1(net1843),
    .X(_00149_));
 sky130_fd_sc_hd__o32ai_2 _12399_ (.A1(net1636),
    .A2(net1621),
    .A3(_04645_),
    .B1(net1317),
    .B2(\coreWBInterface.readDataBuffered[20] ),
    .Y(_07113_));
 sky130_fd_sc_hd__nand2_1 _12400_ (.A(net582),
    .B(_07113_),
    .Y(_07114_));
 sky130_fd_sc_hd__o211a_1 _12401_ (.A1(net1777),
    .A2(net582),
    .B1(_07114_),
    .C1(net1858),
    .X(_00150_));
 sky130_fd_sc_hd__o32ai_2 _12402_ (.A1(net1637),
    .A2(net1621),
    .A3(_04559_),
    .B1(net1316),
    .B2(\coreWBInterface.readDataBuffered[21] ),
    .Y(_07115_));
 sky130_fd_sc_hd__nand2_1 _12403_ (.A(net581),
    .B(_07115_),
    .Y(_07116_));
 sky130_fd_sc_hd__o211a_1 _12404_ (.A1(net1775),
    .A2(net581),
    .B1(_07116_),
    .C1(net1858),
    .X(_00151_));
 sky130_fd_sc_hd__o32ai_2 _12405_ (.A1(net1636),
    .A2(net1621),
    .A3(_04474_),
    .B1(net1316),
    .B2(\coreWBInterface.readDataBuffered[22] ),
    .Y(_07117_));
 sky130_fd_sc_hd__nand2_1 _12406_ (.A(net581),
    .B(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__o211a_1 _12407_ (.A1(net1766),
    .A2(net581),
    .B1(_07118_),
    .C1(net1858),
    .X(_00152_));
 sky130_fd_sc_hd__or2_1 _12408_ (.A(net1761),
    .B(net579),
    .X(_07119_));
 sky130_fd_sc_hd__o32a_1 _12409_ (.A1(net1635),
    .A2(net1622),
    .A3(_03996_),
    .B1(net1315),
    .B2(\coreWBInterface.readDataBuffered[23] ),
    .X(_07120_));
 sky130_fd_sc_hd__o311a_1 _12410_ (.A1(\core.pipe0_fetch.currentPipeStall ),
    .A2(net597),
    .A3(_07120_),
    .B1(_07119_),
    .C1(net1836),
    .X(_00153_));
 sky130_fd_sc_hd__o32ai_4 _12411_ (.A1(net1636),
    .A2(net1623),
    .A3(_04308_),
    .B1(net1317),
    .B2(\coreWBInterface.readDataBuffered[24] ),
    .Y(_07121_));
 sky130_fd_sc_hd__nand2_1 _12412_ (.A(net582),
    .B(_07121_),
    .Y(_07122_));
 sky130_fd_sc_hd__o211a_1 _12413_ (.A1(net1759),
    .A2(net582),
    .B1(_07122_),
    .C1(net1858),
    .X(_00154_));
 sky130_fd_sc_hd__a2bb2o_1 _12414_ (.A1_N(\coreWBInterface.readDataBuffered[25] ),
    .A2_N(net1316),
    .B1(_04220_),
    .B2(net1746),
    .X(_07123_));
 sky130_fd_sc_hd__nand2_1 _12415_ (.A(net583),
    .B(_07123_),
    .Y(_07124_));
 sky130_fd_sc_hd__o211a_1 _12416_ (.A1(\core.pipe0_currentInstruction[25] ),
    .A2(net583),
    .B1(_07124_),
    .C1(net1843),
    .X(_00155_));
 sky130_fd_sc_hd__o32ai_2 _12417_ (.A1(net1636),
    .A2(net1623),
    .A3(_04134_),
    .B1(net1317),
    .B2(\coreWBInterface.readDataBuffered[26] ),
    .Y(_07125_));
 sky130_fd_sc_hd__nand2_1 _12418_ (.A(net583),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__o211a_1 _12419_ (.A1(\core.pipe0_currentInstruction[26] ),
    .A2(net583),
    .B1(_07126_),
    .C1(net1843),
    .X(_00156_));
 sky130_fd_sc_hd__o32ai_4 _12420_ (.A1(net1637),
    .A2(net1624),
    .A3(_03976_),
    .B1(net1318),
    .B2(\coreWBInterface.readDataBuffered[27] ),
    .Y(_07127_));
 sky130_fd_sc_hd__nand2_1 _12421_ (.A(net580),
    .B(_07127_),
    .Y(_07128_));
 sky130_fd_sc_hd__o211a_1 _12422_ (.A1(\core.pipe0_currentInstruction[27] ),
    .A2(net580),
    .B1(_07128_),
    .C1(net1843),
    .X(_00157_));
 sky130_fd_sc_hd__o32ai_4 _12423_ (.A1(net1636),
    .A2(net1623),
    .A3(_04643_),
    .B1(net1316),
    .B2(\coreWBInterface.readDataBuffered[28] ),
    .Y(_07129_));
 sky130_fd_sc_hd__nand2_1 _12424_ (.A(net583),
    .B(_07129_),
    .Y(_07130_));
 sky130_fd_sc_hd__o211a_1 _12425_ (.A1(\core.pipe0_currentInstruction[28] ),
    .A2(net580),
    .B1(_07130_),
    .C1(net1843),
    .X(_00158_));
 sky130_fd_sc_hd__o32ai_4 _12426_ (.A1(net1636),
    .A2(net1624),
    .A3(_04557_),
    .B1(net1316),
    .B2(\coreWBInterface.readDataBuffered[29] ),
    .Y(_07131_));
 sky130_fd_sc_hd__nand2_1 _12427_ (.A(net583),
    .B(_07131_),
    .Y(_07132_));
 sky130_fd_sc_hd__o211a_1 _12428_ (.A1(\core.pipe0_currentInstruction[29] ),
    .A2(net583),
    .B1(_07132_),
    .C1(net1843),
    .X(_00159_));
 sky130_fd_sc_hd__o32ai_4 _12429_ (.A1(net1636),
    .A2(net1623),
    .A3(_04472_),
    .B1(net1316),
    .B2(\coreWBInterface.readDataBuffered[30] ),
    .Y(_07133_));
 sky130_fd_sc_hd__nand2_1 _12430_ (.A(net581),
    .B(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__o211a_1 _12431_ (.A1(net1752),
    .A2(net581),
    .B1(_07134_),
    .C1(net1858),
    .X(_00160_));
 sky130_fd_sc_hd__o32a_1 _12432_ (.A1(net1635),
    .A2(net1624),
    .A3(_03992_),
    .B1(net1315),
    .B2(\coreWBInterface.readDataBuffered[31] ),
    .X(_07135_));
 sky130_fd_sc_hd__or3_1 _12433_ (.A(\core.pipe0_fetch.currentPipeStall ),
    .B(net597),
    .C(_07135_),
    .X(_07136_));
 sky130_fd_sc_hd__o211a_1 _12434_ (.A1(net1751),
    .A2(net579),
    .B1(_07136_),
    .C1(net1836),
    .X(_00161_));
 sky130_fd_sc_hd__nor2_8 _12435_ (.A(_03861_),
    .B(net1275),
    .Y(_07137_));
 sky130_fd_sc_hd__and2_1 _12436_ (.A(_03863_),
    .B(_07137_),
    .X(_07138_));
 sky130_fd_sc_hd__nand2_1 _12437_ (.A(_03863_),
    .B(_07137_),
    .Y(_07139_));
 sky130_fd_sc_hd__or2_2 _12438_ (.A(\core.pipe0_currentInstruction[6] ),
    .B(_03860_),
    .X(_07140_));
 sky130_fd_sc_hd__nor2_4 _12439_ (.A(_03877_),
    .B(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__and2_2 _12440_ (.A(net1794),
    .B(_04059_),
    .X(_07142_));
 sky130_fd_sc_hd__nand2_1 _12441_ (.A(net1794),
    .B(_04059_),
    .Y(_07143_));
 sky130_fd_sc_hd__and4_2 _12442_ (.A(net1752),
    .B(net1629),
    .C(net1234),
    .D(net1218),
    .X(_07144_));
 sky130_fd_sc_hd__or4_4 _12443_ (.A(_03858_),
    .B(_04061_),
    .C(_07140_),
    .D(_07144_),
    .X(_07145_));
 sky130_fd_sc_hd__and2_4 _12444_ (.A(_04065_),
    .B(_07145_),
    .X(_07146_));
 sky130_fd_sc_hd__nand2_4 _12445_ (.A(_04065_),
    .B(_07145_),
    .Y(_07147_));
 sky130_fd_sc_hd__a211o_1 _12446_ (.A1(net1629),
    .A2(_04061_),
    .B1(_04055_),
    .C1(_03860_),
    .X(_07148_));
 sky130_fd_sc_hd__o21ai_4 _12447_ (.A1(_07144_),
    .A2(_07148_),
    .B1(_04065_),
    .Y(_07149_));
 sky130_fd_sc_hd__or4_4 _12448_ (.A(net1266),
    .B(net1133),
    .C(net1220),
    .D(_07147_),
    .X(_07150_));
 sky130_fd_sc_hd__o31a_2 _12449_ (.A1(net1151),
    .A2(net1122),
    .A3(_07150_),
    .B1(net1719),
    .X(_07151_));
 sky130_fd_sc_hd__o31ai_2 _12450_ (.A1(net1151),
    .A2(net1122),
    .A3(_07150_),
    .B1(net1719),
    .Y(_07152_));
 sky130_fd_sc_hd__and2_1 _12451_ (.A(net1794),
    .B(_07137_),
    .X(_07153_));
 sky130_fd_sc_hd__nand2_1 _12452_ (.A(net1795),
    .B(_07137_),
    .Y(_07154_));
 sky130_fd_sc_hd__mux2_1 _12453_ (.A0(net1793),
    .A1(_05049_),
    .S(net1114),
    .X(_07155_));
 sky130_fd_sc_hd__and2_2 _12454_ (.A(_04059_),
    .B(_07137_),
    .X(_07156_));
 sky130_fd_sc_hd__nand2_2 _12455_ (.A(_04059_),
    .B(_07137_),
    .Y(_07157_));
 sky130_fd_sc_hd__o21ai_2 _12456_ (.A1(_07037_),
    .A2(_07041_),
    .B1(net1713),
    .Y(_07158_));
 sky130_fd_sc_hd__nand2b_2 _12457_ (.A_N(_07021_),
    .B(_07023_),
    .Y(_07159_));
 sky130_fd_sc_hd__nor2_1 _12458_ (.A(_07158_),
    .B(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__or2_2 _12459_ (.A(_07158_),
    .B(_07159_),
    .X(_07161_));
 sky130_fd_sc_hd__nor2_1 _12460_ (.A(_03828_),
    .B(net1121),
    .Y(_07162_));
 sky130_fd_sc_hd__nand2_4 _12461_ (.A(net1719),
    .B(net1122),
    .Y(_07163_));
 sky130_fd_sc_hd__a21oi_4 _12462_ (.A1(net1726),
    .A2(net1071),
    .B1(net1021),
    .Y(_07164_));
 sky130_fd_sc_hd__a21o_4 _12463_ (.A1(net1725),
    .A2(net1071),
    .B1(net1021),
    .X(_07165_));
 sky130_fd_sc_hd__nand2_1 _12464_ (.A(net1714),
    .B(_07028_),
    .Y(_07166_));
 sky130_fd_sc_hd__a21bo_2 _12465_ (.A1(net1725),
    .A2(net1762),
    .B1_N(_07166_),
    .X(_07167_));
 sky130_fd_sc_hd__mux2_2 _12466_ (.A0(net1766),
    .A1(_07029_),
    .S(net1714),
    .X(_07168_));
 sky130_fd_sc_hd__nor2_4 _12467_ (.A(_07167_),
    .B(_07168_),
    .Y(_07169_));
 sky130_fd_sc_hd__nand2_2 _12468_ (.A(net1725),
    .B(net1690),
    .Y(_07170_));
 sky130_fd_sc_hd__o21a_4 _12469_ (.A1(net1725),
    .A2(_07033_),
    .B1(_07170_),
    .X(_07171_));
 sky130_fd_sc_hd__o21ai_4 _12470_ (.A1(net1725),
    .A2(_07033_),
    .B1(_07170_),
    .Y(_07172_));
 sky130_fd_sc_hd__mux2_8 _12471_ (.A0(net1775),
    .A1(_07032_),
    .S(net1714),
    .X(_07173_));
 sky130_fd_sc_hd__nor2_4 _12472_ (.A(_07171_),
    .B(_07173_),
    .Y(_07174_));
 sky130_fd_sc_hd__nand2_8 _12473_ (.A(_07169_),
    .B(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__nor2_2 _12474_ (.A(net1729),
    .B(_07013_),
    .Y(_07176_));
 sky130_fd_sc_hd__a21o_1 _12475_ (.A1(net1724),
    .A2(\core.pipe0_currentInstruction[28] ),
    .B1(_07176_),
    .X(_07177_));
 sky130_fd_sc_hd__nor2_1 _12476_ (.A(net1729),
    .B(_07015_),
    .Y(_07178_));
 sky130_fd_sc_hd__a21o_1 _12477_ (.A1(net1724),
    .A2(\core.pipe0_currentInstruction[29] ),
    .B1(_07178_),
    .X(_07179_));
 sky130_fd_sc_hd__nor2_2 _12478_ (.A(net1729),
    .B(_07017_),
    .Y(_07180_));
 sky130_fd_sc_hd__a21oi_1 _12479_ (.A1(net1726),
    .A2(_03833_),
    .B1(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__a21o_1 _12480_ (.A1(net1725),
    .A2(_03833_),
    .B1(_07180_),
    .X(_07182_));
 sky130_fd_sc_hd__or3_1 _12481_ (.A(_07177_),
    .B(_07179_),
    .C(_07181_),
    .X(_07183_));
 sky130_fd_sc_hd__mux2_2 _12482_ (.A0(\core.pipe0_currentInstruction[31] ),
    .A1(_07016_),
    .S(net1714),
    .X(_07184_));
 sky130_fd_sc_hd__nor2_2 _12483_ (.A(net1729),
    .B(_07014_),
    .Y(_07185_));
 sky130_fd_sc_hd__a21o_2 _12484_ (.A1(net1724),
    .A2(\core.pipe0_currentInstruction[30] ),
    .B1(_07185_),
    .X(_07186_));
 sky130_fd_sc_hd__nand2_1 _12485_ (.A(_07184_),
    .B(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__and2_1 _12486_ (.A(net1716),
    .B(_07022_),
    .X(_07188_));
 sky130_fd_sc_hd__a21o_1 _12487_ (.A1(net1724),
    .A2(\core.pipe0_currentInstruction[25] ),
    .B1(_07188_),
    .X(_07189_));
 sky130_fd_sc_hd__nand2_1 _12488_ (.A(net1724),
    .B(net1711),
    .Y(_07190_));
 sky130_fd_sc_hd__o21ai_2 _12489_ (.A1(net1724),
    .A2(_07024_),
    .B1(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__nand2b_2 _12490_ (.A_N(_07189_),
    .B(_07191_),
    .Y(_07192_));
 sky130_fd_sc_hd__or3_4 _12491_ (.A(_07183_),
    .B(_07187_),
    .C(_07192_),
    .X(_07193_));
 sky130_fd_sc_hd__and2_2 _12492_ (.A(net1716),
    .B(_07018_),
    .X(_07194_));
 sky130_fd_sc_hd__a21o_4 _12493_ (.A1(net1724),
    .A2(\core.pipe0_currentInstruction[27] ),
    .B1(_07194_),
    .X(_07195_));
 sky130_fd_sc_hd__or2_4 _12494_ (.A(_07193_),
    .B(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__nor2_4 _12495_ (.A(_07175_),
    .B(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__nand2b_4 _12496_ (.A_N(_07193_),
    .B(_07195_),
    .Y(_07198_));
 sky130_fd_sc_hd__nor2_4 _12497_ (.A(_07175_),
    .B(_07198_),
    .Y(_07199_));
 sky130_fd_sc_hd__a22o_1 _12498_ (.A1(\core.csr.cycleTimer.currentValue[0] ),
    .A2(net726),
    .B1(net722),
    .B2(\core.csr.cycleTimer.currentValue[32] ),
    .X(_07200_));
 sky130_fd_sc_hd__or4_4 _12499_ (.A(_07167_),
    .B(_07168_),
    .C(_07172_),
    .D(_07173_),
    .X(_07201_));
 sky130_fd_sc_hd__or2_4 _12500_ (.A(_07164_),
    .B(_07201_),
    .X(_07202_));
 sky130_fd_sc_hd__nand2_2 _12501_ (.A(_07177_),
    .B(_07179_),
    .Y(_07203_));
 sky130_fd_sc_hd__or2_1 _12502_ (.A(_07181_),
    .B(_07195_),
    .X(_07204_));
 sky130_fd_sc_hd__nor2_1 _12503_ (.A(_07203_),
    .B(_07204_),
    .Y(_07205_));
 sky130_fd_sc_hd__or4b_4 _12504_ (.A(_07187_),
    .B(_07189_),
    .C(_07191_),
    .D_N(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__nor2_4 _12505_ (.A(_07202_),
    .B(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__or2_4 _12506_ (.A(_07202_),
    .B(_07206_),
    .X(_07208_));
 sky130_fd_sc_hd__nand2_4 _12507_ (.A(_07169_),
    .B(_07173_),
    .Y(_07209_));
 sky130_fd_sc_hd__or2_4 _12508_ (.A(_07171_),
    .B(_07209_),
    .X(_07210_));
 sky130_fd_sc_hd__or2_4 _12509_ (.A(_07164_),
    .B(_07210_),
    .X(_07211_));
 sky130_fd_sc_hd__or2_4 _12510_ (.A(_07193_),
    .B(_07211_),
    .X(_07212_));
 sky130_fd_sc_hd__nor4_4 _12511_ (.A(_07184_),
    .B(_07186_),
    .C(_07192_),
    .D(_07203_),
    .Y(_07213_));
 sky130_fd_sc_hd__nand2b_4 _12512_ (.A_N(_07204_),
    .B(_07213_),
    .Y(_07214_));
 sky130_fd_sc_hd__and2b_1 _12513_ (.A_N(_07167_),
    .B(_07168_),
    .X(_07215_));
 sky130_fd_sc_hd__nand2_4 _12514_ (.A(_07174_),
    .B(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__or2_4 _12515_ (.A(_07164_),
    .B(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__nor2_1 _12516_ (.A(_07214_),
    .B(_07217_),
    .Y(_07218_));
 sky130_fd_sc_hd__or2_4 _12517_ (.A(_07214_),
    .B(_07217_),
    .X(_07219_));
 sky130_fd_sc_hd__or3b_4 _12518_ (.A(_07182_),
    .B(_07195_),
    .C_N(_07213_),
    .X(_07220_));
 sky130_fd_sc_hd__nor2_1 _12519_ (.A(_07217_),
    .B(_07220_),
    .Y(_07221_));
 sky130_fd_sc_hd__or2_4 _12520_ (.A(_07172_),
    .B(_07209_),
    .X(_07222_));
 sky130_fd_sc_hd__and3_1 _12521_ (.A(\core.csr.traps.mip.csrReadData[0] ),
    .B(_07221_),
    .C(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__a2111oi_1 _12522_ (.A1(_03809_),
    .A2(_07171_),
    .B1(_07209_),
    .C1(_07220_),
    .D1(_07164_),
    .Y(_07224_));
 sky130_fd_sc_hd__or2_4 _12523_ (.A(_07164_),
    .B(_07175_),
    .X(_07225_));
 sky130_fd_sc_hd__nor2_1 _12524_ (.A(_07220_),
    .B(_07225_),
    .Y(_07226_));
 sky130_fd_sc_hd__a21o_1 _12525_ (.A1(_07202_),
    .A2(_07225_),
    .B1(_07220_),
    .X(_07227_));
 sky130_fd_sc_hd__or3_1 _12526_ (.A(\core.csr.traps.mcause.csrReadData[0] ),
    .B(_07211_),
    .C(_07220_),
    .X(_07228_));
 sky130_fd_sc_hd__o211a_1 _12527_ (.A1(_07223_),
    .A2(_07224_),
    .B1(_07227_),
    .C1(_07228_),
    .X(_07229_));
 sky130_fd_sc_hd__or4b_4 _12528_ (.A(_07164_),
    .B(_07172_),
    .C(_07173_),
    .D_N(_07215_),
    .X(_07230_));
 sky130_fd_sc_hd__nor2_8 _12529_ (.A(_07214_),
    .B(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__a221o_1 _12530_ (.A1(\core.csr.traps.mscratch.currentValue[0] ),
    .A2(_07226_),
    .B1(_07231_),
    .B2(\core.csr.traps.mtvec.csrReadData[0] ),
    .C1(_07218_),
    .X(_07232_));
 sky130_fd_sc_hd__o22a_1 _12531_ (.A1(\core.csr.traps.mie.currentValue[0] ),
    .A2(_07219_),
    .B1(_07229_),
    .B2(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__nor2_2 _12532_ (.A(_07206_),
    .B(_07230_),
    .Y(_07234_));
 sky130_fd_sc_hd__nor2_1 _12533_ (.A(_07206_),
    .B(_07217_),
    .Y(_07235_));
 sky130_fd_sc_hd__a221o_4 _12534_ (.A1(\core.csr.mconfigptr.currentValue[0] ),
    .A2(net717),
    .B1(_07235_),
    .B2(net1),
    .C1(_07233_),
    .X(_07236_));
 sky130_fd_sc_hd__or2_4 _12535_ (.A(_07164_),
    .B(_07206_),
    .X(_07237_));
 sky130_fd_sc_hd__nor2_8 _12536_ (.A(_07210_),
    .B(_07237_),
    .Y(_07238_));
 sky130_fd_sc_hd__or2_4 _12537_ (.A(_07209_),
    .B(_07237_),
    .X(_07239_));
 sky130_fd_sc_hd__nor2_2 _12538_ (.A(_07172_),
    .B(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__a221o_1 _12539_ (.A1(net264),
    .A2(_07238_),
    .B1(_07240_),
    .B2(net280),
    .C1(_07207_),
    .X(_07241_));
 sky130_fd_sc_hd__o221a_1 _12540_ (.A1(net253),
    .A2(_07208_),
    .B1(_07236_),
    .B2(_07241_),
    .C1(_07212_),
    .X(_07242_));
 sky130_fd_sc_hd__nor2_1 _12541_ (.A(_07198_),
    .B(_07202_),
    .Y(_07243_));
 sky130_fd_sc_hd__nor2_1 _12542_ (.A(_07196_),
    .B(_07202_),
    .Y(_07244_));
 sky130_fd_sc_hd__or2_4 _12543_ (.A(_07196_),
    .B(_07202_),
    .X(_07245_));
 sky130_fd_sc_hd__nor2_4 _12544_ (.A(_07196_),
    .B(_07210_),
    .Y(_07246_));
 sky130_fd_sc_hd__nor2_4 _12545_ (.A(_07198_),
    .B(_07210_),
    .Y(_07247_));
 sky130_fd_sc_hd__a22o_1 _12546_ (.A1(\core.csr.instretTimer.currentValue[0] ),
    .A2(net702),
    .B1(net698),
    .B2(\core.csr.instretTimer.currentValue[32] ),
    .X(_07248_));
 sky130_fd_sc_hd__a221o_1 _12547_ (.A1(\core.csr.cycleTimer.currentValue[32] ),
    .A2(net716),
    .B1(_07248_),
    .B2(net978),
    .C1(net712),
    .X(_07249_));
 sky130_fd_sc_hd__or2_4 _12548_ (.A(_07193_),
    .B(_07225_),
    .X(_07250_));
 sky130_fd_sc_hd__o221a_1 _12549_ (.A1(\core.csr.cycleTimer.currentValue[0] ),
    .A2(net708),
    .B1(_07249_),
    .B2(_07242_),
    .C1(_07250_),
    .X(_07251_));
 sky130_fd_sc_hd__a21o_4 _12550_ (.A1(net978),
    .A2(_07200_),
    .B1(_07251_),
    .X(_07252_));
 sky130_fd_sc_hd__nor2_2 _12551_ (.A(_07216_),
    .B(_07237_),
    .Y(_07253_));
 sky130_fd_sc_hd__or2_2 _12552_ (.A(_07216_),
    .B(_07237_),
    .X(_07254_));
 sky130_fd_sc_hd__or4_1 _12553_ (.A(_07184_),
    .B(_07186_),
    .C(_07192_),
    .D(_07203_),
    .X(_07255_));
 sky130_fd_sc_hd__or3_4 _12554_ (.A(_07182_),
    .B(_07195_),
    .C(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__nor2_1 _12555_ (.A(_07211_),
    .B(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__nor2_1 _12556_ (.A(_07225_),
    .B(_07256_),
    .Y(_07258_));
 sky130_fd_sc_hd__or2_1 _12557_ (.A(_07225_),
    .B(_07256_),
    .X(_07259_));
 sky130_fd_sc_hd__nor2_1 _12558_ (.A(_07202_),
    .B(_07256_),
    .Y(_07260_));
 sky130_fd_sc_hd__or2_1 _12559_ (.A(_07202_),
    .B(_07256_),
    .X(_07261_));
 sky130_fd_sc_hd__nand2_1 _12560_ (.A(net693),
    .B(net687),
    .Y(_07262_));
 sky130_fd_sc_hd__or2_1 _12561_ (.A(_07164_),
    .B(_07256_),
    .X(_07263_));
 sky130_fd_sc_hd__or2_1 _12562_ (.A(_07222_),
    .B(_07263_),
    .X(_07264_));
 sky130_fd_sc_hd__or2_4 _12563_ (.A(_07204_),
    .B(_07255_),
    .X(_07265_));
 sky130_fd_sc_hd__nor2_1 _12564_ (.A(_07217_),
    .B(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__or2_1 _12565_ (.A(_07217_),
    .B(_07265_),
    .X(_07267_));
 sky130_fd_sc_hd__nor2_1 _12566_ (.A(_07230_),
    .B(_07265_),
    .Y(_07268_));
 sky130_fd_sc_hd__nor2_2 _12567_ (.A(_07225_),
    .B(_07265_),
    .Y(_07269_));
 sky130_fd_sc_hd__inv_2 _12568_ (.A(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__a21oi_1 _12569_ (.A1(_07216_),
    .A2(_07222_),
    .B1(_07263_),
    .Y(_07271_));
 sky130_fd_sc_hd__or4_1 _12570_ (.A(net666),
    .B(_07262_),
    .C(net684),
    .D(_07269_),
    .X(_07272_));
 sky130_fd_sc_hd__o31a_1 _12571_ (.A1(net678),
    .A2(net660),
    .A3(_07272_),
    .B1(_07270_),
    .X(_07273_));
 sky130_fd_sc_hd__or4b_4 _12572_ (.A(_07187_),
    .B(_07189_),
    .C(_07191_),
    .D_N(_07205_),
    .X(_07274_));
 sky130_fd_sc_hd__or2_2 _12573_ (.A(_07164_),
    .B(_07274_),
    .X(_07275_));
 sky130_fd_sc_hd__nor2_4 _12574_ (.A(_07201_),
    .B(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__nor2_8 _12575_ (.A(_07211_),
    .B(_07274_),
    .Y(_07277_));
 sky130_fd_sc_hd__or2_4 _12576_ (.A(_07209_),
    .B(_07275_),
    .X(_07278_));
 sky130_fd_sc_hd__or2_4 _12577_ (.A(_07164_),
    .B(_07220_),
    .X(_07279_));
 sky130_fd_sc_hd__nor2_4 _12578_ (.A(_07175_),
    .B(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__nor2_8 _12579_ (.A(_07210_),
    .B(_07279_),
    .Y(_07281_));
 sky130_fd_sc_hd__nor2_1 _12580_ (.A(_07222_),
    .B(_07279_),
    .Y(_07282_));
 sky130_fd_sc_hd__nor2_8 _12581_ (.A(_07201_),
    .B(_07279_),
    .Y(_07283_));
 sky130_fd_sc_hd__or2_4 _12582_ (.A(_07201_),
    .B(_07279_),
    .X(_07284_));
 sky130_fd_sc_hd__nor2_8 _12583_ (.A(_07230_),
    .B(_07274_),
    .Y(_07285_));
 sky130_fd_sc_hd__nor2_2 _12584_ (.A(_07217_),
    .B(_07274_),
    .Y(_07286_));
 sky130_fd_sc_hd__a21o_1 _12585_ (.A1(net1111),
    .A2(_07252_),
    .B1(_07155_),
    .X(_07287_));
 sky130_fd_sc_hd__and2_4 _12586_ (.A(_04049_),
    .B(_07137_),
    .X(_07288_));
 sky130_fd_sc_hd__nand2_2 _12587_ (.A(_04049_),
    .B(_07137_),
    .Y(_07289_));
 sky130_fd_sc_hd__o21ai_2 _12588_ (.A1(_04051_),
    .A2(_04059_),
    .B1(_07137_),
    .Y(_07290_));
 sky130_fd_sc_hd__o21a_1 _12589_ (.A1(_04051_),
    .A2(_04059_),
    .B1(_07137_),
    .X(_07291_));
 sky130_fd_sc_hd__o21ai_1 _12590_ (.A1(_07155_),
    .A2(net1108),
    .B1(net1107),
    .Y(_07292_));
 sky130_fd_sc_hd__a31o_1 _12591_ (.A1(net1122),
    .A2(_07287_),
    .A3(_07292_),
    .B1(net1151),
    .X(_07293_));
 sky130_fd_sc_hd__o21a_1 _12592_ (.A1(_04068_),
    .A2(net671),
    .B1(_07293_),
    .X(_07294_));
 sky130_fd_sc_hd__nor2_1 _12593_ (.A(_06050_),
    .B(_06661_),
    .Y(_07295_));
 sky130_fd_sc_hd__or2_1 _12594_ (.A(_06014_),
    .B(_06046_),
    .X(_07296_));
 sky130_fd_sc_hd__nor2_2 _12595_ (.A(_06247_),
    .B(_06278_),
    .Y(_07297_));
 sky130_fd_sc_hd__nor2_2 _12596_ (.A(_06323_),
    .B(_06354_),
    .Y(_07298_));
 sky130_fd_sc_hd__nor2_1 _12597_ (.A(_06400_),
    .B(_06430_),
    .Y(_07299_));
 sky130_fd_sc_hd__or2_1 _12598_ (.A(_04045_),
    .B(_04130_),
    .X(_07300_));
 sky130_fd_sc_hd__nand2_1 _12599_ (.A(_04180_),
    .B(_04214_),
    .Y(_07301_));
 sky130_fd_sc_hd__and2_1 _12600_ (.A(_04268_),
    .B(_04303_),
    .X(_07302_));
 sky130_fd_sc_hd__nand2_1 _12601_ (.A(net748),
    .B(_04802_),
    .Y(_07303_));
 sky130_fd_sc_hd__or2_1 _12602_ (.A(_04852_),
    .B(_04883_),
    .X(_07304_));
 sky130_fd_sc_hd__or2_2 _12603_ (.A(net885),
    .B(_05050_),
    .X(_07305_));
 sky130_fd_sc_hd__nand2_1 _12604_ (.A(_04972_),
    .B(_07305_),
    .Y(_07306_));
 sky130_fd_sc_hd__a22oi_4 _12605_ (.A1(net889),
    .A2(_04969_),
    .B1(_04972_),
    .B2(_07305_),
    .Y(_07307_));
 sky130_fd_sc_hd__o21a_2 _12606_ (.A1(_06712_),
    .A2(_07307_),
    .B1(_07304_),
    .X(_07308_));
 sky130_fd_sc_hd__o21a_1 _12607_ (.A1(_06714_),
    .A2(_07308_),
    .B1(_07303_),
    .X(_07309_));
 sky130_fd_sc_hd__a21o_1 _12608_ (.A1(_04721_),
    .A2(_04723_),
    .B1(_07309_),
    .X(_07310_));
 sky130_fd_sc_hd__nand2_1 _12609_ (.A(_04687_),
    .B(_04720_),
    .Y(_07311_));
 sky130_fd_sc_hd__nand2_1 _12610_ (.A(_07310_),
    .B(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__or2_1 _12611_ (.A(_06719_),
    .B(_06721_),
    .X(_07313_));
 sky130_fd_sc_hd__nand2b_1 _12612_ (.A_N(_04461_),
    .B(_04424_),
    .Y(_07314_));
 sky130_fd_sc_hd__nand2b_1 _12613_ (.A_N(_04547_),
    .B(_04513_),
    .Y(_07315_));
 sky130_fd_sc_hd__nand2b_1 _12614_ (.A_N(_04632_),
    .B(_04598_),
    .Y(_07316_));
 sky130_fd_sc_hd__or4bb_2 _12615_ (.A(_07313_),
    .B(_07309_),
    .C_N(_04724_),
    .D_N(_04636_),
    .X(_07317_));
 sky130_fd_sc_hd__o21a_1 _12616_ (.A1(_04635_),
    .A2(_07311_),
    .B1(_07316_),
    .X(_07318_));
 sky130_fd_sc_hd__o221a_1 _12617_ (.A1(_06721_),
    .A2(_07315_),
    .B1(_07318_),
    .B2(_07313_),
    .C1(_07314_),
    .X(_07319_));
 sky130_fd_sc_hd__a21oi_2 _12618_ (.A1(_07317_),
    .A2(_07319_),
    .B1(_04391_),
    .Y(_07320_));
 sky130_fd_sc_hd__o21ba_1 _12619_ (.A1(_04353_),
    .A2(_04354_),
    .B1_N(_04388_),
    .X(_07321_));
 sky130_fd_sc_hd__o21a_1 _12620_ (.A1(_07320_),
    .A2(_07321_),
    .B1(_04306_),
    .X(_07322_));
 sky130_fd_sc_hd__o21ai_2 _12621_ (.A1(_07302_),
    .A2(_07322_),
    .B1(_04218_),
    .Y(_07323_));
 sky130_fd_sc_hd__nand2_1 _12622_ (.A(_07301_),
    .B(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__a21o_1 _12623_ (.A1(_07301_),
    .A2(_07323_),
    .B1(_04133_),
    .X(_07325_));
 sky130_fd_sc_hd__nand2_1 _12624_ (.A(_07300_),
    .B(_07325_),
    .Y(_07326_));
 sky130_fd_sc_hd__nor2_1 _12625_ (.A(_06477_),
    .B(_06507_),
    .Y(_07327_));
 sky130_fd_sc_hd__or4_1 _12626_ (.A(_06281_),
    .B(_06357_),
    .C(_06434_),
    .D(_06511_),
    .X(_07328_));
 sky130_fd_sc_hd__a21o_2 _12627_ (.A1(_07300_),
    .A2(_07325_),
    .B1(_07328_),
    .X(_07329_));
 sky130_fd_sc_hd__o21a_1 _12628_ (.A1(_06432_),
    .A2(_06433_),
    .B1(_07327_),
    .X(_07330_));
 sky130_fd_sc_hd__o211a_1 _12629_ (.A1(_07299_),
    .A2(_07330_),
    .B1(_06282_),
    .C1(_06358_),
    .X(_07331_));
 sky130_fd_sc_hd__a211oi_4 _12630_ (.A1(_06282_),
    .A2(_07298_),
    .B1(_07331_),
    .C1(_07297_),
    .Y(_07332_));
 sky130_fd_sc_hd__a21oi_4 _12631_ (.A1(_07329_),
    .A2(_07332_),
    .B1(_06203_),
    .Y(_07333_));
 sky130_fd_sc_hd__o32a_1 _12632_ (.A1(_06127_),
    .A2(_06169_),
    .A3(_06200_),
    .B1(_06124_),
    .B2(_06092_),
    .X(_07334_));
 sky130_fd_sc_hd__o21a_1 _12633_ (.A1(_06050_),
    .A2(_07334_),
    .B1(_07296_),
    .X(_07335_));
 sky130_fd_sc_hd__or2_1 _12634_ (.A(_06661_),
    .B(_07335_),
    .X(_07336_));
 sky130_fd_sc_hd__o21ai_1 _12635_ (.A1(_05938_),
    .A2(_05970_),
    .B1(_07336_),
    .Y(_07337_));
 sky130_fd_sc_hd__a31o_2 _12636_ (.A1(_06128_),
    .A2(_07295_),
    .A3(_07333_),
    .B1(_07337_),
    .X(_07338_));
 sky130_fd_sc_hd__nand2b_1 _12637_ (.A_N(_05897_),
    .B(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__nor4_1 _12638_ (.A(_05742_),
    .B(_05897_),
    .C(_06525_),
    .D(_06529_),
    .Y(_07340_));
 sky130_fd_sc_hd__nand2b_2 _12639_ (.A_N(_05704_),
    .B(_05739_),
    .Y(_07341_));
 sky130_fd_sc_hd__nand2b_1 _12640_ (.A_N(_05782_),
    .B(_05817_),
    .Y(_07342_));
 sky130_fd_sc_hd__or2_1 _12641_ (.A(_05862_),
    .B(_05894_),
    .X(_07343_));
 sky130_fd_sc_hd__o21ai_1 _12642_ (.A1(_06525_),
    .A2(_07343_),
    .B1(_07342_),
    .Y(_07344_));
 sky130_fd_sc_hd__nand2_1 _12643_ (.A(_05743_),
    .B(_07344_),
    .Y(_07345_));
 sky130_fd_sc_hd__a21oi_1 _12644_ (.A1(_07341_),
    .A2(_07345_),
    .B1(_06529_),
    .Y(_07346_));
 sky130_fd_sc_hd__a21o_1 _12645_ (.A1(_05628_),
    .A2(_05663_),
    .B1(_07346_),
    .X(_07347_));
 sky130_fd_sc_hd__a21o_4 _12646_ (.A1(_07338_),
    .A2(_07340_),
    .B1(_07347_),
    .X(_07348_));
 sky130_fd_sc_hd__nor3_1 _12647_ (.A(_05591_),
    .B(_06533_),
    .C(_06538_),
    .Y(_07349_));
 sky130_fd_sc_hd__and2b_1 _12648_ (.A_N(_05404_),
    .B(_05439_),
    .X(_07350_));
 sky130_fd_sc_hd__and2b_1 _12649_ (.A_N(_05478_),
    .B(_05513_),
    .X(_07351_));
 sky130_fd_sc_hd__and2b_1 _12650_ (.A_N(_05553_),
    .B(_05588_),
    .X(_07352_));
 sky130_fd_sc_hd__a21o_1 _12651_ (.A1(_06534_),
    .A2(_07352_),
    .B1(_07351_),
    .X(_07353_));
 sky130_fd_sc_hd__a21oi_1 _12652_ (.A1(_05442_),
    .A2(_07353_),
    .B1(_07350_),
    .Y(_07354_));
 sky130_fd_sc_hd__nand2b_1 _12653_ (.A_N(_05331_),
    .B(_05366_),
    .Y(_07355_));
 sky130_fd_sc_hd__o21ai_1 _12654_ (.A1(_06538_),
    .A2(_07354_),
    .B1(_07355_),
    .Y(_07356_));
 sky130_fd_sc_hd__a31o_4 _12655_ (.A1(_05442_),
    .A2(_07348_),
    .A3(_07349_),
    .B1(_07356_),
    .X(_07357_));
 sky130_fd_sc_hd__and4_1 _12656_ (.A(_05148_),
    .B(_06617_),
    .C(_06622_),
    .D(_06624_),
    .X(_07358_));
 sky130_fd_sc_hd__nand2b_1 _12657_ (.A_N(_05185_),
    .B(_05218_),
    .Y(_07359_));
 sky130_fd_sc_hd__nand2b_1 _12658_ (.A_N(_05260_),
    .B(_05293_),
    .Y(_07360_));
 sky130_fd_sc_hd__o21ai_2 _12659_ (.A1(_06621_),
    .A2(_07360_),
    .B1(_07359_),
    .Y(_07361_));
 sky130_fd_sc_hd__and2b_1 _12660_ (.A_N(_05110_),
    .B(_05145_),
    .X(_07362_));
 sky130_fd_sc_hd__a21o_1 _12661_ (.A1(_05148_),
    .A2(_07361_),
    .B1(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__a22oi_4 _12662_ (.A1(_07357_),
    .A2(_07358_),
    .B1(_07363_),
    .B2(_06616_),
    .Y(_07364_));
 sky130_fd_sc_hd__nand2b_1 _12663_ (.A_N(_06615_),
    .B(_07364_),
    .Y(_07365_));
 sky130_fd_sc_hd__a21oi_2 _12664_ (.A1(_06616_),
    .A2(_07364_),
    .B1(_06615_),
    .Y(_07366_));
 sky130_fd_sc_hd__or3_1 _12665_ (.A(_03843_),
    .B(_04052_),
    .C(_07365_),
    .X(_07367_));
 sky130_fd_sc_hd__nor2_4 _12666_ (.A(net1794),
    .B(_04060_),
    .Y(_07368_));
 sky130_fd_sc_hd__or2_4 _12667_ (.A(net1794),
    .B(_04060_),
    .X(_07369_));
 sky130_fd_sc_hd__mux2_1 _12668_ (.A0(_04214_),
    .A1(_05817_),
    .S(net1214),
    .X(_07370_));
 sky130_fd_sc_hd__mux2_2 _12669_ (.A0(_04046_),
    .A1(_05893_),
    .S(net1213),
    .X(_07371_));
 sky130_fd_sc_hd__mux2_1 _12670_ (.A0(_07371_),
    .A1(_07370_),
    .S(net881),
    .X(_07372_));
 sky130_fd_sc_hd__or2_1 _12671_ (.A(_05662_),
    .B(net1209),
    .X(_07373_));
 sky130_fd_sc_hd__o21ai_1 _12672_ (.A1(_04388_),
    .A2(net1214),
    .B1(_07373_),
    .Y(_07374_));
 sky130_fd_sc_hd__mux2_1 _12673_ (.A0(_04303_),
    .A1(_05739_),
    .S(net1214),
    .X(_07375_));
 sky130_fd_sc_hd__mux2_1 _12674_ (.A0(_07375_),
    .A1(_07374_),
    .S(net883),
    .X(_07376_));
 sky130_fd_sc_hd__mux2_1 _12675_ (.A0(_07372_),
    .A1(_07376_),
    .S(net886),
    .X(_07377_));
 sky130_fd_sc_hd__mux2_1 _12676_ (.A0(_06124_),
    .A1(_06354_),
    .S(net1209),
    .X(_07378_));
 sky130_fd_sc_hd__mux2_1 _12677_ (.A0(_06200_),
    .A1(_06278_),
    .S(net1209),
    .X(_07379_));
 sky130_fd_sc_hd__mux2_1 _12678_ (.A0(_07379_),
    .A1(_07378_),
    .S(net882),
    .X(_07380_));
 sky130_fd_sc_hd__mux2_4 _12679_ (.A0(_05970_),
    .A1(_06507_),
    .S(net1210),
    .X(_07381_));
 sky130_fd_sc_hd__inv_2 _12680_ (.A(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__mux2_4 _12681_ (.A0(_06046_),
    .A1(_06430_),
    .S(net1211),
    .X(_07383_));
 sky130_fd_sc_hd__mux2_1 _12682_ (.A0(_07383_),
    .A1(_07381_),
    .S(net881),
    .X(_07384_));
 sky130_fd_sc_hd__or2_1 _12683_ (.A(net744),
    .B(_07384_),
    .X(_07385_));
 sky130_fd_sc_hd__o21ai_1 _12684_ (.A1(net886),
    .A2(_07380_),
    .B1(_07385_),
    .Y(_07386_));
 sky130_fd_sc_hd__mux2_1 _12685_ (.A0(_07377_),
    .A1(_07386_),
    .S(net893),
    .X(_07387_));
 sky130_fd_sc_hd__mux2_1 _12686_ (.A0(_04884_),
    .A1(_05218_),
    .S(net1213),
    .X(_07388_));
 sky130_fd_sc_hd__mux2_2 _12687_ (.A0(_04802_),
    .A1(_05293_),
    .S(net1213),
    .X(_07389_));
 sky130_fd_sc_hd__mux2_2 _12688_ (.A0(_07389_),
    .A1(_07388_),
    .S(net885),
    .X(_07390_));
 sky130_fd_sc_hd__mux2_1 _12689_ (.A0(_04969_),
    .A1(_05145_),
    .S(net1213),
    .X(_07391_));
 sky130_fd_sc_hd__mux2_1 _12690_ (.A0(_05050_),
    .A1(_06614_),
    .S(net1213),
    .X(_07392_));
 sky130_fd_sc_hd__mux2_1 _12691_ (.A0(_07391_),
    .A1(_07392_),
    .S(net885),
    .X(_07393_));
 sky130_fd_sc_hd__mux2_1 _12692_ (.A0(_07390_),
    .A1(_07393_),
    .S(net887),
    .X(_07394_));
 sky130_fd_sc_hd__mux2_1 _12693_ (.A0(_04513_),
    .A1(_05513_),
    .S(net1214),
    .X(_07395_));
 sky130_fd_sc_hd__mux2_1 _12694_ (.A0(_04424_),
    .A1(_05588_),
    .S(net1214),
    .X(_07396_));
 sky130_fd_sc_hd__mux2_1 _12695_ (.A0(_07396_),
    .A1(_07395_),
    .S(net883),
    .X(_07397_));
 sky130_fd_sc_hd__mux2_1 _12696_ (.A0(_04720_),
    .A1(_05366_),
    .S(net1213),
    .X(_07398_));
 sky130_fd_sc_hd__mux2_1 _12697_ (.A0(_04598_),
    .A1(_05439_),
    .S(net1214),
    .X(_07399_));
 sky130_fd_sc_hd__mux2_1 _12698_ (.A0(_07399_),
    .A1(_07398_),
    .S(net883),
    .X(_07400_));
 sky130_fd_sc_hd__mux2_1 _12699_ (.A0(_07397_),
    .A1(_07400_),
    .S(net887),
    .X(_07401_));
 sky130_fd_sc_hd__mux2_1 _12700_ (.A0(_07394_),
    .A1(_07401_),
    .S(net894),
    .X(_07402_));
 sky130_fd_sc_hd__mux2_2 _12701_ (.A0(_07387_),
    .A1(_07402_),
    .S(net746),
    .X(_07403_));
 sky130_fd_sc_hd__inv_2 _12702_ (.A(_07403_),
    .Y(_07404_));
 sky130_fd_sc_hd__mux2_1 _12703_ (.A0(_04802_),
    .A1(_05293_),
    .S(net1210),
    .X(_07405_));
 sky130_fd_sc_hd__mux2_1 _12704_ (.A0(_04884_),
    .A1(_05218_),
    .S(net1210),
    .X(_07406_));
 sky130_fd_sc_hd__mux2_1 _12705_ (.A0(_07406_),
    .A1(_07405_),
    .S(net884),
    .X(_07407_));
 sky130_fd_sc_hd__or2_1 _12706_ (.A(_06613_),
    .B(net1213),
    .X(_07408_));
 sky130_fd_sc_hd__a21bo_1 _12707_ (.A1(_05050_),
    .A2(net1213),
    .B1_N(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__mux2_1 _12708_ (.A0(_04969_),
    .A1(_05145_),
    .S(net1211),
    .X(_07410_));
 sky130_fd_sc_hd__mux2_1 _12709_ (.A0(_07409_),
    .A1(_07410_),
    .S(net884),
    .X(_07411_));
 sky130_fd_sc_hd__mux2_1 _12710_ (.A0(_07407_),
    .A1(_07411_),
    .S(net745),
    .X(_07412_));
 sky130_fd_sc_hd__mux2_1 _12711_ (.A0(_04598_),
    .A1(_05439_),
    .S(net1207),
    .X(_07413_));
 sky130_fd_sc_hd__mux2_1 _12712_ (.A0(_04720_),
    .A1(_05366_),
    .S(net1208),
    .X(_07414_));
 sky130_fd_sc_hd__mux2_1 _12713_ (.A0(_07414_),
    .A1(_07413_),
    .S(net884),
    .X(_07415_));
 sky130_fd_sc_hd__mux2_1 _12714_ (.A0(_04424_),
    .A1(_05588_),
    .S(net1209),
    .X(_07416_));
 sky130_fd_sc_hd__mux2_1 _12715_ (.A0(_04513_),
    .A1(_05513_),
    .S(net1209),
    .X(_07417_));
 sky130_fd_sc_hd__mux2_1 _12716_ (.A0(_07417_),
    .A1(_07416_),
    .S(net883),
    .X(_07418_));
 sky130_fd_sc_hd__mux2_1 _12717_ (.A0(_07415_),
    .A1(_07418_),
    .S(net888),
    .X(_07419_));
 sky130_fd_sc_hd__mux2_1 _12718_ (.A0(_07412_),
    .A1(_07419_),
    .S(net891),
    .X(_07420_));
 sky130_fd_sc_hd__or2_1 _12719_ (.A(net747),
    .B(_07420_),
    .X(_07421_));
 sky130_fd_sc_hd__mux2_4 _12720_ (.A0(_06045_),
    .A1(_06431_),
    .S(_07368_),
    .X(_07422_));
 sky130_fd_sc_hd__mux2_4 _12721_ (.A0(_05969_),
    .A1(_06508_),
    .S(_07368_),
    .X(_07423_));
 sky130_fd_sc_hd__mux2_1 _12722_ (.A0(_07423_),
    .A1(_07422_),
    .S(net881),
    .X(_07424_));
 sky130_fd_sc_hd__mux2_1 _12723_ (.A0(_06200_),
    .A1(_06278_),
    .S(net1214),
    .X(_07425_));
 sky130_fd_sc_hd__mux2_1 _12724_ (.A0(_06124_),
    .A1(_06354_),
    .S(net1214),
    .X(_07426_));
 sky130_fd_sc_hd__mux2_1 _12725_ (.A0(_07426_),
    .A1(_07425_),
    .S(net882),
    .X(_07427_));
 sky130_fd_sc_hd__inv_2 _12726_ (.A(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__mux2_1 _12727_ (.A0(_07424_),
    .A1(_07428_),
    .S(net886),
    .X(_07429_));
 sky130_fd_sc_hd__mux2_1 _12728_ (.A0(_04303_),
    .A1(_05739_),
    .S(net1209),
    .X(_07430_));
 sky130_fd_sc_hd__or2_1 _12729_ (.A(_05662_),
    .B(net1214),
    .X(_07431_));
 sky130_fd_sc_hd__o21ai_1 _12730_ (.A1(_04388_),
    .A2(net1209),
    .B1(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__mux2_1 _12731_ (.A0(_07432_),
    .A1(_07430_),
    .S(net881),
    .X(_07433_));
 sky130_fd_sc_hd__mux2_2 _12732_ (.A0(_04045_),
    .A1(_05894_),
    .S(net1207),
    .X(_07434_));
 sky130_fd_sc_hd__mux2_1 _12733_ (.A0(_04214_),
    .A1(_05817_),
    .S(net1209),
    .X(_07435_));
 sky130_fd_sc_hd__nor2_1 _12734_ (.A(net882),
    .B(_07435_),
    .Y(_07436_));
 sky130_fd_sc_hd__a21oi_1 _12735_ (.A1(net881),
    .A2(_07434_),
    .B1(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__mux2_1 _12736_ (.A0(_07433_),
    .A1(_07437_),
    .S(net886),
    .X(_07438_));
 sky130_fd_sc_hd__mux2_2 _12737_ (.A0(_07429_),
    .A1(_07438_),
    .S(net893),
    .X(_07439_));
 sky130_fd_sc_hd__o21ai_2 _12738_ (.A1(net750),
    .A2(_07439_),
    .B1(_07421_),
    .Y(_07440_));
 sky130_fd_sc_hd__mux2_2 _12739_ (.A0(_07404_),
    .A1(_07440_),
    .S(net756),
    .X(_07441_));
 sky130_fd_sc_hd__or3_2 _12740_ (.A(_04058_),
    .B(_04060_),
    .C(_04064_),
    .X(_07442_));
 sky130_fd_sc_hd__a21oi_1 _12741_ (.A1(_07145_),
    .A2(_07442_),
    .B1(_04063_),
    .Y(_07443_));
 sky130_fd_sc_hd__a21o_4 _12742_ (.A1(_07145_),
    .A2(_07442_),
    .B1(_04063_),
    .X(_07444_));
 sky130_fd_sc_hd__nor2_2 _12743_ (.A(_07408_),
    .B(net1060),
    .Y(_07445_));
 sky130_fd_sc_hd__nor2_1 _12744_ (.A(net753),
    .B(_07445_),
    .Y(_07446_));
 sky130_fd_sc_hd__or2_4 _12745_ (.A(net747),
    .B(_07445_),
    .X(_07447_));
 sky130_fd_sc_hd__or2_2 _12746_ (.A(net892),
    .B(_07445_),
    .X(_07448_));
 sky130_fd_sc_hd__o21ai_2 _12747_ (.A1(net884),
    .A2(net1064),
    .B1(_07409_),
    .Y(_07449_));
 sky130_fd_sc_hd__inv_2 _12748_ (.A(_07449_),
    .Y(_07450_));
 sky130_fd_sc_hd__mux2_1 _12749_ (.A0(_07445_),
    .A1(_07450_),
    .S(net888),
    .X(_07451_));
 sky130_fd_sc_hd__o21a_1 _12750_ (.A1(net895),
    .A2(_07451_),
    .B1(_07448_),
    .X(_07452_));
 sky130_fd_sc_hd__o21ai_2 _12751_ (.A1(net750),
    .A2(_07452_),
    .B1(_07447_),
    .Y(_07453_));
 sky130_fd_sc_hd__a21o_1 _12752_ (.A1(net753),
    .A2(_07453_),
    .B1(net631),
    .X(_07454_));
 sky130_fd_sc_hd__and2_2 _12753_ (.A(net1795),
    .B(_04051_),
    .X(_07455_));
 sky130_fd_sc_hd__nand2_2 _12754_ (.A(net1795),
    .B(_04051_),
    .Y(_07456_));
 sky130_fd_sc_hd__and2_2 _12755_ (.A(net1795),
    .B(_04049_),
    .X(_07457_));
 sky130_fd_sc_hd__nand2_8 _12756_ (.A(net1794),
    .B(_04049_),
    .Y(_07458_));
 sky130_fd_sc_hd__o22a_1 _12757_ (.A1(net1218),
    .A2(_07441_),
    .B1(_07454_),
    .B2(net1211),
    .X(_07459_));
 sky130_fd_sc_hd__o221a_1 _12758_ (.A1(_06636_),
    .A2(net1204),
    .B1(_07458_),
    .B2(_05052_),
    .C1(_07459_),
    .X(_07460_));
 sky130_fd_sc_hd__o22a_1 _12759_ (.A1(net669),
    .A2(_06645_),
    .B1(_07366_),
    .B2(_04053_),
    .X(_07461_));
 sky130_fd_sc_hd__a31oi_2 _12760_ (.A1(_07367_),
    .A2(_07460_),
    .A3(_07461_),
    .B1(_07146_),
    .Y(_07462_));
 sky130_fd_sc_hd__or4_2 _12761_ (.A(net1266),
    .B(net1133),
    .C(_07294_),
    .D(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__nor2_2 _12762_ (.A(_07141_),
    .B(net983),
    .Y(_07464_));
 sky130_fd_sc_hd__a31o_1 _12763_ (.A1(net1262),
    .A2(net1226),
    .A3(net1181),
    .B1(net450),
    .X(_07465_));
 sky130_fd_sc_hd__a32o_1 _12764_ (.A1(_07463_),
    .A2(net825),
    .A3(_07465_),
    .B1(net984),
    .B2(\core.pipe1_resultRegister[0] ),
    .X(_07466_));
 sky130_fd_sc_hd__and2_1 _12765_ (.A(net1822),
    .B(_07466_),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _12766_ (.A0(net1666),
    .A1(_04968_),
    .S(net1114),
    .X(_07467_));
 sky130_fd_sc_hd__a22o_1 _12767_ (.A1(\core.csr.cycleTimer.currentValue[1] ),
    .A2(net726),
    .B1(net722),
    .B2(\core.csr.cycleTimer.currentValue[33] ),
    .X(_07468_));
 sky130_fd_sc_hd__or2_1 _12768_ (.A(_07214_),
    .B(_07225_),
    .X(_07469_));
 sky130_fd_sc_hd__a22o_1 _12769_ (.A1(\core.csr.instretTimer.currentValue[1] ),
    .A2(net703),
    .B1(net699),
    .B2(\core.csr.instretTimer.currentValue[33] ),
    .X(_07470_));
 sky130_fd_sc_hd__and2_1 _12770_ (.A(net281),
    .B(_07171_),
    .X(_07471_));
 sky130_fd_sc_hd__or2_4 _12771_ (.A(_07221_),
    .B(net657),
    .X(_07472_));
 sky130_fd_sc_hd__mux2_1 _12772_ (.A0(\core.csr.traps.mip.csrReadData[1] ),
    .A1(\core.csr.traps.mtval.csrReadData[1] ),
    .S(net656),
    .X(_07473_));
 sky130_fd_sc_hd__a221o_1 _12773_ (.A1(\core.csr.traps.mcause.csrReadData[1] ),
    .A2(_07281_),
    .B1(_07472_),
    .B2(_07473_),
    .C1(_07283_),
    .X(_07474_));
 sky130_fd_sc_hd__o21a_1 _12774_ (.A1(\core.csr.trapReturnVector[1] ),
    .A2(_07284_),
    .B1(_07474_),
    .X(_07475_));
 sky130_fd_sc_hd__a221o_1 _12775_ (.A1(\core.csr.traps.mtvec.csrReadData[1] ),
    .A2(_07231_),
    .B1(_07280_),
    .B2(\core.csr.traps.mscratch.currentValue[1] ),
    .C1(_07475_),
    .X(_07476_));
 sky130_fd_sc_hd__mux2_2 _12776_ (.A0(\core.csr.traps.mie.currentValue[1] ),
    .A1(_07476_),
    .S(_07219_),
    .X(_07477_));
 sky130_fd_sc_hd__a221o_4 _12777_ (.A1(\core.csr.mconfigptr.currentValue[1] ),
    .A2(_07285_),
    .B1(_07286_),
    .B2(net2),
    .C1(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__mux2_1 _12778_ (.A0(_07471_),
    .A1(_07478_),
    .S(_07278_),
    .X(_07479_));
 sky130_fd_sc_hd__a21o_1 _12779_ (.A1(net271),
    .A2(_07277_),
    .B1(_07479_),
    .X(_07480_));
 sky130_fd_sc_hd__mux2_1 _12780_ (.A0(_07480_),
    .A1(net255),
    .S(_07276_),
    .X(_07481_));
 sky130_fd_sc_hd__a221o_1 _12781_ (.A1(\core.csr.cycleTimer.currentValue[33] ),
    .A2(net716),
    .B1(_07470_),
    .B2(net979),
    .C1(_07481_),
    .X(_07482_));
 sky130_fd_sc_hd__mux2_2 _12782_ (.A0(\core.csr.cycleTimer.currentValue[1] ),
    .A1(_07482_),
    .S(net707),
    .X(_07483_));
 sky130_fd_sc_hd__a21oi_4 _12783_ (.A1(net979),
    .A2(_07468_),
    .B1(_07483_),
    .Y(_07484_));
 sky130_fd_sc_hd__o21ai_1 _12784_ (.A1(net1112),
    .A2(_07484_),
    .B1(_07467_),
    .Y(_07485_));
 sky130_fd_sc_hd__a21o_1 _12785_ (.A1(net1109),
    .A2(_07467_),
    .B1(net1104),
    .X(_07486_));
 sky130_fd_sc_hd__a21o_4 _12786_ (.A1(\core.pipe0_currentInstruction[1] ),
    .A2(\core.pipe0_currentInstruction[0] ),
    .B1(net1634),
    .X(_07487_));
 sky130_fd_sc_hd__nor2_2 _12787_ (.A(net461),
    .B(net1300),
    .Y(_07488_));
 sky130_fd_sc_hd__and2_1 _12788_ (.A(net461),
    .B(net1300),
    .X(_07489_));
 sky130_fd_sc_hd__nor2_1 _12789_ (.A(_07488_),
    .B(_07489_),
    .Y(_07490_));
 sky130_fd_sc_hd__inv_2 _12790_ (.A(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__a221o_1 _12791_ (.A1(net1151),
    .A2(net635),
    .B1(net1133),
    .B2(_07491_),
    .C1(net1266),
    .X(_07492_));
 sky130_fd_sc_hd__a31o_1 _12792_ (.A1(net1122),
    .A2(_07485_),
    .A3(_07486_),
    .B1(_07492_),
    .X(_07493_));
 sky130_fd_sc_hd__mux2_1 _12793_ (.A0(_07374_),
    .A1(_07396_),
    .S(net883),
    .X(_07494_));
 sky130_fd_sc_hd__mux2_1 _12794_ (.A0(_07395_),
    .A1(_07399_),
    .S(net883),
    .X(_07495_));
 sky130_fd_sc_hd__mux2_1 _12795_ (.A0(_07494_),
    .A1(_07495_),
    .S(net887),
    .X(_07496_));
 sky130_fd_sc_hd__mux2_2 _12796_ (.A0(_07388_),
    .A1(_07391_),
    .S(net885),
    .X(_07497_));
 sky130_fd_sc_hd__mux2_1 _12797_ (.A0(_07398_),
    .A1(_07389_),
    .S(net883),
    .X(_07498_));
 sky130_fd_sc_hd__mux2_1 _12798_ (.A0(_07497_),
    .A1(_07498_),
    .S(net744),
    .X(_07499_));
 sky130_fd_sc_hd__mux2_1 _12799_ (.A0(_07496_),
    .A1(_07499_),
    .S(net890),
    .X(_07500_));
 sky130_fd_sc_hd__mux2_1 _12800_ (.A0(_07425_),
    .A1(_07379_),
    .S(net882),
    .X(_07501_));
 sky130_fd_sc_hd__mux2_1 _12801_ (.A0(_07378_),
    .A1(_07383_),
    .S(net882),
    .X(_07502_));
 sky130_fd_sc_hd__mux2_1 _12802_ (.A0(_07501_),
    .A1(_07502_),
    .S(net886),
    .X(_07503_));
 sky130_fd_sc_hd__inv_2 _12803_ (.A(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__mux2_1 _12804_ (.A0(_07382_),
    .A1(_07371_),
    .S(net882),
    .X(_07505_));
 sky130_fd_sc_hd__mux2_1 _12805_ (.A0(_07370_),
    .A1(_07375_),
    .S(net881),
    .X(_07506_));
 sky130_fd_sc_hd__mux2_1 _12806_ (.A0(_07505_),
    .A1(_07506_),
    .S(net887),
    .X(_07507_));
 sky130_fd_sc_hd__mux2_1 _12807_ (.A0(_07504_),
    .A1(_07507_),
    .S(net890),
    .X(_07508_));
 sky130_fd_sc_hd__mux2_1 _12808_ (.A0(_07500_),
    .A1(_07508_),
    .S(net749),
    .X(_07509_));
 sky130_fd_sc_hd__mux2_1 _12809_ (.A0(_07410_),
    .A1(_07406_),
    .S(net884),
    .X(_07510_));
 sky130_fd_sc_hd__inv_2 _12810_ (.A(_07510_),
    .Y(_07511_));
 sky130_fd_sc_hd__mux2_1 _12811_ (.A0(_07449_),
    .A1(_07511_),
    .S(net888),
    .X(_07512_));
 sky130_fd_sc_hd__mux2_1 _12812_ (.A0(_07405_),
    .A1(_07414_),
    .S(net884),
    .X(_07513_));
 sky130_fd_sc_hd__mux2_1 _12813_ (.A0(_07413_),
    .A1(_07417_),
    .S(net884),
    .X(_07514_));
 sky130_fd_sc_hd__mux2_1 _12814_ (.A0(_07513_),
    .A1(_07514_),
    .S(net888),
    .X(_07515_));
 sky130_fd_sc_hd__inv_2 _12815_ (.A(_07515_),
    .Y(_07516_));
 sky130_fd_sc_hd__mux2_1 _12816_ (.A0(_07512_),
    .A1(_07516_),
    .S(net891),
    .X(_07517_));
 sky130_fd_sc_hd__inv_2 _12817_ (.A(_07517_),
    .Y(_07518_));
 sky130_fd_sc_hd__mux2_1 _12818_ (.A0(_07416_),
    .A1(_07432_),
    .S(net883),
    .X(_07519_));
 sky130_fd_sc_hd__mux2_1 _12819_ (.A0(_07430_),
    .A1(_07435_),
    .S(net881),
    .X(_07520_));
 sky130_fd_sc_hd__mux2_1 _12820_ (.A0(_07519_),
    .A1(_07520_),
    .S(net886),
    .X(_07521_));
 sky130_fd_sc_hd__nor2_1 _12821_ (.A(net881),
    .B(_07434_),
    .Y(_07522_));
 sky130_fd_sc_hd__a21oi_2 _12822_ (.A1(net881),
    .A2(_07423_),
    .B1(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__nand2_1 _12823_ (.A(net882),
    .B(_07426_),
    .Y(_07524_));
 sky130_fd_sc_hd__o21ai_1 _12824_ (.A1(net881),
    .A2(_07422_),
    .B1(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__mux2_1 _12825_ (.A0(_07523_),
    .A1(_07525_),
    .S(net886),
    .X(_07526_));
 sky130_fd_sc_hd__inv_2 _12826_ (.A(_07526_),
    .Y(_07527_));
 sky130_fd_sc_hd__mux2_1 _12827_ (.A0(_07521_),
    .A1(_07527_),
    .S(net890),
    .X(_07528_));
 sky130_fd_sc_hd__mux2_2 _12828_ (.A0(_07518_),
    .A1(_07528_),
    .S(net746),
    .X(_07529_));
 sky130_fd_sc_hd__mux2_4 _12829_ (.A0(_07509_),
    .A1(_07529_),
    .S(net755),
    .X(_07530_));
 sky130_fd_sc_hd__mux2_1 _12830_ (.A0(_07411_),
    .A1(_07445_),
    .S(net745),
    .X(_07531_));
 sky130_fd_sc_hd__o21ai_2 _12831_ (.A1(net895),
    .A2(_07531_),
    .B1(_07448_),
    .Y(_07532_));
 sky130_fd_sc_hd__a21boi_1 _12832_ (.A1(net747),
    .A2(_07532_),
    .B1_N(_07447_),
    .Y(_07533_));
 sky130_fd_sc_hd__inv_2 _12833_ (.A(_07533_),
    .Y(_07534_));
 sky130_fd_sc_hd__a21o_1 _12834_ (.A1(net753),
    .A2(_07534_),
    .B1(net632),
    .X(_07535_));
 sky130_fd_sc_hd__nor2_1 _12835_ (.A(net1211),
    .B(_07535_),
    .Y(_07536_));
 sky130_fd_sc_hd__nor2_8 _12836_ (.A(_04062_),
    .B(_06645_),
    .Y(_07537_));
 sky130_fd_sc_hd__or2_1 _12837_ (.A(_04062_),
    .B(_06645_),
    .X(_07538_));
 sky130_fd_sc_hd__mux2_1 _12838_ (.A0(_07537_),
    .A1(net1200),
    .S(_04970_),
    .X(_07539_));
 sky130_fd_sc_hd__o22a_1 _12839_ (.A1(net745),
    .A2(_04969_),
    .B1(net1205),
    .B2(_07539_),
    .X(_07540_));
 sky130_fd_sc_hd__a2111o_4 _12840_ (.A1(_07142_),
    .A2(_07530_),
    .B1(_07536_),
    .C1(_07540_),
    .D1(net1274),
    .X(_07541_));
 sky130_fd_sc_hd__a21o_1 _12841_ (.A1(net635),
    .A2(net1061),
    .B1(net1234),
    .X(_07542_));
 sky130_fd_sc_hd__or2_1 _12842_ (.A(_04972_),
    .B(_07305_),
    .X(_07543_));
 sky130_fd_sc_hd__a31o_2 _12843_ (.A1(_07306_),
    .A2(net1065),
    .A3(_07543_),
    .B1(_07542_),
    .X(_07544_));
 sky130_fd_sc_hd__a31o_1 _12844_ (.A1(_07147_),
    .A2(_07541_),
    .A3(_07544_),
    .B1(_07493_),
    .X(_07545_));
 sky130_fd_sc_hd__a32o_1 _12845_ (.A1(_04936_),
    .A2(net825),
    .A3(_07545_),
    .B1(net984),
    .B2(\core.pipe1_resultRegister[1] ),
    .X(_07546_));
 sky130_fd_sc_hd__and2_1 _12846_ (.A(net1821),
    .B(_07546_),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _12847_ (.A0(net1669),
    .A1(_04882_),
    .S(net1115),
    .X(_07547_));
 sky130_fd_sc_hd__a22o_1 _12848_ (.A1(\core.csr.cycleTimer.currentValue[2] ),
    .A2(net726),
    .B1(net722),
    .B2(\core.csr.cycleTimer.currentValue[34] ),
    .X(_07548_));
 sky130_fd_sc_hd__o31a_1 _12849_ (.A1(\core.csr.traps.mtvec.csrReadData[2] ),
    .A2(_07214_),
    .A3(_07230_),
    .B1(_07219_),
    .X(_07549_));
 sky130_fd_sc_hd__a22o_1 _12850_ (.A1(\core.csr.instretTimer.currentValue[2] ),
    .A2(net703),
    .B1(net699),
    .B2(\core.csr.instretTimer.currentValue[34] ),
    .X(_07550_));
 sky130_fd_sc_hd__and2_1 _12851_ (.A(net282),
    .B(_07171_),
    .X(_07551_));
 sky130_fd_sc_hd__mux2_1 _12852_ (.A0(\core.csr.traps.mip.csrReadData[2] ),
    .A1(\core.csr.traps.mtval.csrReadData[2] ),
    .S(net657),
    .X(_07552_));
 sky130_fd_sc_hd__a221o_1 _12853_ (.A1(\core.csr.traps.mcause.csrReadData[2] ),
    .A2(_07281_),
    .B1(_07472_),
    .B2(_07552_),
    .C1(_07283_),
    .X(_07553_));
 sky130_fd_sc_hd__o21ba_1 _12854_ (.A1(\core.csr.trapReturnVector[2] ),
    .A2(_07284_),
    .B1_N(_07280_),
    .X(_07554_));
 sky130_fd_sc_hd__a221o_1 _12855_ (.A1(\core.csr.traps.mscratch.currentValue[2] ),
    .A2(_07280_),
    .B1(_07553_),
    .B2(_07554_),
    .C1(_07231_),
    .X(_07555_));
 sky130_fd_sc_hd__a22o_1 _12856_ (.A1(\core.csr.traps.mie.currentValue[2] ),
    .A2(_07218_),
    .B1(_07549_),
    .B2(_07555_),
    .X(_07556_));
 sky130_fd_sc_hd__mux2_2 _12857_ (.A0(\core.csr.traps.machineInterruptEnable ),
    .A1(_07556_),
    .S(_07469_),
    .X(_07557_));
 sky130_fd_sc_hd__a221o_4 _12858_ (.A1(\core.csr.mconfigptr.currentValue[2] ),
    .A2(_07285_),
    .B1(_07286_),
    .B2(net3),
    .C1(_07557_),
    .X(_07558_));
 sky130_fd_sc_hd__mux2_1 _12859_ (.A0(_07551_),
    .A1(_07558_),
    .S(_07278_),
    .X(_07559_));
 sky130_fd_sc_hd__a21o_1 _12860_ (.A1(net272),
    .A2(_07277_),
    .B1(_07559_),
    .X(_07560_));
 sky130_fd_sc_hd__mux2_1 _12861_ (.A0(_07560_),
    .A1(net256),
    .S(_07276_),
    .X(_07561_));
 sky130_fd_sc_hd__a221o_1 _12862_ (.A1(\core.csr.cycleTimer.currentValue[34] ),
    .A2(net716),
    .B1(_07550_),
    .B2(net980),
    .C1(_07561_),
    .X(_07562_));
 sky130_fd_sc_hd__mux2_2 _12863_ (.A0(\core.csr.cycleTimer.currentValue[2] ),
    .A1(_07562_),
    .S(net707),
    .X(_07563_));
 sky130_fd_sc_hd__a21oi_4 _12864_ (.A1(net980),
    .A2(_07548_),
    .B1(_07563_),
    .Y(_07564_));
 sky130_fd_sc_hd__inv_2 _12865_ (.A(_07564_),
    .Y(_07565_));
 sky130_fd_sc_hd__o21ai_1 _12866_ (.A1(net1112),
    .A2(_07564_),
    .B1(_07547_),
    .Y(_07566_));
 sky130_fd_sc_hd__a21o_1 _12867_ (.A1(net1109),
    .A2(_07547_),
    .B1(net1104),
    .X(_07567_));
 sky130_fd_sc_hd__xnor2_2 _12868_ (.A(net472),
    .B(_07488_),
    .Y(_07568_));
 sky130_fd_sc_hd__inv_2 _12869_ (.A(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__a221o_1 _12870_ (.A1(net1151),
    .A2(_06713_),
    .B1(net1133),
    .B2(_07568_),
    .C1(net1266),
    .X(_07570_));
 sky130_fd_sc_hd__a31o_1 _12871_ (.A1(net1123),
    .A2(_07566_),
    .A3(_07567_),
    .B1(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__nand2_1 _12872_ (.A(net744),
    .B(_07384_),
    .Y(_07572_));
 sky130_fd_sc_hd__o21ai_1 _12873_ (.A1(net744),
    .A2(_07372_),
    .B1(_07572_),
    .Y(_07573_));
 sky130_fd_sc_hd__mux2_1 _12874_ (.A0(_07380_),
    .A1(_07427_),
    .S(net744),
    .X(_07574_));
 sky130_fd_sc_hd__mux2_1 _12875_ (.A0(_07573_),
    .A1(_07574_),
    .S(net893),
    .X(_07575_));
 sky130_fd_sc_hd__mux2_1 _12876_ (.A0(_07376_),
    .A1(_07397_),
    .S(net887),
    .X(_07576_));
 sky130_fd_sc_hd__inv_2 _12877_ (.A(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__mux2_1 _12878_ (.A0(_07390_),
    .A1(_07400_),
    .S(net745),
    .X(_07578_));
 sky130_fd_sc_hd__nor2_1 _12879_ (.A(net894),
    .B(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__a211o_1 _12880_ (.A1(net894),
    .A2(_07577_),
    .B1(_07579_),
    .C1(net749),
    .X(_07580_));
 sky130_fd_sc_hd__mux2_1 _12881_ (.A0(_07407_),
    .A1(_07415_),
    .S(net888),
    .X(_07581_));
 sky130_fd_sc_hd__mux2_1 _12882_ (.A0(_07531_),
    .A1(_07581_),
    .S(net892),
    .X(_07582_));
 sky130_fd_sc_hd__inv_2 _12883_ (.A(_07582_),
    .Y(_07583_));
 sky130_fd_sc_hd__mux2_1 _12884_ (.A0(_07424_),
    .A1(_07437_),
    .S(net744),
    .X(_07584_));
 sky130_fd_sc_hd__inv_2 _12885_ (.A(_07584_),
    .Y(_07585_));
 sky130_fd_sc_hd__mux2_1 _12886_ (.A0(_07418_),
    .A1(_07433_),
    .S(net887),
    .X(_07586_));
 sky130_fd_sc_hd__mux2_1 _12887_ (.A0(_07584_),
    .A1(_07586_),
    .S(net893),
    .X(_07587_));
 sky130_fd_sc_hd__inv_2 _12888_ (.A(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__mux2_1 _12889_ (.A0(_07583_),
    .A1(_07588_),
    .S(net748),
    .X(_07589_));
 sky130_fd_sc_hd__o211a_1 _12890_ (.A1(net746),
    .A2(_07575_),
    .B1(_07580_),
    .C1(net752),
    .X(_07590_));
 sky130_fd_sc_hd__a21o_1 _12891_ (.A1(net756),
    .A2(_07589_),
    .B1(_07590_),
    .X(_07591_));
 sky130_fd_sc_hd__o21ai_1 _12892_ (.A1(_04885_),
    .A2(net1198),
    .B1(net1204),
    .Y(_07592_));
 sky130_fd_sc_hd__a22o_1 _12893_ (.A1(_04885_),
    .A2(net1202),
    .B1(_07592_),
    .B2(_04886_),
    .X(_07593_));
 sky130_fd_sc_hd__a21bo_1 _12894_ (.A1(net892),
    .A2(_07512_),
    .B1_N(_07448_),
    .X(_07594_));
 sky130_fd_sc_hd__inv_2 _12895_ (.A(_07594_),
    .Y(_07595_));
 sky130_fd_sc_hd__o21ai_1 _12896_ (.A1(net751),
    .A2(_07595_),
    .B1(_07447_),
    .Y(_07596_));
 sky130_fd_sc_hd__a21o_1 _12897_ (.A1(net752),
    .A2(_07596_),
    .B1(net631),
    .X(_07597_));
 sky130_fd_sc_hd__o22a_2 _12898_ (.A1(net1215),
    .A2(_07591_),
    .B1(_07597_),
    .B2(net1207),
    .X(_07598_));
 sky130_fd_sc_hd__or3b_2 _12899_ (.A(net1274),
    .B(_07593_),
    .C_N(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__xor2_2 _12900_ (.A(_06712_),
    .B(_07307_),
    .X(_07600_));
 sky130_fd_sc_hd__and2_1 _12901_ (.A(net1065),
    .B(_07600_),
    .X(_07601_));
 sky130_fd_sc_hd__a211o_1 _12902_ (.A1(_06713_),
    .A2(net1061),
    .B1(_07601_),
    .C1(net1234),
    .X(_07602_));
 sky130_fd_sc_hd__a31o_1 _12903_ (.A1(_07147_),
    .A2(_07599_),
    .A3(_07602_),
    .B1(_07571_),
    .X(_07603_));
 sky130_fd_sc_hd__a32o_1 _12904_ (.A1(_04854_),
    .A2(net825),
    .A3(_07603_),
    .B1(net984),
    .B2(\core.pipe1_resultRegister[2] ),
    .X(_07604_));
 sky130_fd_sc_hd__and2_1 _12905_ (.A(net1821),
    .B(_07604_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _12906_ (.A0(_03839_),
    .A1(_04801_),
    .S(net1114),
    .X(_07605_));
 sky130_fd_sc_hd__a22o_1 _12907_ (.A1(\core.csr.cycleTimer.currentValue[3] ),
    .A2(net726),
    .B1(net722),
    .B2(\core.csr.cycleTimer.currentValue[35] ),
    .X(_07606_));
 sky130_fd_sc_hd__a22o_1 _12908_ (.A1(\core.csr.instretTimer.currentValue[3] ),
    .A2(net703),
    .B1(net699),
    .B2(\core.csr.instretTimer.currentValue[35] ),
    .X(_07607_));
 sky130_fd_sc_hd__a21o_1 _12909_ (.A1(net283),
    .A2(_07171_),
    .B1(_07278_),
    .X(_07608_));
 sky130_fd_sc_hd__mux2_1 _12910_ (.A0(\core.csr.traps.mip.csrReadData[3] ),
    .A1(\core.csr.traps.mtval.csrReadData[3] ),
    .S(net656),
    .X(_07609_));
 sky130_fd_sc_hd__a221o_1 _12911_ (.A1(\core.csr.traps.mcause.csrReadData[3] ),
    .A2(_07281_),
    .B1(_07472_),
    .B2(_07609_),
    .C1(_07283_),
    .X(_07610_));
 sky130_fd_sc_hd__o21a_2 _12912_ (.A1(\core.csr.trapReturnVector[3] ),
    .A2(_07284_),
    .B1(_07610_),
    .X(_07611_));
 sky130_fd_sc_hd__a221o_1 _12913_ (.A1(\core.csr.traps.mtvec.csrReadData[3] ),
    .A2(_07231_),
    .B1(_07280_),
    .B2(\core.csr.traps.mscratch.currentValue[3] ),
    .C1(_07611_),
    .X(_07612_));
 sky130_fd_sc_hd__mux2_2 _12914_ (.A0(\core.csr.traps.mie.currentValue[3] ),
    .A1(_07612_),
    .S(_07219_),
    .X(_07613_));
 sky130_fd_sc_hd__a2bb2o_1 _12915_ (.A1_N(_07222_),
    .A2_N(_07275_),
    .B1(_07286_),
    .B2(net4),
    .X(_07614_));
 sky130_fd_sc_hd__a211o_4 _12916_ (.A1(\core.csr.mconfigptr.currentValue[3] ),
    .A2(_07285_),
    .B1(_07613_),
    .C1(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__a22o_1 _12917_ (.A1(net273),
    .A2(_07277_),
    .B1(_07608_),
    .B2(_07615_),
    .X(_07616_));
 sky130_fd_sc_hd__mux2_1 _12918_ (.A0(_07616_),
    .A1(net257),
    .S(_07276_),
    .X(_07617_));
 sky130_fd_sc_hd__a221o_1 _12919_ (.A1(\core.csr.cycleTimer.currentValue[35] ),
    .A2(net716),
    .B1(_07607_),
    .B2(net980),
    .C1(_07617_),
    .X(_07618_));
 sky130_fd_sc_hd__mux2_2 _12920_ (.A0(\core.csr.cycleTimer.currentValue[3] ),
    .A1(_07618_),
    .S(net708),
    .X(_07619_));
 sky130_fd_sc_hd__a21oi_4 _12921_ (.A1(net980),
    .A2(_07606_),
    .B1(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__inv_2 _12922_ (.A(_07620_),
    .Y(_07621_));
 sky130_fd_sc_hd__o21ai_1 _12923_ (.A1(net1112),
    .A2(_07620_),
    .B1(_07605_),
    .Y(_07622_));
 sky130_fd_sc_hd__a21o_1 _12924_ (.A1(net1109),
    .A2(_07605_),
    .B1(net1104),
    .X(_07623_));
 sky130_fd_sc_hd__o211a_4 _12925_ (.A1(net461),
    .A2(net1300),
    .B1(net475),
    .C1(net472),
    .X(_07624_));
 sky130_fd_sc_hd__o21ba_1 _12926_ (.A1(_03827_),
    .A2(_07488_),
    .B1_N(net475),
    .X(_07625_));
 sky130_fd_sc_hd__nor2_1 _12927_ (.A(_07624_),
    .B(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__a221o_1 _12928_ (.A1(net1151),
    .A2(_06715_),
    .B1(net1133),
    .B2(_07626_),
    .C1(net1266),
    .X(_07627_));
 sky130_fd_sc_hd__a31o_1 _12929_ (.A1(net1123),
    .A2(_07622_),
    .A3(_07623_),
    .B1(_07627_),
    .X(_07628_));
 sky130_fd_sc_hd__mux2_1 _12930_ (.A0(_07510_),
    .A1(_07513_),
    .S(net888),
    .X(_07629_));
 sky130_fd_sc_hd__mux2_2 _12931_ (.A0(_07451_),
    .A1(_07629_),
    .S(net892),
    .X(_07630_));
 sky130_fd_sc_hd__or2_1 _12932_ (.A(net747),
    .B(_07630_),
    .X(_07631_));
 sky130_fd_sc_hd__nor2_1 _12933_ (.A(net886),
    .B(_07520_),
    .Y(_07632_));
 sky130_fd_sc_hd__a21oi_2 _12934_ (.A1(net886),
    .A2(_07523_),
    .B1(_07632_),
    .Y(_07633_));
 sky130_fd_sc_hd__mux2_1 _12935_ (.A0(_07514_),
    .A1(_07519_),
    .S(net888),
    .X(_07634_));
 sky130_fd_sc_hd__mux2_1 _12936_ (.A0(_07633_),
    .A1(_07634_),
    .S(net895),
    .X(_07635_));
 sky130_fd_sc_hd__o21ai_1 _12937_ (.A1(net751),
    .A2(_07635_),
    .B1(_07631_),
    .Y(_07636_));
 sky130_fd_sc_hd__nand2_1 _12938_ (.A(net744),
    .B(_07502_),
    .Y(_07637_));
 sky130_fd_sc_hd__o21ai_1 _12939_ (.A1(net744),
    .A2(_07505_),
    .B1(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__mux2_1 _12940_ (.A0(_07501_),
    .A1(_07525_),
    .S(net744),
    .X(_07639_));
 sky130_fd_sc_hd__mux2_2 _12941_ (.A0(_07638_),
    .A1(_07639_),
    .S(net893),
    .X(_07640_));
 sky130_fd_sc_hd__mux2_1 _12942_ (.A0(_07494_),
    .A1(_07506_),
    .S(net744),
    .X(_07641_));
 sky130_fd_sc_hd__mux2_1 _12943_ (.A0(_07495_),
    .A1(_07498_),
    .S(net887),
    .X(_07642_));
 sky130_fd_sc_hd__mux2_1 _12944_ (.A0(_07641_),
    .A1(_07642_),
    .S(net890),
    .X(_07643_));
 sky130_fd_sc_hd__nand2_1 _12945_ (.A(net746),
    .B(_07643_),
    .Y(_07644_));
 sky130_fd_sc_hd__o211a_1 _12946_ (.A1(net746),
    .A2(_07640_),
    .B1(_07644_),
    .C1(net752),
    .X(_07645_));
 sky130_fd_sc_hd__a21o_2 _12947_ (.A1(net755),
    .A2(_07636_),
    .B1(_07645_),
    .X(_07646_));
 sky130_fd_sc_hd__o21a_1 _12948_ (.A1(_04806_),
    .A2(net1198),
    .B1(net1204),
    .X(_07647_));
 sky130_fd_sc_hd__o2bb2a_2 _12949_ (.A1_N(_04806_),
    .A2_N(net1202),
    .B1(_07647_),
    .B2(_04804_),
    .X(_07648_));
 sky130_fd_sc_hd__o21ai_1 _12950_ (.A1(net895),
    .A2(_07412_),
    .B1(_07448_),
    .Y(_07649_));
 sky130_fd_sc_hd__a21boi_1 _12951_ (.A1(net747),
    .A2(_07649_),
    .B1_N(_07447_),
    .Y(_07650_));
 sky130_fd_sc_hd__inv_2 _12952_ (.A(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__a21o_1 _12953_ (.A1(net753),
    .A2(_07651_),
    .B1(net631),
    .X(_07652_));
 sky130_fd_sc_hd__o211a_1 _12954_ (.A1(net1210),
    .A2(_07652_),
    .B1(_07648_),
    .C1(_07000_),
    .X(_07653_));
 sky130_fd_sc_hd__o21ai_4 _12955_ (.A1(net1217),
    .A2(_07646_),
    .B1(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__and2_1 _12956_ (.A(_06715_),
    .B(net1061),
    .X(_07655_));
 sky130_fd_sc_hd__xor2_4 _12957_ (.A(_06714_),
    .B(_07308_),
    .X(_07656_));
 sky130_fd_sc_hd__a211o_1 _12958_ (.A1(net1066),
    .A2(_07656_),
    .B1(_07655_),
    .C1(net1235),
    .X(_07657_));
 sky130_fd_sc_hd__a31o_1 _12959_ (.A1(_07147_),
    .A2(_07654_),
    .A3(_07657_),
    .B1(_07628_),
    .X(_07658_));
 sky130_fd_sc_hd__a32o_1 _12960_ (.A1(_04768_),
    .A2(net825),
    .A3(_07658_),
    .B1(net984),
    .B2(\core.pipe1_resultRegister[3] ),
    .X(_07659_));
 sky130_fd_sc_hd__and2_1 _12961_ (.A(net1821),
    .B(_07659_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _12962_ (.A0(net1783),
    .A1(_04719_),
    .S(net1114),
    .X(_07660_));
 sky130_fd_sc_hd__a22o_1 _12963_ (.A1(\core.csr.cycleTimer.currentValue[4] ),
    .A2(net727),
    .B1(net723),
    .B2(\core.csr.cycleTimer.currentValue[36] ),
    .X(_07661_));
 sky130_fd_sc_hd__a21o_1 _12964_ (.A1(net274),
    .A2(_07238_),
    .B1(_07207_),
    .X(_07662_));
 sky130_fd_sc_hd__a22o_1 _12965_ (.A1(\core.csr.instretTimer.currentValue[4] ),
    .A2(net703),
    .B1(net699),
    .B2(\core.csr.instretTimer.currentValue[36] ),
    .X(_07663_));
 sky130_fd_sc_hd__or2_1 _12966_ (.A(\core.csr.cycleTimer.currentValue[4] ),
    .B(net707),
    .X(_07664_));
 sky130_fd_sc_hd__a21o_1 _12967_ (.A1(\core.csr.mconfigptr.currentValue[4] ),
    .A2(net719),
    .B1(_07253_),
    .X(_07665_));
 sky130_fd_sc_hd__or2_1 _12968_ (.A(\core.csr.traps.mip.csrReadData[4] ),
    .B(net656),
    .X(_07666_));
 sky130_fd_sc_hd__o211a_1 _12969_ (.A1(\core.csr.traps.mtval.csrReadData[4] ),
    .A2(net663),
    .B1(net660),
    .C1(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__a21o_1 _12970_ (.A1(\core.csr.traps.mcause.csrReadData[4] ),
    .A2(net666),
    .B1(net690),
    .X(_07668_));
 sky130_fd_sc_hd__o221a_1 _12971_ (.A1(\core.csr.trapReturnVector[4] ),
    .A2(net687),
    .B1(_07667_),
    .B2(_07668_),
    .C1(net693),
    .X(_07669_));
 sky130_fd_sc_hd__a221o_1 _12972_ (.A1(\core.csr.traps.mscratch.currentValue[4] ),
    .A2(net696),
    .B1(net678),
    .B2(\core.csr.traps.mtvec.csrReadData[4] ),
    .C1(net684),
    .X(_07670_));
 sky130_fd_sc_hd__o221a_4 _12973_ (.A1(\core.csr.traps.mie.currentValue[4] ),
    .A2(net681),
    .B1(_07669_),
    .B2(_07670_),
    .C1(net609),
    .X(_07671_));
 sky130_fd_sc_hd__o221a_2 _12974_ (.A1(net5),
    .A2(_07254_),
    .B1(_07665_),
    .B2(_07671_),
    .C1(_07239_),
    .X(_07672_));
 sky130_fd_sc_hd__o221a_1 _12975_ (.A1(net258),
    .A2(_07208_),
    .B1(_07662_),
    .B2(_07672_),
    .C1(_07212_),
    .X(_07673_));
 sky130_fd_sc_hd__a221o_1 _12976_ (.A1(\core.csr.cycleTimer.currentValue[36] ),
    .A2(net715),
    .B1(_07663_),
    .B2(net980),
    .C1(net711),
    .X(_07674_));
 sky130_fd_sc_hd__or2_1 _12977_ (.A(_07673_),
    .B(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__a22o_4 _12978_ (.A1(net980),
    .A2(_07661_),
    .B1(_07664_),
    .B2(_07675_),
    .X(_07676_));
 sky130_fd_sc_hd__a21o_1 _12979_ (.A1(net1111),
    .A2(_07676_),
    .B1(_07660_),
    .X(_07677_));
 sky130_fd_sc_hd__o21ai_1 _12980_ (.A1(net1108),
    .A2(_07660_),
    .B1(net1107),
    .Y(_07678_));
 sky130_fd_sc_hd__xnor2_4 _12981_ (.A(net1748),
    .B(_07624_),
    .Y(_07679_));
 sky130_fd_sc_hd__nor2_1 _12982_ (.A(net1136),
    .B(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__a211o_1 _12983_ (.A1(net1151),
    .A2(_06716_),
    .B1(_07680_),
    .C1(net1267),
    .X(_07681_));
 sky130_fd_sc_hd__a31o_1 _12984_ (.A1(net1122),
    .A2(_07677_),
    .A3(_07678_),
    .B1(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__xnor2_1 _12985_ (.A(_04724_),
    .B(_07309_),
    .Y(_07683_));
 sky130_fd_sc_hd__o21a_1 _12986_ (.A1(_06716_),
    .A2(net1065),
    .B1(net1275),
    .X(_07684_));
 sky130_fd_sc_hd__o21ai_1 _12987_ (.A1(net1061),
    .A2(_07683_),
    .B1(_07684_),
    .Y(_07685_));
 sky130_fd_sc_hd__or2_2 _12988_ (.A(net893),
    .B(_07438_),
    .X(_07686_));
 sky130_fd_sc_hd__o21ai_2 _12989_ (.A1(net891),
    .A2(_07419_),
    .B1(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__or2_1 _12990_ (.A(net747),
    .B(_07649_),
    .X(_07688_));
 sky130_fd_sc_hd__o21ai_1 _12991_ (.A1(net751),
    .A2(_07687_),
    .B1(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__inv_2 _12992_ (.A(_07689_),
    .Y(_07690_));
 sky130_fd_sc_hd__mux2_2 _12993_ (.A0(_07386_),
    .A1(_07429_),
    .S(net893),
    .X(_07691_));
 sky130_fd_sc_hd__inv_2 _12994_ (.A(_07691_),
    .Y(_07692_));
 sky130_fd_sc_hd__mux2_1 _12995_ (.A0(_07377_),
    .A1(_07401_),
    .S(net890),
    .X(_07693_));
 sky130_fd_sc_hd__mux2_1 _12996_ (.A0(_07691_),
    .A1(_07693_),
    .S(net746),
    .X(_07694_));
 sky130_fd_sc_hd__inv_2 _12997_ (.A(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__mux2_2 _12998_ (.A0(_07690_),
    .A1(_07695_),
    .S(net753),
    .X(_07696_));
 sky130_fd_sc_hd__mux2_2 _12999_ (.A0(net1202),
    .A1(_07537_),
    .S(_04721_),
    .X(_07697_));
 sky130_fd_sc_hd__o21ai_4 _13000_ (.A1(net1205),
    .A2(_07697_),
    .B1(_04723_),
    .Y(_07698_));
 sky130_fd_sc_hd__o21ai_4 _13001_ (.A1(net751),
    .A2(_07630_),
    .B1(_07447_),
    .Y(_07699_));
 sky130_fd_sc_hd__a21o_1 _13002_ (.A1(net753),
    .A2(_07699_),
    .B1(net632),
    .X(_07700_));
 sky130_fd_sc_hd__o221a_4 _13003_ (.A1(net1216),
    .A2(_07696_),
    .B1(_07700_),
    .B2(net1210),
    .C1(_07698_),
    .X(_07701_));
 sky130_fd_sc_hd__a21oi_2 _13004_ (.A1(_07685_),
    .A2(_07701_),
    .B1(_07146_),
    .Y(_07702_));
 sky130_fd_sc_hd__o221a_1 _13005_ (.A1(net1748),
    .A2(net1260),
    .B1(_07682_),
    .B2(_07702_),
    .C1(net825),
    .X(_07703_));
 sky130_fd_sc_hd__a21oi_1 _13006_ (.A1(\core.pipe1_resultRegister[4] ),
    .A2(net985),
    .B1(_07703_),
    .Y(_07704_));
 sky130_fd_sc_hd__nor2_1 _13007_ (.A(net1906),
    .B(_07704_),
    .Y(_00166_));
 sky130_fd_sc_hd__nor2_1 _13008_ (.A(_04597_),
    .B(net1117),
    .Y(_07705_));
 sky130_fd_sc_hd__a22o_1 _13009_ (.A1(\core.csr.cycleTimer.currentValue[5] ),
    .A2(net727),
    .B1(net723),
    .B2(\core.csr.cycleTimer.currentValue[37] ),
    .X(_07706_));
 sky130_fd_sc_hd__a21o_1 _13010_ (.A1(net275),
    .A2(_07238_),
    .B1(_07207_),
    .X(_07707_));
 sky130_fd_sc_hd__a22o_1 _13011_ (.A1(\core.csr.instretTimer.currentValue[5] ),
    .A2(net703),
    .B1(net699),
    .B2(\core.csr.instretTimer.currentValue[37] ),
    .X(_07708_));
 sky130_fd_sc_hd__or2_1 _13012_ (.A(\core.csr.cycleTimer.currentValue[5] ),
    .B(net707),
    .X(_07709_));
 sky130_fd_sc_hd__a21o_1 _13013_ (.A1(\core.csr.mconfigptr.currentValue[5] ),
    .A2(net719),
    .B1(_07253_),
    .X(_07710_));
 sky130_fd_sc_hd__or2_1 _13014_ (.A(\core.csr.traps.mip.csrReadData[5] ),
    .B(net656),
    .X(_07711_));
 sky130_fd_sc_hd__o211a_1 _13015_ (.A1(\core.csr.traps.mtval.csrReadData[5] ),
    .A2(net663),
    .B1(net660),
    .C1(_07711_),
    .X(_07712_));
 sky130_fd_sc_hd__a21o_1 _13016_ (.A1(\core.csr.traps.mcause.csrReadData[5] ),
    .A2(net666),
    .B1(net690),
    .X(_07713_));
 sky130_fd_sc_hd__o221a_1 _13017_ (.A1(\core.csr.trapReturnVector[5] ),
    .A2(net687),
    .B1(_07712_),
    .B2(_07713_),
    .C1(net693),
    .X(_07714_));
 sky130_fd_sc_hd__a221o_1 _13018_ (.A1(\core.csr.traps.mscratch.currentValue[5] ),
    .A2(net696),
    .B1(net678),
    .B2(\core.csr.traps.mtvec.csrReadData[5] ),
    .C1(net684),
    .X(_07715_));
 sky130_fd_sc_hd__o221a_4 _13019_ (.A1(\core.csr.traps.mie.currentValue[5] ),
    .A2(net681),
    .B1(_07714_),
    .B2(_07715_),
    .C1(net609),
    .X(_07716_));
 sky130_fd_sc_hd__o221a_2 _13020_ (.A1(net6),
    .A2(_07254_),
    .B1(_07710_),
    .B2(_07716_),
    .C1(_07239_),
    .X(_07717_));
 sky130_fd_sc_hd__o221a_1 _13021_ (.A1(net259),
    .A2(_07208_),
    .B1(_07707_),
    .B2(_07717_),
    .C1(_07212_),
    .X(_07718_));
 sky130_fd_sc_hd__a221o_1 _13022_ (.A1(\core.csr.cycleTimer.currentValue[37] ),
    .A2(net715),
    .B1(_07708_),
    .B2(net980),
    .C1(net711),
    .X(_07719_));
 sky130_fd_sc_hd__or2_1 _13023_ (.A(_07718_),
    .B(_07719_),
    .X(_07720_));
 sky130_fd_sc_hd__a22o_4 _13024_ (.A1(net980),
    .A2(_07706_),
    .B1(_07709_),
    .B2(_07720_),
    .X(_07721_));
 sky130_fd_sc_hd__a21o_1 _13025_ (.A1(net1111),
    .A2(_07721_),
    .B1(_07705_),
    .X(_07722_));
 sky130_fd_sc_hd__o21ai_1 _13026_ (.A1(net1108),
    .A2(_07705_),
    .B1(net1107),
    .Y(_07723_));
 sky130_fd_sc_hd__and3_1 _13027_ (.A(net1122),
    .B(_07722_),
    .C(_07723_),
    .X(_07724_));
 sky130_fd_sc_hd__and3_1 _13028_ (.A(net477),
    .B(net1748),
    .C(_07624_),
    .X(_07725_));
 sky130_fd_sc_hd__a21oi_1 _13029_ (.A1(net1748),
    .A2(_07624_),
    .B1(net477),
    .Y(_07726_));
 sky130_fd_sc_hd__nor2_1 _13030_ (.A(_07725_),
    .B(_07726_),
    .Y(_07727_));
 sky130_fd_sc_hd__a221o_1 _13031_ (.A1(net1152),
    .A2(_06718_),
    .B1(net1133),
    .B2(_07727_),
    .C1(net1267),
    .X(_07728_));
 sky130_fd_sc_hd__nor2_1 _13032_ (.A(_04636_),
    .B(_07312_),
    .Y(_07729_));
 sky130_fd_sc_hd__nand2_1 _13033_ (.A(_04636_),
    .B(_07312_),
    .Y(_07730_));
 sky130_fd_sc_hd__and2b_1 _13034_ (.A_N(_07729_),
    .B(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__nor2_1 _13035_ (.A(net1061),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__a211o_1 _13036_ (.A1(_06717_),
    .A2(net1061),
    .B1(_07732_),
    .C1(net1235),
    .X(_07733_));
 sky130_fd_sc_hd__mux2_1 _13037_ (.A0(_07503_),
    .A1(_07526_),
    .S(net893),
    .X(_07734_));
 sky130_fd_sc_hd__nand2_1 _13038_ (.A(net749),
    .B(_07734_),
    .Y(_07735_));
 sky130_fd_sc_hd__mux2_1 _13039_ (.A0(_07496_),
    .A1(_07507_),
    .S(net894),
    .X(_07736_));
 sky130_fd_sc_hd__o211a_1 _13040_ (.A1(net749),
    .A2(_07736_),
    .B1(_07735_),
    .C1(net752),
    .X(_07737_));
 sky130_fd_sc_hd__mux2_1 _13041_ (.A0(_07515_),
    .A1(_07521_),
    .S(net891),
    .X(_07738_));
 sky130_fd_sc_hd__mux2_1 _13042_ (.A0(_07595_),
    .A1(_07738_),
    .S(net747),
    .X(_07739_));
 sky130_fd_sc_hd__a21oi_2 _13043_ (.A1(net755),
    .A2(_07739_),
    .B1(_07737_),
    .Y(_07740_));
 sky130_fd_sc_hd__mux2_1 _13044_ (.A0(net1199),
    .A1(_07458_),
    .S(_04633_),
    .X(_07741_));
 sky130_fd_sc_hd__a21o_2 _13045_ (.A1(net1204),
    .A2(_07741_),
    .B1(_04634_),
    .X(_07742_));
 sky130_fd_sc_hd__o21a_1 _13046_ (.A1(net751),
    .A2(_07582_),
    .B1(_07447_),
    .X(_07743_));
 sky130_fd_sc_hd__inv_2 _13047_ (.A(_07743_),
    .Y(_07744_));
 sky130_fd_sc_hd__a21o_1 _13048_ (.A1(net754),
    .A2(_07744_),
    .B1(net631),
    .X(_07745_));
 sky130_fd_sc_hd__o221a_4 _13049_ (.A1(net1216),
    .A2(_07740_),
    .B1(_07745_),
    .B2(net1208),
    .C1(_07742_),
    .X(_07746_));
 sky130_fd_sc_hd__a21oi_1 _13050_ (.A1(_07733_),
    .A2(_07746_),
    .B1(_07146_),
    .Y(_07747_));
 sky130_fd_sc_hd__or3_1 _13051_ (.A(_07724_),
    .B(_07728_),
    .C(_07747_),
    .X(_07748_));
 sky130_fd_sc_hd__a32o_1 _13052_ (.A1(_04550_),
    .A2(net825),
    .A3(_07748_),
    .B1(net984),
    .B2(\core.pipe1_resultRegister[5] ),
    .X(_07749_));
 sky130_fd_sc_hd__and2_1 _13053_ (.A(net1821),
    .B(_07749_),
    .X(_00167_));
 sky130_fd_sc_hd__and2_1 _13054_ (.A(net478),
    .B(_07725_),
    .X(_07750_));
 sky130_fd_sc_hd__nor2_1 _13055_ (.A(net478),
    .B(_07725_),
    .Y(_07751_));
 sky130_fd_sc_hd__or2_2 _13056_ (.A(_07750_),
    .B(_07751_),
    .X(_07752_));
 sky130_fd_sc_hd__o21ai_1 _13057_ (.A1(net1136),
    .A2(_07752_),
    .B1(net1262),
    .Y(_07753_));
 sky130_fd_sc_hd__or2_1 _13058_ (.A(_04512_),
    .B(net1117),
    .X(_07754_));
 sky130_fd_sc_hd__a22o_1 _13059_ (.A1(\core.csr.cycleTimer.currentValue[6] ),
    .A2(net727),
    .B1(net723),
    .B2(\core.csr.cycleTimer.currentValue[38] ),
    .X(_07755_));
 sky130_fd_sc_hd__a21o_1 _13060_ (.A1(net276),
    .A2(_07238_),
    .B1(_07207_),
    .X(_07756_));
 sky130_fd_sc_hd__a22o_1 _13061_ (.A1(\core.csr.instretTimer.currentValue[6] ),
    .A2(net703),
    .B1(net699),
    .B2(\core.csr.instretTimer.currentValue[38] ),
    .X(_07757_));
 sky130_fd_sc_hd__a21oi_1 _13062_ (.A1(_03810_),
    .A2(net678),
    .B1(net684),
    .Y(_07758_));
 sky130_fd_sc_hd__o21a_1 _13063_ (.A1(\core.csr.trapReturnVector[6] ),
    .A2(net687),
    .B1(net693),
    .X(_07759_));
 sky130_fd_sc_hd__or2_1 _13064_ (.A(\core.csr.traps.mtval.csrReadData[6] ),
    .B(net663),
    .X(_07760_));
 sky130_fd_sc_hd__o21a_1 _13065_ (.A1(\core.csr.traps.mip.csrReadData[6] ),
    .A2(net657),
    .B1(net660),
    .X(_07761_));
 sky130_fd_sc_hd__a221o_1 _13066_ (.A1(\core.csr.traps.mcause.csrReadData[6] ),
    .A2(net666),
    .B1(_07760_),
    .B2(_07761_),
    .C1(net690),
    .X(_07762_));
 sky130_fd_sc_hd__a221o_1 _13067_ (.A1(\core.csr.traps.mscratch.currentValue[6] ),
    .A2(net696),
    .B1(_07759_),
    .B2(_07762_),
    .C1(net678),
    .X(_07763_));
 sky130_fd_sc_hd__a221o_2 _13068_ (.A1(\core.csr.traps.mie.currentValue[6] ),
    .A2(net684),
    .B1(_07758_),
    .B2(_07763_),
    .C1(_07269_),
    .X(_07764_));
 sky130_fd_sc_hd__o32a_2 _13069_ (.A1(net678),
    .A2(net660),
    .A3(_07272_),
    .B1(_07270_),
    .B2(\core.csr.traps.machinePreviousInterruptEnable ),
    .X(_07765_));
 sky130_fd_sc_hd__a221o_2 _13070_ (.A1(\core.csr.mconfigptr.currentValue[6] ),
    .A2(net717),
    .B1(_07764_),
    .B2(_07765_),
    .C1(_07253_),
    .X(_07766_));
 sky130_fd_sc_hd__o211a_2 _13071_ (.A1(net7),
    .A2(_07254_),
    .B1(_07766_),
    .C1(_07239_),
    .X(_07767_));
 sky130_fd_sc_hd__o221a_1 _13072_ (.A1(net260),
    .A2(_07208_),
    .B1(_07756_),
    .B2(_07767_),
    .C1(_07212_),
    .X(_07768_));
 sky130_fd_sc_hd__a221o_1 _13073_ (.A1(\core.csr.cycleTimer.currentValue[38] ),
    .A2(net715),
    .B1(_07757_),
    .B2(net980),
    .C1(net711),
    .X(_07769_));
 sky130_fd_sc_hd__o221a_2 _13074_ (.A1(\core.csr.cycleTimer.currentValue[6] ),
    .A2(net708),
    .B1(_07768_),
    .B2(_07769_),
    .C1(_07250_),
    .X(_07770_));
 sky130_fd_sc_hd__a21oi_4 _13075_ (.A1(net978),
    .A2(_07755_),
    .B1(_07770_),
    .Y(_07771_));
 sky130_fd_sc_hd__inv_2 _13076_ (.A(_07771_),
    .Y(_07772_));
 sky130_fd_sc_hd__o21ai_1 _13077_ (.A1(net1112),
    .A2(_07771_),
    .B1(_07754_),
    .Y(_07773_));
 sky130_fd_sc_hd__a21o_1 _13078_ (.A1(net1109),
    .A2(_07754_),
    .B1(net1105),
    .X(_07774_));
 sky130_fd_sc_hd__and3_1 _13079_ (.A(net1123),
    .B(_07773_),
    .C(_07774_),
    .X(_07775_));
 sky130_fd_sc_hd__a211o_1 _13080_ (.A1(net1152),
    .A2(_06720_),
    .B1(_07753_),
    .C1(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__and2_1 _13081_ (.A(_06720_),
    .B(net1061),
    .X(_07777_));
 sky130_fd_sc_hd__a21o_1 _13082_ (.A1(_07316_),
    .A2(_07730_),
    .B1(_06719_),
    .X(_07778_));
 sky130_fd_sc_hd__nand3_1 _13083_ (.A(_06719_),
    .B(_07316_),
    .C(_07730_),
    .Y(_07779_));
 sky130_fd_sc_hd__and2_1 _13084_ (.A(_07778_),
    .B(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__a211o_1 _13085_ (.A1(net1065),
    .A2(_07780_),
    .B1(_07777_),
    .C1(net1235),
    .X(_07781_));
 sky130_fd_sc_hd__mux2_1 _13086_ (.A0(_07574_),
    .A1(_07585_),
    .S(net893),
    .X(_07782_));
 sky130_fd_sc_hd__mux2_1 _13087_ (.A0(_07573_),
    .A1(_07577_),
    .S(net890),
    .X(_07783_));
 sky130_fd_sc_hd__mux2_1 _13088_ (.A0(_07782_),
    .A1(_07783_),
    .S(net746),
    .X(_07784_));
 sky130_fd_sc_hd__or2_1 _13089_ (.A(net893),
    .B(_07586_),
    .X(_07785_));
 sky130_fd_sc_hd__o21ai_1 _13090_ (.A1(net891),
    .A2(_07581_),
    .B1(_07785_),
    .Y(_07786_));
 sky130_fd_sc_hd__mux2_1 _13091_ (.A0(_07532_),
    .A1(_07786_),
    .S(net747),
    .X(_07787_));
 sky130_fd_sc_hd__mux2_2 _13092_ (.A0(_07784_),
    .A1(_07787_),
    .S(net755),
    .X(_07788_));
 sky130_fd_sc_hd__o21ai_1 _13093_ (.A1(net750),
    .A2(_07518_),
    .B1(_07447_),
    .Y(_07789_));
 sky130_fd_sc_hd__a21o_1 _13094_ (.A1(net752),
    .A2(_07789_),
    .B1(net631),
    .X(_07790_));
 sky130_fd_sc_hd__a221oi_4 _13095_ (.A1(_04548_),
    .A2(net1200),
    .B1(_07537_),
    .B2(_06719_),
    .C1(net1275),
    .Y(_07791_));
 sky130_fd_sc_hd__o221a_4 _13096_ (.A1(net1215),
    .A2(_07788_),
    .B1(_07790_),
    .B2(net1207),
    .C1(_07791_),
    .X(_07792_));
 sky130_fd_sc_hd__a21bo_1 _13097_ (.A1(_04549_),
    .A2(net1205),
    .B1_N(_07792_),
    .X(_07793_));
 sky130_fd_sc_hd__a31o_1 _13098_ (.A1(_07149_),
    .A2(_07781_),
    .A3(_07793_),
    .B1(_07776_),
    .X(_07794_));
 sky130_fd_sc_hd__a32o_1 _13099_ (.A1(_04464_),
    .A2(net825),
    .A3(_07794_),
    .B1(net984),
    .B2(\core.pipe1_resultRegister[6] ),
    .X(_07795_));
 sky130_fd_sc_hd__and2_1 _13100_ (.A(net1821),
    .B(_07795_),
    .X(_00168_));
 sky130_fd_sc_hd__nand2_1 _13101_ (.A(_04423_),
    .B(net1114),
    .Y(_07796_));
 sky130_fd_sc_hd__a22o_1 _13102_ (.A1(\core.csr.cycleTimer.currentValue[7] ),
    .A2(net727),
    .B1(net723),
    .B2(\core.csr.cycleTimer.currentValue[39] ),
    .X(_07797_));
 sky130_fd_sc_hd__a21o_1 _13103_ (.A1(net277),
    .A2(_07238_),
    .B1(_07207_),
    .X(_07798_));
 sky130_fd_sc_hd__a22o_1 _13104_ (.A1(\core.csr.instretTimer.currentValue[7] ),
    .A2(net704),
    .B1(net700),
    .B2(\core.csr.instretTimer.currentValue[39] ),
    .X(_07799_));
 sky130_fd_sc_hd__nor2_1 _13105_ (.A(\core.csr.cycleTimer.currentValue[7] ),
    .B(net708),
    .Y(_07800_));
 sky130_fd_sc_hd__a21o_1 _13106_ (.A1(\core.csr.mconfigptr.currentValue[7] ),
    .A2(net719),
    .B1(_07253_),
    .X(_07801_));
 sky130_fd_sc_hd__or2_1 _13107_ (.A(\core.csr.traps.mip.csrReadData[7] ),
    .B(net656),
    .X(_07802_));
 sky130_fd_sc_hd__o211a_1 _13108_ (.A1(\core.csr.traps.mtval.csrReadData[7] ),
    .A2(net663),
    .B1(net660),
    .C1(_07802_),
    .X(_07803_));
 sky130_fd_sc_hd__a21o_1 _13109_ (.A1(\core.csr.traps.mcause.csrReadData[7] ),
    .A2(net666),
    .B1(net690),
    .X(_07804_));
 sky130_fd_sc_hd__o221a_2 _13110_ (.A1(\core.csr.trapReturnVector[7] ),
    .A2(net687),
    .B1(_07803_),
    .B2(_07804_),
    .C1(net693),
    .X(_07805_));
 sky130_fd_sc_hd__a221o_1 _13111_ (.A1(\core.csr.traps.mscratch.currentValue[7] ),
    .A2(net696),
    .B1(net678),
    .B2(\core.csr.traps.mtvec.csrReadData[7] ),
    .C1(net684),
    .X(_07806_));
 sky130_fd_sc_hd__o221a_4 _13112_ (.A1(\core.csr.traps.mie.currentValue[7] ),
    .A2(net681),
    .B1(_07805_),
    .B2(_07806_),
    .C1(net609),
    .X(_07807_));
 sky130_fd_sc_hd__o221a_2 _13113_ (.A1(net8),
    .A2(_07254_),
    .B1(_07801_),
    .B2(_07807_),
    .C1(_07239_),
    .X(_07808_));
 sky130_fd_sc_hd__o221a_1 _13114_ (.A1(net261),
    .A2(_07208_),
    .B1(_07798_),
    .B2(_07808_),
    .C1(_07212_),
    .X(_07809_));
 sky130_fd_sc_hd__a221o_1 _13115_ (.A1(\core.csr.cycleTimer.currentValue[39] ),
    .A2(net715),
    .B1(_07799_),
    .B2(net979),
    .C1(net712),
    .X(_07810_));
 sky130_fd_sc_hd__nor2_1 _13116_ (.A(_07809_),
    .B(_07810_),
    .Y(_07811_));
 sky130_fd_sc_hd__o2bb2a_4 _13117_ (.A1_N(net979),
    .A2_N(_07797_),
    .B1(_07800_),
    .B2(_07811_),
    .X(_07812_));
 sky130_fd_sc_hd__inv_2 _13118_ (.A(_07812_),
    .Y(_07813_));
 sky130_fd_sc_hd__o21ai_1 _13119_ (.A1(_07156_),
    .A2(_07812_),
    .B1(_07796_),
    .Y(_07814_));
 sky130_fd_sc_hd__a21o_1 _13120_ (.A1(net1109),
    .A2(_07796_),
    .B1(net1105),
    .X(_07815_));
 sky130_fd_sc_hd__xnor2_1 _13121_ (.A(net479),
    .B(_07750_),
    .Y(_07816_));
 sky130_fd_sc_hd__inv_2 _13122_ (.A(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__a32o_1 _13123_ (.A1(net1123),
    .A2(_07814_),
    .A3(_07815_),
    .B1(_06722_),
    .B2(net1152),
    .X(_07818_));
 sky130_fd_sc_hd__a211o_1 _13124_ (.A1(net1134),
    .A2(_07817_),
    .B1(_07818_),
    .C1(net1266),
    .X(_07819_));
 sky130_fd_sc_hd__and2_1 _13125_ (.A(_06722_),
    .B(net1061),
    .X(_07820_));
 sky130_fd_sc_hd__nand2_1 _13126_ (.A(_07315_),
    .B(_07778_),
    .Y(_07821_));
 sky130_fd_sc_hd__xnor2_2 _13127_ (.A(_06721_),
    .B(_07821_),
    .Y(_07822_));
 sky130_fd_sc_hd__a211o_1 _13128_ (.A1(net1066),
    .A2(_07822_),
    .B1(_07820_),
    .C1(net1234),
    .X(_07823_));
 sky130_fd_sc_hd__nor2_1 _13129_ (.A(net890),
    .B(_07638_),
    .Y(_07824_));
 sky130_fd_sc_hd__nand2_1 _13130_ (.A(net890),
    .B(_07639_),
    .Y(_07825_));
 sky130_fd_sc_hd__o21a_1 _13131_ (.A1(net890),
    .A2(_07633_),
    .B1(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__a21o_1 _13132_ (.A1(net890),
    .A2(_07641_),
    .B1(net749),
    .X(_07827_));
 sky130_fd_sc_hd__o22a_1 _13133_ (.A1(net746),
    .A2(_07826_),
    .B1(_07827_),
    .B2(_07824_),
    .X(_07828_));
 sky130_fd_sc_hd__mux2_1 _13134_ (.A0(_07629_),
    .A1(_07634_),
    .S(net892),
    .X(_07829_));
 sky130_fd_sc_hd__mux2_1 _13135_ (.A0(_07452_),
    .A1(_07829_),
    .S(net746),
    .X(_07830_));
 sky130_fd_sc_hd__mux2_1 _13136_ (.A0(_07828_),
    .A1(_07830_),
    .S(net755),
    .X(_07831_));
 sky130_fd_sc_hd__inv_2 _13137_ (.A(_07831_),
    .Y(_07832_));
 sky130_fd_sc_hd__o21a_1 _13138_ (.A1(net750),
    .A2(_07420_),
    .B1(_07447_),
    .X(_07833_));
 sky130_fd_sc_hd__inv_2 _13139_ (.A(_07833_),
    .Y(_07834_));
 sky130_fd_sc_hd__a21o_1 _13140_ (.A1(net752),
    .A2(_07834_),
    .B1(net631),
    .X(_07835_));
 sky130_fd_sc_hd__a221oi_4 _13141_ (.A1(_04462_),
    .A2(net1200),
    .B1(_07537_),
    .B2(_06721_),
    .C1(net1275),
    .Y(_07836_));
 sky130_fd_sc_hd__o221a_4 _13142_ (.A1(net1215),
    .A2(_07832_),
    .B1(_07835_),
    .B2(net1207),
    .C1(_07836_),
    .X(_07837_));
 sky130_fd_sc_hd__o21ai_1 _13143_ (.A1(_04463_),
    .A2(net1204),
    .B1(_07837_),
    .Y(_07838_));
 sky130_fd_sc_hd__a31o_1 _13144_ (.A1(_07147_),
    .A2(_07823_),
    .A3(_07838_),
    .B1(_07819_),
    .X(_07839_));
 sky130_fd_sc_hd__a32o_1 _13145_ (.A1(_04393_),
    .A2(net825),
    .A3(_07839_),
    .B1(net984),
    .B2(\core.pipe1_resultRegister[7] ),
    .X(_07840_));
 sky130_fd_sc_hd__and2_1 _13146_ (.A(net1822),
    .B(_07840_),
    .X(_00169_));
 sky130_fd_sc_hd__nor2_1 _13147_ (.A(_06723_),
    .B(net1066),
    .Y(_07841_));
 sky130_fd_sc_hd__and3_1 _13148_ (.A(_04391_),
    .B(_07317_),
    .C(_07319_),
    .X(_07842_));
 sky130_fd_sc_hd__or2_1 _13149_ (.A(_07320_),
    .B(_07842_),
    .X(_07843_));
 sky130_fd_sc_hd__a211o_1 _13150_ (.A1(net1066),
    .A2(_07843_),
    .B1(_07841_),
    .C1(net1234),
    .X(_07844_));
 sky130_fd_sc_hd__mux2_1 _13151_ (.A0(_07387_),
    .A1(_07439_),
    .S(net749),
    .X(_07845_));
 sky130_fd_sc_hd__inv_2 _13152_ (.A(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__mux2_2 _13153_ (.A0(_07834_),
    .A1(_07846_),
    .S(net752),
    .X(_07847_));
 sky130_fd_sc_hd__mux2_2 _13154_ (.A0(net1200),
    .A1(_07537_),
    .S(_04389_),
    .X(_07848_));
 sky130_fd_sc_hd__o21ai_4 _13155_ (.A1(net1206),
    .A2(_07848_),
    .B1(_04390_),
    .Y(_07849_));
 sky130_fd_sc_hd__o21bai_2 _13156_ (.A1(net755),
    .A2(_07830_),
    .B1_N(net631),
    .Y(_07850_));
 sky130_fd_sc_hd__o221a_4 _13157_ (.A1(net1215),
    .A2(_07847_),
    .B1(_07850_),
    .B2(net1207),
    .C1(_07849_),
    .X(_07851_));
 sky130_fd_sc_hd__a21oi_1 _13158_ (.A1(_07844_),
    .A2(_07851_),
    .B1(_07146_),
    .Y(_07852_));
 sky130_fd_sc_hd__and3_1 _13159_ (.A(net480),
    .B(net479),
    .C(_07750_),
    .X(_07853_));
 sky130_fd_sc_hd__a21oi_1 _13160_ (.A1(net479),
    .A2(_07750_),
    .B1(net480),
    .Y(_07854_));
 sky130_fd_sc_hd__or2_1 _13161_ (.A(_07853_),
    .B(_07854_),
    .X(_07855_));
 sky130_fd_sc_hd__nor2_1 _13162_ (.A(net1136),
    .B(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__nand2_1 _13163_ (.A(_04387_),
    .B(net1114),
    .Y(_07857_));
 sky130_fd_sc_hd__a22o_1 _13164_ (.A1(\core.csr.cycleTimer.currentValue[8] ),
    .A2(net727),
    .B1(net723),
    .B2(\core.csr.cycleTimer.currentValue[40] ),
    .X(_07858_));
 sky130_fd_sc_hd__or3_2 _13165_ (.A(\core.csr.mconfigptr.currentValue[8] ),
    .B(_07206_),
    .C(_07230_),
    .X(_07859_));
 sky130_fd_sc_hd__a22o_1 _13166_ (.A1(\core.csr.instretTimer.currentValue[8] ),
    .A2(net704),
    .B1(net700),
    .B2(\core.csr.instretTimer.currentValue[40] ),
    .X(_07860_));
 sky130_fd_sc_hd__nor2_1 _13167_ (.A(_07202_),
    .B(_07265_),
    .Y(_07861_));
 sky130_fd_sc_hd__or2_1 _13168_ (.A(\core.csr.traps.mip.csrReadData[8] ),
    .B(net656),
    .X(_07862_));
 sky130_fd_sc_hd__o211a_1 _13169_ (.A1(\core.csr.traps.mtval.csrReadData[8] ),
    .A2(net663),
    .B1(net660),
    .C1(_07862_),
    .X(_07863_));
 sky130_fd_sc_hd__a21o_1 _13170_ (.A1(\core.csr.traps.mcause.csrReadData[8] ),
    .A2(net666),
    .B1(net690),
    .X(_07864_));
 sky130_fd_sc_hd__o22a_1 _13171_ (.A1(\core.csr.trapReturnVector[8] ),
    .A2(net687),
    .B1(_07863_),
    .B2(_07864_),
    .X(_07865_));
 sky130_fd_sc_hd__a221o_1 _13172_ (.A1(\core.csr.traps.mscratch.currentValue[8] ),
    .A2(net696),
    .B1(net678),
    .B2(\core.csr.traps.mtvec.csrReadData[8] ),
    .C1(net684),
    .X(_07866_));
 sky130_fd_sc_hd__o221a_2 _13173_ (.A1(\core.csr.traps.mie.currentValue[8] ),
    .A2(net681),
    .B1(_07865_),
    .B2(_07866_),
    .C1(net609),
    .X(_07867_));
 sky130_fd_sc_hd__or3_4 _13174_ (.A(net717),
    .B(_07861_),
    .C(_07867_),
    .X(_07868_));
 sky130_fd_sc_hd__a221o_1 _13175_ (.A1(net278),
    .A2(_07238_),
    .B1(_07859_),
    .B2(_07868_),
    .C1(_07207_),
    .X(_07869_));
 sky130_fd_sc_hd__o211a_1 _13176_ (.A1(net262),
    .A2(_07208_),
    .B1(_07212_),
    .C1(_07869_),
    .X(_07870_));
 sky130_fd_sc_hd__a221o_1 _13177_ (.A1(\core.csr.cycleTimer.currentValue[40] ),
    .A2(net715),
    .B1(_07860_),
    .B2(net978),
    .C1(net711),
    .X(_07871_));
 sky130_fd_sc_hd__o221a_2 _13178_ (.A1(\core.csr.cycleTimer.currentValue[8] ),
    .A2(net708),
    .B1(_07870_),
    .B2(_07871_),
    .C1(_07250_),
    .X(_07872_));
 sky130_fd_sc_hd__a21oi_4 _13179_ (.A1(net978),
    .A2(_07858_),
    .B1(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__inv_2 _13180_ (.A(_07873_),
    .Y(_07874_));
 sky130_fd_sc_hd__o21bai_1 _13181_ (.A1(_07202_),
    .A2(_07214_),
    .B1_N(_07285_),
    .Y(_07875_));
 sky130_fd_sc_hd__o21ai_1 _13182_ (.A1(net1112),
    .A2(_07873_),
    .B1(_07857_),
    .Y(_07876_));
 sky130_fd_sc_hd__a21o_1 _13183_ (.A1(_07288_),
    .A2(_07857_),
    .B1(net1105),
    .X(_07877_));
 sky130_fd_sc_hd__a32o_1 _13184_ (.A1(net1123),
    .A2(_07876_),
    .A3(_07877_),
    .B1(_06723_),
    .B2(net1152),
    .X(_07878_));
 sky130_fd_sc_hd__or4_1 _13185_ (.A(net1266),
    .B(_07852_),
    .C(_07856_),
    .D(_07878_),
    .X(_07879_));
 sky130_fd_sc_hd__a32o_1 _13186_ (.A1(_04355_),
    .A2(_07464_),
    .A3(_07879_),
    .B1(net984),
    .B2(\core.pipe1_resultRegister[8] ),
    .X(_07880_));
 sky130_fd_sc_hd__and2_1 _13187_ (.A(net1822),
    .B(_07880_),
    .X(_00170_));
 sky130_fd_sc_hd__nor3_1 _13188_ (.A(_04306_),
    .B(_07320_),
    .C(_07321_),
    .Y(_07881_));
 sky130_fd_sc_hd__nor2_1 _13189_ (.A(_07322_),
    .B(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__o21ai_1 _13190_ (.A1(net1061),
    .A2(_07882_),
    .B1(net1275),
    .Y(_07883_));
 sky130_fd_sc_hd__a21o_1 _13191_ (.A1(_06724_),
    .A2(_07444_),
    .B1(_07883_),
    .X(_07884_));
 sky130_fd_sc_hd__mux2_1 _13192_ (.A0(_07508_),
    .A1(_07528_),
    .S(net749),
    .X(_07885_));
 sky130_fd_sc_hd__inv_2 _13193_ (.A(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__mux2_2 _13194_ (.A0(_07789_),
    .A1(_07886_),
    .S(net752),
    .X(_07887_));
 sky130_fd_sc_hd__mux2_2 _13195_ (.A0(net1200),
    .A1(_07537_),
    .S(_04304_),
    .X(_07888_));
 sky130_fd_sc_hd__o21ai_4 _13196_ (.A1(net1206),
    .A2(_07888_),
    .B1(_04305_),
    .Y(_07889_));
 sky130_fd_sc_hd__a21o_1 _13197_ (.A1(net752),
    .A2(_07787_),
    .B1(net631),
    .X(_07890_));
 sky130_fd_sc_hd__o221a_4 _13198_ (.A1(net1215),
    .A2(_07887_),
    .B1(_07890_),
    .B2(net1209),
    .C1(_07889_),
    .X(_07891_));
 sky130_fd_sc_hd__a21o_1 _13199_ (.A1(_07884_),
    .A2(_07891_),
    .B1(_07146_),
    .X(_07892_));
 sky130_fd_sc_hd__and2_2 _13200_ (.A(net481),
    .B(_07853_),
    .X(_07893_));
 sky130_fd_sc_hd__nor2_1 _13201_ (.A(net481),
    .B(_07853_),
    .Y(_07894_));
 sky130_fd_sc_hd__or2_2 _13202_ (.A(_07893_),
    .B(_07894_),
    .X(_07895_));
 sky130_fd_sc_hd__inv_2 _13203_ (.A(_07895_),
    .Y(_07896_));
 sky130_fd_sc_hd__and2_1 _13204_ (.A(_04301_),
    .B(net1114),
    .X(_07897_));
 sky130_fd_sc_hd__a22o_1 _13205_ (.A1(\core.csr.cycleTimer.currentValue[9] ),
    .A2(net726),
    .B1(net722),
    .B2(\core.csr.cycleTimer.currentValue[41] ),
    .X(_07898_));
 sky130_fd_sc_hd__a221o_1 _13206_ (.A1(\core.csr.mconfigptr.currentValue[9] ),
    .A2(net719),
    .B1(_07238_),
    .B2(net279),
    .C1(_07207_),
    .X(_07899_));
 sky130_fd_sc_hd__a22o_1 _13207_ (.A1(\core.csr.instretTimer.currentValue[9] ),
    .A2(net704),
    .B1(net700),
    .B2(\core.csr.instretTimer.currentValue[41] ),
    .X(_07900_));
 sky130_fd_sc_hd__or2_1 _13208_ (.A(\core.csr.traps.mip.csrReadData[9] ),
    .B(net655),
    .X(_07901_));
 sky130_fd_sc_hd__o211a_1 _13209_ (.A1(\core.csr.traps.mtval.csrReadData[9] ),
    .A2(net662),
    .B1(net659),
    .C1(_07901_),
    .X(_07902_));
 sky130_fd_sc_hd__a21o_1 _13210_ (.A1(\core.csr.traps.mcause.csrReadData[9] ),
    .A2(net666),
    .B1(net690),
    .X(_07903_));
 sky130_fd_sc_hd__o221a_1 _13211_ (.A1(\core.csr.trapReturnVector[9] ),
    .A2(net687),
    .B1(_07902_),
    .B2(_07903_),
    .C1(net693),
    .X(_07904_));
 sky130_fd_sc_hd__a221o_1 _13212_ (.A1(\core.csr.traps.mscratch.currentValue[9] ),
    .A2(net696),
    .B1(net677),
    .B2(\core.csr.traps.mtvec.csrReadData[9] ),
    .C1(net683),
    .X(_07905_));
 sky130_fd_sc_hd__o221a_4 _13213_ (.A1(\core.csr.traps.mie.currentValue[9] ),
    .A2(net680),
    .B1(_07904_),
    .B2(_07905_),
    .C1(net608),
    .X(_07906_));
 sky130_fd_sc_hd__o221a_1 _13214_ (.A1(net263),
    .A2(_07208_),
    .B1(_07899_),
    .B2(_07906_),
    .C1(_07212_),
    .X(_07907_));
 sky130_fd_sc_hd__a221o_1 _13215_ (.A1(\core.csr.cycleTimer.currentValue[41] ),
    .A2(net715),
    .B1(_07900_),
    .B2(net978),
    .C1(net711),
    .X(_07908_));
 sky130_fd_sc_hd__o22a_1 _13216_ (.A1(\core.csr.cycleTimer.currentValue[9] ),
    .A2(net707),
    .B1(_07907_),
    .B2(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__a21o_4 _13217_ (.A1(net978),
    .A2(_07898_),
    .B1(_07909_),
    .X(_07910_));
 sky130_fd_sc_hd__a21oi_1 _13218_ (.A1(net1111),
    .A2(_07910_),
    .B1(_07897_),
    .Y(_07911_));
 sky130_fd_sc_hd__o21a_1 _13219_ (.A1(net1108),
    .A2(_07897_),
    .B1(net1107),
    .X(_07912_));
 sky130_fd_sc_hd__o32a_1 _13220_ (.A1(net1121),
    .A2(_07911_),
    .A3(_07912_),
    .B1(_06724_),
    .B2(_04068_),
    .X(_07913_));
 sky130_fd_sc_hd__o2111ai_2 _13221_ (.A1(net1136),
    .A2(_07895_),
    .B1(_07913_),
    .C1(_07892_),
    .D1(net1262),
    .Y(_07914_));
 sky130_fd_sc_hd__a32o_1 _13222_ (.A1(_04269_),
    .A2(net825),
    .A3(_07914_),
    .B1(net984),
    .B2(\core.pipe1_resultRegister[9] ),
    .X(_07915_));
 sky130_fd_sc_hd__and2_1 _13223_ (.A(net1823),
    .B(_07915_),
    .X(_00171_));
 sky130_fd_sc_hd__nor2_1 _13224_ (.A(_06726_),
    .B(net1066),
    .Y(_07916_));
 sky130_fd_sc_hd__or3_1 _13225_ (.A(_04218_),
    .B(_07302_),
    .C(_07322_),
    .X(_07917_));
 sky130_fd_sc_hd__nand2_1 _13226_ (.A(_07323_),
    .B(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__a211o_1 _13227_ (.A1(net1066),
    .A2(_07918_),
    .B1(_07916_),
    .C1(net1235),
    .X(_07919_));
 sky130_fd_sc_hd__mux2_1 _13228_ (.A0(_07575_),
    .A1(_07588_),
    .S(net749),
    .X(_07920_));
 sky130_fd_sc_hd__mux2_1 _13229_ (.A0(_07744_),
    .A1(_07920_),
    .S(net754),
    .X(_07921_));
 sky130_fd_sc_hd__mux2_1 _13230_ (.A0(_07537_),
    .A1(net1202),
    .S(_04216_),
    .X(_07922_));
 sky130_fd_sc_hd__o21ai_1 _13231_ (.A1(net1206),
    .A2(_07922_),
    .B1(_04217_),
    .Y(_07923_));
 sky130_fd_sc_hd__o21bai_1 _13232_ (.A1(net755),
    .A2(_07739_),
    .B1_N(net631),
    .Y(_07924_));
 sky130_fd_sc_hd__o22a_2 _13233_ (.A1(net1216),
    .A2(_07921_),
    .B1(_07924_),
    .B2(net1208),
    .X(_07925_));
 sky130_fd_sc_hd__a31o_1 _13234_ (.A1(_07919_),
    .A2(_07923_),
    .A3(_07925_),
    .B1(_07146_),
    .X(_07926_));
 sky130_fd_sc_hd__xnor2_2 _13235_ (.A(net451),
    .B(_07893_),
    .Y(_07927_));
 sky130_fd_sc_hd__inv_2 _13236_ (.A(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__o21ai_1 _13237_ (.A1(net1136),
    .A2(_07927_),
    .B1(net1262),
    .Y(_07929_));
 sky130_fd_sc_hd__and2_1 _13238_ (.A(_04213_),
    .B(net1114),
    .X(_07930_));
 sky130_fd_sc_hd__a22o_1 _13239_ (.A1(\core.csr.cycleTimer.currentValue[10] ),
    .A2(net726),
    .B1(net722),
    .B2(\core.csr.cycleTimer.currentValue[42] ),
    .X(_07931_));
 sky130_fd_sc_hd__a221o_1 _13240_ (.A1(\core.csr.mconfigptr.currentValue[10] ),
    .A2(_07234_),
    .B1(_07238_),
    .B2(net265),
    .C1(_07207_),
    .X(_07932_));
 sky130_fd_sc_hd__a22o_2 _13241_ (.A1(\core.csr.instretTimer.currentValue[10] ),
    .A2(net704),
    .B1(net700),
    .B2(\core.csr.instretTimer.currentValue[42] ),
    .X(_07933_));
 sky130_fd_sc_hd__or2_1 _13242_ (.A(\core.csr.traps.mip.csrReadData[10] ),
    .B(net656),
    .X(_07934_));
 sky130_fd_sc_hd__o211a_1 _13243_ (.A1(\core.csr.traps.mtval.csrReadData[10] ),
    .A2(net663),
    .B1(net660),
    .C1(_07934_),
    .X(_07935_));
 sky130_fd_sc_hd__a21o_1 _13244_ (.A1(\core.csr.traps.mcause.csrReadData[10] ),
    .A2(net666),
    .B1(net690),
    .X(_07936_));
 sky130_fd_sc_hd__o221a_1 _13245_ (.A1(\core.csr.trapReturnVector[10] ),
    .A2(net687),
    .B1(_07935_),
    .B2(_07936_),
    .C1(net693),
    .X(_07937_));
 sky130_fd_sc_hd__a221o_1 _13246_ (.A1(\core.csr.traps.mscratch.currentValue[10] ),
    .A2(net696),
    .B1(net678),
    .B2(\core.csr.traps.mtvec.csrReadData[10] ),
    .C1(net684),
    .X(_07938_));
 sky130_fd_sc_hd__o221a_4 _13247_ (.A1(\core.csr.traps.mie.currentValue[10] ),
    .A2(net681),
    .B1(_07937_),
    .B2(_07938_),
    .C1(net609),
    .X(_07939_));
 sky130_fd_sc_hd__o221a_1 _13248_ (.A1(net254),
    .A2(_07208_),
    .B1(_07932_),
    .B2(_07939_),
    .C1(_07212_),
    .X(_07940_));
 sky130_fd_sc_hd__a221o_1 _13249_ (.A1(\core.csr.cycleTimer.currentValue[42] ),
    .A2(net715),
    .B1(_07933_),
    .B2(net978),
    .C1(net711),
    .X(_07941_));
 sky130_fd_sc_hd__o22a_1 _13250_ (.A1(\core.csr.cycleTimer.currentValue[10] ),
    .A2(net707),
    .B1(_07940_),
    .B2(_07941_),
    .X(_07942_));
 sky130_fd_sc_hd__a21o_4 _13251_ (.A1(net975),
    .A2(_07931_),
    .B1(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__a21o_1 _13252_ (.A1(_07157_),
    .A2(_07943_),
    .B1(_07930_),
    .X(_07944_));
 sky130_fd_sc_hd__o21ai_1 _13253_ (.A1(_07289_),
    .A2(_07930_),
    .B1(net1107),
    .Y(_07945_));
 sky130_fd_sc_hd__a32o_1 _13254_ (.A1(net1122),
    .A2(_07944_),
    .A3(_07945_),
    .B1(_06726_),
    .B2(net1152),
    .X(_07946_));
 sky130_fd_sc_hd__or3b_1 _13255_ (.A(_07929_),
    .B(_07946_),
    .C_N(_07926_),
    .X(_07947_));
 sky130_fd_sc_hd__a32o_1 _13256_ (.A1(_04181_),
    .A2(_07464_),
    .A3(_07947_),
    .B1(net984),
    .B2(\core.pipe1_resultRegister[10] ),
    .X(_07948_));
 sky130_fd_sc_hd__and2_1 _13257_ (.A(net1822),
    .B(_07948_),
    .X(_00172_));
 sky130_fd_sc_hd__nor2_1 _13258_ (.A(_05068_),
    .B(net1065),
    .Y(_07949_));
 sky130_fd_sc_hd__and2_4 _13259_ (.A(net1275),
    .B(_07050_),
    .X(_07950_));
 sky130_fd_sc_hd__nand2_1 _13260_ (.A(net1275),
    .B(_07050_),
    .Y(_07951_));
 sky130_fd_sc_hd__xor2_1 _13261_ (.A(_04133_),
    .B(_07324_),
    .X(_07952_));
 sky130_fd_sc_hd__a211o_1 _13262_ (.A1(net1065),
    .A2(_07952_),
    .B1(net1178),
    .C1(_07949_),
    .X(_07953_));
 sky130_fd_sc_hd__nor2_1 _13263_ (.A(net748),
    .B(_07635_),
    .Y(_07954_));
 sky130_fd_sc_hd__a211o_1 _13264_ (.A1(net748),
    .A2(_07640_),
    .B1(_07954_),
    .C1(net756),
    .X(_07955_));
 sky130_fd_sc_hd__o21ai_4 _13265_ (.A1(net753),
    .A2(_07699_),
    .B1(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__a21o_2 _13266_ (.A1(net753),
    .A2(_07690_),
    .B1(net632),
    .X(_07957_));
 sky130_fd_sc_hd__nand2_1 _13267_ (.A(_04132_),
    .B(net1200),
    .Y(_07958_));
 sky130_fd_sc_hd__o211a_1 _13268_ (.A1(_04132_),
    .A2(net1199),
    .B1(_07958_),
    .C1(net1204),
    .X(_07959_));
 sky130_fd_sc_hd__o221a_1 _13269_ (.A1(net1212),
    .A2(_07957_),
    .B1(_07959_),
    .B2(_04131_),
    .C1(_07953_),
    .X(_07960_));
 sky130_fd_sc_hd__a21bo_1 _13270_ (.A1(_07142_),
    .A2(_07956_),
    .B1_N(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__and3_1 _13271_ (.A(net452),
    .B(net451),
    .C(_07893_),
    .X(_07962_));
 sky130_fd_sc_hd__a21oi_1 _13272_ (.A1(net451),
    .A2(_07893_),
    .B1(net452),
    .Y(_07963_));
 sky130_fd_sc_hd__nor2_1 _13273_ (.A(_07962_),
    .B(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__nand2_1 _13274_ (.A(_04044_),
    .B(net1115),
    .Y(_07965_));
 sky130_fd_sc_hd__a22o_1 _13275_ (.A1(\core.csr.cycleTimer.currentValue[11] ),
    .A2(net726),
    .B1(net722),
    .B2(\core.csr.cycleTimer.currentValue[43] ),
    .X(_07966_));
 sky130_fd_sc_hd__a22o_1 _13276_ (.A1(\core.csr.instretTimer.currentValue[11] ),
    .A2(net704),
    .B1(net700),
    .B2(\core.csr.instretTimer.currentValue[43] ),
    .X(_07967_));
 sky130_fd_sc_hd__mux2_1 _13277_ (.A0(\core.csr.traps.mip.csrReadData[11] ),
    .A1(\core.csr.traps.mtval.csrReadData[11] ),
    .S(net657),
    .X(_07968_));
 sky130_fd_sc_hd__a221o_1 _13278_ (.A1(\core.csr.traps.mcause.csrReadData[11] ),
    .A2(_07281_),
    .B1(_07472_),
    .B2(_07968_),
    .C1(_07283_),
    .X(_07969_));
 sky130_fd_sc_hd__o21a_1 _13279_ (.A1(\core.csr.trapReturnVector[11] ),
    .A2(_07284_),
    .B1(_07969_),
    .X(_07970_));
 sky130_fd_sc_hd__a221o_1 _13280_ (.A1(\core.csr.traps.mtvec.csrReadData[11] ),
    .A2(_07231_),
    .B1(_07280_),
    .B2(\core.csr.traps.mscratch.currentValue[11] ),
    .C1(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__mux2_2 _13281_ (.A0(\core.csr.traps.mie.currentValue[11] ),
    .A1(_07971_),
    .S(_07219_),
    .X(_07972_));
 sky130_fd_sc_hd__a22o_2 _13282_ (.A1(net266),
    .A2(_07277_),
    .B1(_07967_),
    .B2(net981),
    .X(_07973_));
 sky130_fd_sc_hd__a211o_1 _13283_ (.A1(\core.csr.mconfigptr.currentValue[11] ),
    .A2(_07285_),
    .B1(_07972_),
    .C1(_07973_),
    .X(_07974_));
 sky130_fd_sc_hd__a211o_1 _13284_ (.A1(\core.csr.cycleTimer.currentValue[43] ),
    .A2(net714),
    .B1(net709),
    .C1(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__o21a_1 _13285_ (.A1(\core.csr.cycleTimer.currentValue[11] ),
    .A2(net707),
    .B1(_07975_),
    .X(_07976_));
 sky130_fd_sc_hd__a21oi_4 _13286_ (.A1(net975),
    .A2(_07966_),
    .B1(_07976_),
    .Y(_07977_));
 sky130_fd_sc_hd__o21ai_1 _13287_ (.A1(net1112),
    .A2(_07977_),
    .B1(_07965_),
    .Y(_07978_));
 sky130_fd_sc_hd__a21oi_1 _13288_ (.A1(net1109),
    .A2(_07965_),
    .B1(net1105),
    .Y(_07979_));
 sky130_fd_sc_hd__nor2_1 _13289_ (.A(net1121),
    .B(_07979_),
    .Y(_07980_));
 sky130_fd_sc_hd__a221o_1 _13290_ (.A1(net1134),
    .A2(_07964_),
    .B1(_07978_),
    .B2(_07980_),
    .C1(net1266),
    .X(_07981_));
 sky130_fd_sc_hd__a221o_1 _13291_ (.A1(net1151),
    .A2(_05068_),
    .B1(_07147_),
    .B2(_07961_),
    .C1(_07981_),
    .X(_07982_));
 sky130_fd_sc_hd__a32o_1 _13292_ (.A1(_03880_),
    .A2(net825),
    .A3(_07982_),
    .B1(net983),
    .B2(\core.pipe1_resultRegister[11] ),
    .X(_07983_));
 sky130_fd_sc_hd__and2_1 _13293_ (.A(net1824),
    .B(_07983_),
    .X(_00173_));
 sky130_fd_sc_hd__or2_1 _13294_ (.A(net1150),
    .B(_06669_),
    .X(_07984_));
 sky130_fd_sc_hd__nand2_1 _13295_ (.A(_06506_),
    .B(net1115),
    .Y(_07985_));
 sky130_fd_sc_hd__a22o_1 _13296_ (.A1(\core.csr.cycleTimer.currentValue[12] ),
    .A2(net725),
    .B1(net721),
    .B2(\core.csr.cycleTimer.currentValue[44] ),
    .X(_07986_));
 sky130_fd_sc_hd__a22o_1 _13297_ (.A1(\core.csr.instretTimer.currentValue[12] ),
    .A2(net703),
    .B1(net699),
    .B2(\core.csr.instretTimer.currentValue[44] ),
    .X(_07987_));
 sky130_fd_sc_hd__mux2_1 _13298_ (.A0(\core.csr.traps.mip.csrReadData[12] ),
    .A1(\core.csr.traps.mtval.csrReadData[12] ),
    .S(net656),
    .X(_07988_));
 sky130_fd_sc_hd__a221o_1 _13299_ (.A1(\core.csr.traps.mcause.csrReadData[12] ),
    .A2(_07281_),
    .B1(_07472_),
    .B2(_07988_),
    .C1(_07283_),
    .X(_07989_));
 sky130_fd_sc_hd__o21a_1 _13300_ (.A1(\core.csr.trapReturnVector[12] ),
    .A2(_07284_),
    .B1(_07989_),
    .X(_07990_));
 sky130_fd_sc_hd__a221o_1 _13301_ (.A1(\core.csr.traps.mtvec.csrReadData[12] ),
    .A2(_07231_),
    .B1(_07280_),
    .B2(\core.csr.traps.mscratch.currentValue[12] ),
    .C1(_07990_),
    .X(_07991_));
 sky130_fd_sc_hd__mux2_2 _13302_ (.A0(\core.csr.traps.mie.currentValue[12] ),
    .A1(_07991_),
    .S(_07219_),
    .X(_07992_));
 sky130_fd_sc_hd__a22o_2 _13303_ (.A1(net267),
    .A2(_07277_),
    .B1(_07987_),
    .B2(net980),
    .X(_07993_));
 sky130_fd_sc_hd__a211o_1 _13304_ (.A1(\core.csr.mconfigptr.currentValue[12] ),
    .A2(_07285_),
    .B1(_07992_),
    .C1(_07993_),
    .X(_07994_));
 sky130_fd_sc_hd__a211o_1 _13305_ (.A1(\core.csr.cycleTimer.currentValue[44] ),
    .A2(net714),
    .B1(net710),
    .C1(_07994_),
    .X(_07995_));
 sky130_fd_sc_hd__o21a_1 _13306_ (.A1(\core.csr.cycleTimer.currentValue[12] ),
    .A2(net706),
    .B1(_07995_),
    .X(_07996_));
 sky130_fd_sc_hd__a21oi_4 _13307_ (.A1(net975),
    .A2(_07986_),
    .B1(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__o21a_1 _13308_ (.A1(net1112),
    .A2(_07997_),
    .B1(_07985_),
    .X(_07998_));
 sky130_fd_sc_hd__a21oi_1 _13309_ (.A1(net1109),
    .A2(_07985_),
    .B1(net1105),
    .Y(_07999_));
 sky130_fd_sc_hd__or2_1 _13310_ (.A(_06669_),
    .B(net1065),
    .X(_08000_));
 sky130_fd_sc_hd__xnor2_1 _13311_ (.A(_06511_),
    .B(_07326_),
    .Y(_08001_));
 sky130_fd_sc_hd__nand2_1 _13312_ (.A(net1065),
    .B(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__a21o_2 _13313_ (.A1(net753),
    .A2(_07636_),
    .B1(net632),
    .X(_08003_));
 sky130_fd_sc_hd__mux2_1 _13314_ (.A0(_07687_),
    .A1(_07692_),
    .S(net747),
    .X(_08004_));
 sky130_fd_sc_hd__mux2_4 _13315_ (.A0(_07651_),
    .A1(_08004_),
    .S(net753),
    .X(_08005_));
 sky130_fd_sc_hd__nand2_1 _13316_ (.A(_06509_),
    .B(net1200),
    .Y(_08006_));
 sky130_fd_sc_hd__o211a_1 _13317_ (.A1(_06509_),
    .A2(net1198),
    .B1(_08006_),
    .C1(net1204),
    .X(_08007_));
 sky130_fd_sc_hd__o221a_1 _13318_ (.A1(net1212),
    .A2(_08003_),
    .B1(_08007_),
    .B2(_06510_),
    .C1(net1234),
    .X(_08008_));
 sky130_fd_sc_hd__o21a_1 _13319_ (.A1(net1218),
    .A2(_08005_),
    .B1(_08008_),
    .X(_08009_));
 sky130_fd_sc_hd__a31o_1 _13320_ (.A1(_07950_),
    .A2(_08000_),
    .A3(_08002_),
    .B1(_08009_),
    .X(_08010_));
 sky130_fd_sc_hd__or3_1 _13321_ (.A(net1120),
    .B(_07998_),
    .C(_07999_),
    .X(_08011_));
 sky130_fd_sc_hd__nor2_4 _13322_ (.A(net1185),
    .B(net1118),
    .Y(_08012_));
 sky130_fd_sc_hd__or2_4 _13323_ (.A(net1185),
    .B(net1118),
    .X(_08013_));
 sky130_fd_sc_hd__a32o_1 _13324_ (.A1(_07984_),
    .A2(_08011_),
    .A3(net1059),
    .B1(_08010_),
    .B2(net1119),
    .X(_08014_));
 sky130_fd_sc_hd__and2_2 _13325_ (.A(net453),
    .B(_07962_),
    .X(_08015_));
 sky130_fd_sc_hd__nor2_1 _13326_ (.A(net453),
    .B(_07962_),
    .Y(_08016_));
 sky130_fd_sc_hd__or2_1 _13327_ (.A(_08015_),
    .B(_08016_),
    .X(_08017_));
 sky130_fd_sc_hd__a22o_1 _13328_ (.A1(net1225),
    .A2(_08014_),
    .B1(_08017_),
    .B2(net1134),
    .X(_08018_));
 sky130_fd_sc_hd__nand2_1 _13329_ (.A(net1259),
    .B(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__nand2_1 _13330_ (.A(net1264),
    .B(_06669_),
    .Y(_08020_));
 sky130_fd_sc_hd__a221o_4 _13331_ (.A1(\core.pipe0_currentInstruction[12] ),
    .A2(net1220),
    .B1(_08019_),
    .B2(_08020_),
    .C1(net985),
    .X(_08021_));
 sky130_fd_sc_hd__o211a_1 _13332_ (.A1(\core.pipe1_resultRegister[12] ),
    .A2(net986),
    .B1(_08021_),
    .C1(net1841),
    .X(_00174_));
 sky130_fd_sc_hd__nand2_1 _13333_ (.A(_06428_),
    .B(net1115),
    .Y(_08022_));
 sky130_fd_sc_hd__a22o_1 _13334_ (.A1(\core.csr.cycleTimer.currentValue[13] ),
    .A2(net725),
    .B1(net721),
    .B2(\core.csr.cycleTimer.currentValue[45] ),
    .X(_08023_));
 sky130_fd_sc_hd__a22o_1 _13335_ (.A1(\core.csr.instretTimer.currentValue[13] ),
    .A2(net703),
    .B1(net699),
    .B2(\core.csr.instretTimer.currentValue[45] ),
    .X(_08024_));
 sky130_fd_sc_hd__mux2_1 _13336_ (.A0(\core.csr.traps.mip.csrReadData[13] ),
    .A1(\core.csr.traps.mtval.csrReadData[13] ),
    .S(net656),
    .X(_08025_));
 sky130_fd_sc_hd__a221o_1 _13337_ (.A1(\core.csr.traps.mcause.csrReadData[13] ),
    .A2(_07281_),
    .B1(_07472_),
    .B2(_08025_),
    .C1(_07283_),
    .X(_08026_));
 sky130_fd_sc_hd__o21a_2 _13338_ (.A1(\core.csr.trapReturnVector[13] ),
    .A2(_07284_),
    .B1(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__a221o_1 _13339_ (.A1(\core.csr.traps.mtvec.csrReadData[13] ),
    .A2(_07231_),
    .B1(_07280_),
    .B2(\core.csr.traps.mscratch.currentValue[13] ),
    .C1(_08027_),
    .X(_08028_));
 sky130_fd_sc_hd__mux2_2 _13340_ (.A0(\core.csr.traps.mie.currentValue[13] ),
    .A1(_08028_),
    .S(_07219_),
    .X(_08029_));
 sky130_fd_sc_hd__a22o_2 _13341_ (.A1(net268),
    .A2(_07277_),
    .B1(_08024_),
    .B2(net981),
    .X(_08030_));
 sky130_fd_sc_hd__a211o_1 _13342_ (.A1(\core.csr.mconfigptr.currentValue[13] ),
    .A2(_07285_),
    .B1(_08029_),
    .C1(_08030_),
    .X(_08031_));
 sky130_fd_sc_hd__a211o_1 _13343_ (.A1(\core.csr.cycleTimer.currentValue[45] ),
    .A2(net714),
    .B1(net710),
    .C1(_08031_),
    .X(_08032_));
 sky130_fd_sc_hd__o21a_1 _13344_ (.A1(\core.csr.cycleTimer.currentValue[13] ),
    .A2(net706),
    .B1(_08032_),
    .X(_08033_));
 sky130_fd_sc_hd__a21oi_4 _13345_ (.A1(net975),
    .A2(_08023_),
    .B1(_08033_),
    .Y(_08034_));
 sky130_fd_sc_hd__o21ai_1 _13346_ (.A1(net1113),
    .A2(_08034_),
    .B1(_08022_),
    .Y(_08035_));
 sky130_fd_sc_hd__a21o_1 _13347_ (.A1(net1109),
    .A2(_08022_),
    .B1(net1104),
    .X(_08036_));
 sky130_fd_sc_hd__a32o_1 _13348_ (.A1(net1124),
    .A2(_08035_),
    .A3(_08036_),
    .B1(_06668_),
    .B2(net1151),
    .X(_08037_));
 sky130_fd_sc_hd__nand2_1 _13349_ (.A(_06668_),
    .B(net1061),
    .Y(_08038_));
 sky130_fd_sc_hd__a21oi_2 _13350_ (.A1(_06512_),
    .A2(_07326_),
    .B1(_07327_),
    .Y(_08039_));
 sky130_fd_sc_hd__xor2_1 _13351_ (.A(_06434_),
    .B(_08039_),
    .X(_08040_));
 sky130_fd_sc_hd__a21oi_1 _13352_ (.A1(net1065),
    .A2(_08040_),
    .B1(net1178),
    .Y(_08041_));
 sky130_fd_sc_hd__a21o_1 _13353_ (.A1(net754),
    .A2(_07589_),
    .B1(net632),
    .X(_08042_));
 sky130_fd_sc_hd__nand2_1 _13354_ (.A(net749),
    .B(_07738_),
    .Y(_08043_));
 sky130_fd_sc_hd__o211a_1 _13355_ (.A1(net749),
    .A2(_07734_),
    .B1(_08043_),
    .C1(net752),
    .X(_08044_));
 sky130_fd_sc_hd__a21o_1 _13356_ (.A1(net756),
    .A2(_07596_),
    .B1(_08044_),
    .X(_08045_));
 sky130_fd_sc_hd__mux2_1 _13357_ (.A0(net1198),
    .A1(_07458_),
    .S(_06432_),
    .X(_08046_));
 sky130_fd_sc_hd__a21o_1 _13358_ (.A1(net1204),
    .A2(_08046_),
    .B1(_06433_),
    .X(_08047_));
 sky130_fd_sc_hd__o221a_1 _13359_ (.A1(net1211),
    .A2(_08042_),
    .B1(_08045_),
    .B2(net1217),
    .C1(_08047_),
    .X(_08048_));
 sky130_fd_sc_hd__a22o_1 _13360_ (.A1(_08038_),
    .A2(_08041_),
    .B1(_08048_),
    .B2(net1234),
    .X(_08049_));
 sky130_fd_sc_hd__a2bb2o_1 _13361_ (.A1_N(_08013_),
    .A2_N(_08037_),
    .B1(_08049_),
    .B2(net1119),
    .X(_08050_));
 sky130_fd_sc_hd__xnor2_2 _13362_ (.A(net454),
    .B(_08015_),
    .Y(_08051_));
 sky130_fd_sc_hd__inv_2 _13363_ (.A(_08051_),
    .Y(_08052_));
 sky130_fd_sc_hd__a22o_1 _13364_ (.A1(net1224),
    .A2(_08050_),
    .B1(_08051_),
    .B2(net1134),
    .X(_08053_));
 sky130_fd_sc_hd__nand2_1 _13365_ (.A(net1259),
    .B(_08053_),
    .Y(_08054_));
 sky130_fd_sc_hd__or2_1 _13366_ (.A(net1259),
    .B(_06668_),
    .X(_08055_));
 sky130_fd_sc_hd__a221o_4 _13367_ (.A1(\core.pipe0_currentInstruction[13] ),
    .A2(net1220),
    .B1(_08054_),
    .B2(_08055_),
    .C1(net983),
    .X(_08056_));
 sky130_fd_sc_hd__o211a_1 _13368_ (.A1(\core.pipe1_resultRegister[13] ),
    .A2(net986),
    .B1(_08056_),
    .C1(net1842),
    .X(_00175_));
 sky130_fd_sc_hd__nand2_1 _13369_ (.A(_06353_),
    .B(net1115),
    .Y(_08057_));
 sky130_fd_sc_hd__a22o_1 _13370_ (.A1(\core.csr.cycleTimer.currentValue[14] ),
    .A2(net725),
    .B1(net721),
    .B2(\core.csr.cycleTimer.currentValue[46] ),
    .X(_08058_));
 sky130_fd_sc_hd__a22o_1 _13371_ (.A1(\core.csr.instretTimer.currentValue[14] ),
    .A2(net704),
    .B1(net700),
    .B2(\core.csr.instretTimer.currentValue[46] ),
    .X(_08059_));
 sky130_fd_sc_hd__mux2_1 _13372_ (.A0(\core.csr.traps.mip.csrReadData[14] ),
    .A1(\core.csr.traps.mtval.csrReadData[14] ),
    .S(net656),
    .X(_08060_));
 sky130_fd_sc_hd__a221o_1 _13373_ (.A1(\core.csr.traps.mcause.csrReadData[14] ),
    .A2(_07281_),
    .B1(_07472_),
    .B2(_08060_),
    .C1(_07283_),
    .X(_08061_));
 sky130_fd_sc_hd__o21a_2 _13374_ (.A1(\core.csr.trapReturnVector[14] ),
    .A2(_07284_),
    .B1(_08061_),
    .X(_08062_));
 sky130_fd_sc_hd__a221o_1 _13375_ (.A1(\core.csr.traps.mtvec.csrReadData[14] ),
    .A2(_07231_),
    .B1(_07280_),
    .B2(\core.csr.traps.mscratch.currentValue[14] ),
    .C1(_08062_),
    .X(_08063_));
 sky130_fd_sc_hd__mux2_2 _13376_ (.A0(\core.csr.traps.mie.currentValue[14] ),
    .A1(_08063_),
    .S(_07219_),
    .X(_08064_));
 sky130_fd_sc_hd__a22o_2 _13377_ (.A1(net269),
    .A2(_07277_),
    .B1(_08059_),
    .B2(net981),
    .X(_08065_));
 sky130_fd_sc_hd__a211o_1 _13378_ (.A1(\core.csr.mconfigptr.currentValue[14] ),
    .A2(_07285_),
    .B1(_08064_),
    .C1(_08065_),
    .X(_08066_));
 sky130_fd_sc_hd__a211o_1 _13379_ (.A1(\core.csr.cycleTimer.currentValue[46] ),
    .A2(net714),
    .B1(net710),
    .C1(_08066_),
    .X(_08067_));
 sky130_fd_sc_hd__o21a_1 _13380_ (.A1(\core.csr.cycleTimer.currentValue[14] ),
    .A2(net706),
    .B1(_08067_),
    .X(_08068_));
 sky130_fd_sc_hd__a21oi_4 _13381_ (.A1(net976),
    .A2(_08058_),
    .B1(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__o21ai_1 _13382_ (.A1(net1113),
    .A2(_08069_),
    .B1(_08057_),
    .Y(_08070_));
 sky130_fd_sc_hd__a21o_1 _13383_ (.A1(net1110),
    .A2(_08057_),
    .B1(net1104),
    .X(_08071_));
 sky130_fd_sc_hd__a32o_1 _13384_ (.A1(net1124),
    .A2(_08070_),
    .A3(_08071_),
    .B1(_06667_),
    .B2(net1153),
    .X(_08072_));
 sky130_fd_sc_hd__nand2_1 _13385_ (.A(_06667_),
    .B(net1060),
    .Y(_08073_));
 sky130_fd_sc_hd__o21ba_1 _13386_ (.A1(_06434_),
    .A2(_08039_),
    .B1_N(_07299_),
    .X(_08074_));
 sky130_fd_sc_hd__xnor2_1 _13387_ (.A(_06358_),
    .B(_08074_),
    .Y(_08075_));
 sky130_fd_sc_hd__a21oi_1 _13388_ (.A1(net1065),
    .A2(_08075_),
    .B1(net1178),
    .Y(_08076_));
 sky130_fd_sc_hd__mux2_1 _13389_ (.A0(_07782_),
    .A1(_07786_),
    .S(net750),
    .X(_08077_));
 sky130_fd_sc_hd__mux2_1 _13390_ (.A0(_07534_),
    .A1(_08077_),
    .S(net754),
    .X(_08078_));
 sky130_fd_sc_hd__o21bai_4 _13391_ (.A1(net755),
    .A2(_07529_),
    .B1_N(net631),
    .Y(_08079_));
 sky130_fd_sc_hd__a21oi_1 _13392_ (.A1(_06355_),
    .A2(net1200),
    .B1(net1206),
    .Y(_08080_));
 sky130_fd_sc_hd__o22a_1 _13393_ (.A1(_06358_),
    .A2(net1198),
    .B1(_08080_),
    .B2(_06356_),
    .X(_08081_));
 sky130_fd_sc_hd__o221a_1 _13394_ (.A1(net1216),
    .A2(_08078_),
    .B1(_08079_),
    .B2(net1210),
    .C1(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__a22o_1 _13395_ (.A1(_08073_),
    .A2(_08076_),
    .B1(_08082_),
    .B2(net1234),
    .X(_08083_));
 sky130_fd_sc_hd__a2bb2o_1 _13396_ (.A1_N(_08013_),
    .A2_N(_08072_),
    .B1(_08083_),
    .B2(net1119),
    .X(_08084_));
 sky130_fd_sc_hd__and3_1 _13397_ (.A(net455),
    .B(net454),
    .C(_08015_),
    .X(_08085_));
 sky130_fd_sc_hd__a21oi_1 _13398_ (.A1(net454),
    .A2(_08015_),
    .B1(net455),
    .Y(_08086_));
 sky130_fd_sc_hd__or2_1 _13399_ (.A(_08085_),
    .B(_08086_),
    .X(_08087_));
 sky130_fd_sc_hd__a22o_1 _13400_ (.A1(net1224),
    .A2(_08084_),
    .B1(_08087_),
    .B2(net1134),
    .X(_08088_));
 sky130_fd_sc_hd__nand2_1 _13401_ (.A(net1259),
    .B(_08088_),
    .Y(_08089_));
 sky130_fd_sc_hd__or2_1 _13402_ (.A(net1259),
    .B(_06667_),
    .X(_08090_));
 sky130_fd_sc_hd__a221o_4 _13403_ (.A1(net1795),
    .A2(net1220),
    .B1(_08089_),
    .B2(_08090_),
    .C1(net983),
    .X(_08091_));
 sky130_fd_sc_hd__o211a_1 _13404_ (.A1(\core.pipe1_resultRegister[14] ),
    .A2(net986),
    .B1(_08091_),
    .C1(net1842),
    .X(_00176_));
 sky130_fd_sc_hd__and2_2 _13405_ (.A(net456),
    .B(_08085_),
    .X(_08092_));
 sky130_fd_sc_hd__nor2_1 _13406_ (.A(net456),
    .B(_08085_),
    .Y(_08093_));
 sky130_fd_sc_hd__or2_1 _13407_ (.A(_08092_),
    .B(_08093_),
    .X(_08094_));
 sky130_fd_sc_hd__inv_2 _13408_ (.A(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__nand2_1 _13409_ (.A(_06666_),
    .B(net1060),
    .Y(_08096_));
 sky130_fd_sc_hd__o21ba_1 _13410_ (.A1(_06357_),
    .A2(_08074_),
    .B1_N(_07298_),
    .X(_08097_));
 sky130_fd_sc_hd__xnor2_2 _13411_ (.A(_06282_),
    .B(_08097_),
    .Y(_08098_));
 sky130_fd_sc_hd__a21oi_1 _13412_ (.A1(net1064),
    .A2(_08098_),
    .B1(net1177),
    .Y(_08099_));
 sky130_fd_sc_hd__a21o_1 _13413_ (.A1(net754),
    .A2(_07440_),
    .B1(net632),
    .X(_08100_));
 sky130_fd_sc_hd__nand2_1 _13414_ (.A(net750),
    .B(_07829_),
    .Y(_08101_));
 sky130_fd_sc_hd__a21oi_1 _13415_ (.A1(net746),
    .A2(_07826_),
    .B1(net755),
    .Y(_08102_));
 sky130_fd_sc_hd__a22o_2 _13416_ (.A1(net755),
    .A2(_07453_),
    .B1(_08101_),
    .B2(_08102_),
    .X(_08103_));
 sky130_fd_sc_hd__a21oi_1 _13417_ (.A1(_06279_),
    .A2(net1200),
    .B1(net1206),
    .Y(_08104_));
 sky130_fd_sc_hd__o22a_1 _13418_ (.A1(_06282_),
    .A2(net1198),
    .B1(_08104_),
    .B2(_06280_),
    .X(_08105_));
 sky130_fd_sc_hd__o221a_1 _13419_ (.A1(net1211),
    .A2(_08100_),
    .B1(_08103_),
    .B2(net1218),
    .C1(_08105_),
    .X(_08106_));
 sky130_fd_sc_hd__a22o_1 _13420_ (.A1(_08096_),
    .A2(_08099_),
    .B1(_08106_),
    .B2(net1233),
    .X(_08107_));
 sky130_fd_sc_hd__nand2_1 _13421_ (.A(net1151),
    .B(_06666_),
    .Y(_08108_));
 sky130_fd_sc_hd__nand2_1 _13422_ (.A(_06277_),
    .B(net1114),
    .Y(_08109_));
 sky130_fd_sc_hd__a22o_1 _13423_ (.A1(\core.csr.cycleTimer.currentValue[15] ),
    .A2(net725),
    .B1(net721),
    .B2(\core.csr.cycleTimer.currentValue[47] ),
    .X(_08110_));
 sky130_fd_sc_hd__o21ai_1 _13424_ (.A1(\core.csr.cycleTimer.currentValue[15] ),
    .A2(net706),
    .B1(_07250_),
    .Y(_08111_));
 sky130_fd_sc_hd__a22o_1 _13425_ (.A1(\core.csr.instretTimer.currentValue[15] ),
    .A2(net704),
    .B1(net700),
    .B2(\core.csr.instretTimer.currentValue[47] ),
    .X(_08112_));
 sky130_fd_sc_hd__a22o_1 _13426_ (.A1(net270),
    .A2(_07238_),
    .B1(net714),
    .B2(\core.csr.cycleTimer.currentValue[47] ),
    .X(_08113_));
 sky130_fd_sc_hd__a21o_2 _13427_ (.A1(net981),
    .A2(_08112_),
    .B1(net711),
    .X(_08114_));
 sky130_fd_sc_hd__or2_1 _13428_ (.A(\core.csr.traps.mip.csrReadData[15] ),
    .B(net655),
    .X(_08115_));
 sky130_fd_sc_hd__o211a_1 _13429_ (.A1(\core.csr.traps.mtval.csrReadData[15] ),
    .A2(net662),
    .B1(net659),
    .C1(_08115_),
    .X(_08116_));
 sky130_fd_sc_hd__a21o_1 _13430_ (.A1(\core.csr.traps.mcause.csrReadData[15] ),
    .A2(net665),
    .B1(net689),
    .X(_08117_));
 sky130_fd_sc_hd__o221a_1 _13431_ (.A1(\core.csr.trapReturnVector[15] ),
    .A2(net686),
    .B1(_08116_),
    .B2(_08117_),
    .C1(net692),
    .X(_08118_));
 sky130_fd_sc_hd__a221o_1 _13432_ (.A1(\core.csr.traps.mscratch.currentValue[15] ),
    .A2(net695),
    .B1(net677),
    .B2(\core.csr.traps.mtvec.csrReadData[15] ),
    .C1(net683),
    .X(_08119_));
 sky130_fd_sc_hd__o221a_4 _13433_ (.A1(\core.csr.traps.mie.currentValue[15] ),
    .A2(net680),
    .B1(_08118_),
    .B2(_08119_),
    .C1(net608),
    .X(_08120_));
 sky130_fd_sc_hd__a2111oi_2 _13434_ (.A1(\core.csr.mconfigptr.currentValue[15] ),
    .A2(net718),
    .B1(_08113_),
    .C1(_08114_),
    .D1(_08120_),
    .Y(_08121_));
 sky130_fd_sc_hd__o2bb2a_4 _13435_ (.A1_N(net974),
    .A2_N(_08110_),
    .B1(_08111_),
    .B2(_08121_),
    .X(_08122_));
 sky130_fd_sc_hd__inv_2 _13436_ (.A(_08122_),
    .Y(_08123_));
 sky130_fd_sc_hd__or2_1 _13437_ (.A(net1112),
    .B(_08122_),
    .X(_08124_));
 sky130_fd_sc_hd__nand2_1 _13438_ (.A(net1109),
    .B(_08109_),
    .Y(_08125_));
 sky130_fd_sc_hd__a221o_1 _13439_ (.A1(_08109_),
    .A2(_08124_),
    .B1(_08125_),
    .B2(net1106),
    .C1(net1121),
    .X(_08126_));
 sky130_fd_sc_hd__a32o_1 _13440_ (.A1(net1059),
    .A2(_08108_),
    .A3(_08126_),
    .B1(_08107_),
    .B2(net1119),
    .X(_08127_));
 sky130_fd_sc_hd__a22o_1 _13441_ (.A1(net1134),
    .A2(_08094_),
    .B1(_08127_),
    .B2(net1224),
    .X(_08128_));
 sky130_fd_sc_hd__nand2_1 _13442_ (.A(net1259),
    .B(_08128_),
    .Y(_08129_));
 sky130_fd_sc_hd__or2_1 _13443_ (.A(net1259),
    .B(_06666_),
    .X(_08130_));
 sky130_fd_sc_hd__a221o_4 _13444_ (.A1(net1793),
    .A2(net1220),
    .B1(_08129_),
    .B2(_08130_),
    .C1(net983),
    .X(_08131_));
 sky130_fd_sc_hd__o211a_1 _13445_ (.A1(\core.pipe1_resultRegister[15] ),
    .A2(net986),
    .B1(_08131_),
    .C1(net1839),
    .X(_00177_));
 sky130_fd_sc_hd__nand2_1 _13446_ (.A(_06198_),
    .B(net1114),
    .Y(_08132_));
 sky130_fd_sc_hd__a22o_1 _13447_ (.A1(\core.csr.cycleTimer.currentValue[16] ),
    .A2(net724),
    .B1(net720),
    .B2(\core.csr.cycleTimer.currentValue[48] ),
    .X(_08133_));
 sky130_fd_sc_hd__a22o_2 _13448_ (.A1(\core.csr.instretTimer.currentValue[16] ),
    .A2(net703),
    .B1(net699),
    .B2(\core.csr.instretTimer.currentValue[48] ),
    .X(_08134_));
 sky130_fd_sc_hd__nor2_1 _13449_ (.A(\core.csr.cycleTimer.currentValue[16] ),
    .B(net705),
    .Y(_08135_));
 sky130_fd_sc_hd__a22o_1 _13450_ (.A1(\core.csr.cycleTimer.currentValue[48] ),
    .A2(net713),
    .B1(_08134_),
    .B2(net974),
    .X(_08136_));
 sky130_fd_sc_hd__or2_1 _13451_ (.A(\core.csr.traps.mip.csrReadData[16] ),
    .B(net654),
    .X(_08137_));
 sky130_fd_sc_hd__o211a_1 _13452_ (.A1(\core.csr.traps.mtval.csrReadData[16] ),
    .A2(net662),
    .B1(net658),
    .C1(_08137_),
    .X(_08138_));
 sky130_fd_sc_hd__a21o_1 _13453_ (.A1(\core.csr.traps.mcause.csrReadData[16] ),
    .A2(net665),
    .B1(net689),
    .X(_08139_));
 sky130_fd_sc_hd__o221a_1 _13454_ (.A1(\core.csr.trapReturnVector[16] ),
    .A2(net686),
    .B1(_08138_),
    .B2(_08139_),
    .C1(net692),
    .X(_08140_));
 sky130_fd_sc_hd__a221o_1 _13455_ (.A1(\core.csr.traps.mscratch.currentValue[16] ),
    .A2(net695),
    .B1(net677),
    .B2(\core.csr.traps.mtvec.csrReadData[16] ),
    .C1(net683),
    .X(_08141_));
 sky130_fd_sc_hd__o221a_4 _13456_ (.A1(\core.csr.traps.mie.currentValue[16] ),
    .A2(net680),
    .B1(_08140_),
    .B2(_08141_),
    .C1(net608),
    .X(_08142_));
 sky130_fd_sc_hd__a2111oi_2 _13457_ (.A1(\core.csr.mconfigptr.currentValue[16] ),
    .A2(net718),
    .B1(net709),
    .C1(_08136_),
    .D1(_08142_),
    .Y(_08143_));
 sky130_fd_sc_hd__o2bb2a_4 _13458_ (.A1_N(net977),
    .A2_N(_08133_),
    .B1(_08135_),
    .B2(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__inv_2 _13459_ (.A(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__o21ai_1 _13460_ (.A1(_07156_),
    .A2(_08144_),
    .B1(_08132_),
    .Y(_08146_));
 sky130_fd_sc_hd__a21o_1 _13461_ (.A1(_07288_),
    .A2(_08132_),
    .B1(net1105),
    .X(_08147_));
 sky130_fd_sc_hd__and3_2 _13462_ (.A(net1122),
    .B(_08146_),
    .C(_08147_),
    .X(_08148_));
 sky130_fd_sc_hd__a211o_1 _13463_ (.A1(net1153),
    .A2(_06665_),
    .B1(_08013_),
    .C1(_08148_),
    .X(_08149_));
 sky130_fd_sc_hd__nand2_1 _13464_ (.A(_06665_),
    .B(net1060),
    .Y(_08150_));
 sky130_fd_sc_hd__and3_1 _13465_ (.A(_06203_),
    .B(_07329_),
    .C(_07332_),
    .X(_08151_));
 sky130_fd_sc_hd__nor2_1 _13466_ (.A(_07333_),
    .B(_08151_),
    .Y(_08152_));
 sky130_fd_sc_hd__a21oi_1 _13467_ (.A1(net1067),
    .A2(_08152_),
    .B1(net1178),
    .Y(_08153_));
 sky130_fd_sc_hd__mux2_1 _13468_ (.A0(net1198),
    .A1(_07458_),
    .S(_06201_),
    .X(_08154_));
 sky130_fd_sc_hd__a21o_1 _13469_ (.A1(net1203),
    .A2(_08154_),
    .B1(_06202_),
    .X(_08155_));
 sky130_fd_sc_hd__o221a_1 _13470_ (.A1(net1218),
    .A2(_08100_),
    .B1(_08103_),
    .B2(net1210),
    .C1(_08155_),
    .X(_08156_));
 sky130_fd_sc_hd__a22o_1 _13471_ (.A1(_08150_),
    .A2(_08153_),
    .B1(_08156_),
    .B2(net1233),
    .X(_08157_));
 sky130_fd_sc_hd__a21bo_1 _13472_ (.A1(_07149_),
    .A2(_08157_),
    .B1_N(_08149_),
    .X(_08158_));
 sky130_fd_sc_hd__xnor2_2 _13473_ (.A(net1747),
    .B(_08092_),
    .Y(_08159_));
 sky130_fd_sc_hd__a22o_1 _13474_ (.A1(net1223),
    .A2(_08158_),
    .B1(_08159_),
    .B2(net1135),
    .X(_08160_));
 sky130_fd_sc_hd__nand2_1 _13475_ (.A(net1255),
    .B(_08160_),
    .Y(_08161_));
 sky130_fd_sc_hd__or2_1 _13476_ (.A(net1259),
    .B(_06665_),
    .X(_08162_));
 sky130_fd_sc_hd__a221o_4 _13477_ (.A1(net1789),
    .A2(net1220),
    .B1(_08161_),
    .B2(_08162_),
    .C1(net983),
    .X(_08163_));
 sky130_fd_sc_hd__o211a_1 _13478_ (.A1(\core.pipe1_resultRegister[16] ),
    .A2(net986),
    .B1(_08163_),
    .C1(net1839),
    .X(_00178_));
 sky130_fd_sc_hd__and3_1 _13479_ (.A(net458),
    .B(net1747),
    .C(_08092_),
    .X(_08164_));
 sky130_fd_sc_hd__a21oi_1 _13480_ (.A1(net1747),
    .A2(_08092_),
    .B1(net458),
    .Y(_08165_));
 sky130_fd_sc_hd__or2_1 _13481_ (.A(_08164_),
    .B(_08165_),
    .X(_08166_));
 sky130_fd_sc_hd__inv_2 _13482_ (.A(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__nand2_1 _13483_ (.A(_06664_),
    .B(_07444_),
    .Y(_08168_));
 sky130_fd_sc_hd__o21bai_1 _13484_ (.A1(_06169_),
    .A2(_06200_),
    .B1_N(_07333_),
    .Y(_08169_));
 sky130_fd_sc_hd__xnor2_1 _13485_ (.A(_06127_),
    .B(_08169_),
    .Y(_08170_));
 sky130_fd_sc_hd__a21oi_1 _13486_ (.A1(net1067),
    .A2(_08170_),
    .B1(net1178),
    .Y(_08171_));
 sky130_fd_sc_hd__mux2_1 _13487_ (.A0(net1198),
    .A1(_07458_),
    .S(_06125_),
    .X(_08172_));
 sky130_fd_sc_hd__a21o_1 _13488_ (.A1(net1203),
    .A2(_08172_),
    .B1(_06126_),
    .X(_08173_));
 sky130_fd_sc_hd__o221a_1 _13489_ (.A1(net1211),
    .A2(_08078_),
    .B1(_08079_),
    .B2(net1216),
    .C1(_08173_),
    .X(_08174_));
 sky130_fd_sc_hd__a22o_1 _13490_ (.A1(_08168_),
    .A2(_08171_),
    .B1(_08174_),
    .B2(net1233),
    .X(_08175_));
 sky130_fd_sc_hd__nand2_1 _13491_ (.A(net1153),
    .B(_06664_),
    .Y(_08176_));
 sky130_fd_sc_hd__or2_1 _13492_ (.A(_06121_),
    .B(net1117),
    .X(_08177_));
 sky130_fd_sc_hd__a22o_1 _13493_ (.A1(\core.csr.cycleTimer.currentValue[17] ),
    .A2(net724),
    .B1(net720),
    .B2(\core.csr.cycleTimer.currentValue[49] ),
    .X(_08178_));
 sky130_fd_sc_hd__o21ai_1 _13494_ (.A1(\core.csr.cycleTimer.currentValue[17] ),
    .A2(net705),
    .B1(_07250_),
    .Y(_08179_));
 sky130_fd_sc_hd__a22o_2 _13495_ (.A1(\core.csr.instretTimer.currentValue[17] ),
    .A2(net703),
    .B1(net699),
    .B2(\core.csr.instretTimer.currentValue[49] ),
    .X(_08180_));
 sky130_fd_sc_hd__a22o_1 _13496_ (.A1(\core.csr.cycleTimer.currentValue[49] ),
    .A2(net713),
    .B1(_08180_),
    .B2(net974),
    .X(_08181_));
 sky130_fd_sc_hd__or2_1 _13497_ (.A(\core.csr.traps.mip.csrReadData[17] ),
    .B(net655),
    .X(_08182_));
 sky130_fd_sc_hd__o211a_1 _13498_ (.A1(\core.csr.traps.mtval.csrReadData[17] ),
    .A2(net662),
    .B1(net659),
    .C1(_08182_),
    .X(_08183_));
 sky130_fd_sc_hd__a21o_1 _13499_ (.A1(\core.csr.traps.mcause.csrReadData[17] ),
    .A2(net665),
    .B1(net689),
    .X(_08184_));
 sky130_fd_sc_hd__o221a_1 _13500_ (.A1(\core.csr.trapReturnVector[17] ),
    .A2(net686),
    .B1(_08183_),
    .B2(_08184_),
    .C1(net692),
    .X(_08185_));
 sky130_fd_sc_hd__a221o_1 _13501_ (.A1(\core.csr.traps.mscratch.currentValue[17] ),
    .A2(net695),
    .B1(net677),
    .B2(\core.csr.traps.mtvec.csrReadData[17] ),
    .C1(net683),
    .X(_08186_));
 sky130_fd_sc_hd__o221a_4 _13502_ (.A1(\core.csr.traps.mie.currentValue[17] ),
    .A2(net680),
    .B1(_08185_),
    .B2(_08186_),
    .C1(net608),
    .X(_08187_));
 sky130_fd_sc_hd__a2111oi_2 _13503_ (.A1(\core.csr.mconfigptr.currentValue[17] ),
    .A2(net717),
    .B1(net709),
    .C1(_08181_),
    .D1(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__o2bb2a_4 _13504_ (.A1_N(net973),
    .A2_N(_08178_),
    .B1(_08179_),
    .B2(_08188_),
    .X(_08189_));
 sky130_fd_sc_hd__inv_2 _13505_ (.A(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__or2_1 _13506_ (.A(net1113),
    .B(_08189_),
    .X(_08191_));
 sky130_fd_sc_hd__nand2_1 _13507_ (.A(net1110),
    .B(_08177_),
    .Y(_08192_));
 sky130_fd_sc_hd__a221o_1 _13508_ (.A1(_08177_),
    .A2(_08191_),
    .B1(_08192_),
    .B2(net1106),
    .C1(net1120),
    .X(_08193_));
 sky130_fd_sc_hd__a32o_1 _13509_ (.A1(_08012_),
    .A2(_08176_),
    .A3(_08193_),
    .B1(_08175_),
    .B2(net1119),
    .X(_08194_));
 sky130_fd_sc_hd__a22o_1 _13510_ (.A1(net1135),
    .A2(_08166_),
    .B1(_08194_),
    .B2(net1223),
    .X(_08195_));
 sky130_fd_sc_hd__nand2_1 _13511_ (.A(net1255),
    .B(_08195_),
    .Y(_08196_));
 sky130_fd_sc_hd__or2_1 _13512_ (.A(net1254),
    .B(_06664_),
    .X(_08197_));
 sky130_fd_sc_hd__a221o_4 _13513_ (.A1(net1784),
    .A2(net1219),
    .B1(_08196_),
    .B2(_08197_),
    .C1(net982),
    .X(_08198_));
 sky130_fd_sc_hd__o211a_1 _13514_ (.A1(\core.pipe1_resultRegister[17] ),
    .A2(net986),
    .B1(_08198_),
    .C1(net1839),
    .X(_00179_));
 sky130_fd_sc_hd__nor2_1 _13515_ (.A(_06043_),
    .B(net1116),
    .Y(_08199_));
 sky130_fd_sc_hd__a22o_1 _13516_ (.A1(\core.csr.cycleTimer.currentValue[18] ),
    .A2(net724),
    .B1(net720),
    .B2(\core.csr.cycleTimer.currentValue[50] ),
    .X(_08200_));
 sky130_fd_sc_hd__o21ai_1 _13517_ (.A1(\core.csr.cycleTimer.currentValue[18] ),
    .A2(net705),
    .B1(_07250_),
    .Y(_08201_));
 sky130_fd_sc_hd__a22o_2 _13518_ (.A1(\core.csr.instretTimer.currentValue[18] ),
    .A2(net702),
    .B1(net698),
    .B2(\core.csr.instretTimer.currentValue[50] ),
    .X(_08202_));
 sky130_fd_sc_hd__a22o_1 _13519_ (.A1(\core.csr.cycleTimer.currentValue[50] ),
    .A2(net713),
    .B1(_08202_),
    .B2(net974),
    .X(_08203_));
 sky130_fd_sc_hd__or2_1 _13520_ (.A(\core.csr.traps.mip.csrReadData[18] ),
    .B(net654),
    .X(_08204_));
 sky130_fd_sc_hd__o211a_1 _13521_ (.A1(\core.csr.traps.mtval.csrReadData[18] ),
    .A2(net662),
    .B1(net658),
    .C1(_08204_),
    .X(_08205_));
 sky130_fd_sc_hd__a21o_1 _13522_ (.A1(\core.csr.traps.mcause.csrReadData[18] ),
    .A2(net665),
    .B1(net689),
    .X(_08206_));
 sky130_fd_sc_hd__o221a_1 _13523_ (.A1(\core.csr.trapReturnVector[18] ),
    .A2(net686),
    .B1(_08205_),
    .B2(_08206_),
    .C1(net692),
    .X(_08207_));
 sky130_fd_sc_hd__a221o_1 _13524_ (.A1(\core.csr.traps.mscratch.currentValue[18] ),
    .A2(net694),
    .B1(net676),
    .B2(\core.csr.traps.mtvec.csrReadData[18] ),
    .C1(net682),
    .X(_08208_));
 sky130_fd_sc_hd__o221a_4 _13525_ (.A1(\core.csr.traps.mie.currentValue[18] ),
    .A2(net679),
    .B1(_08207_),
    .B2(_08208_),
    .C1(net607),
    .X(_08209_));
 sky130_fd_sc_hd__a2111oi_2 _13526_ (.A1(\core.csr.mconfigptr.currentValue[18] ),
    .A2(net717),
    .B1(net709),
    .C1(_08203_),
    .D1(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__a2bb2o_4 _13527_ (.A1_N(_08201_),
    .A2_N(_08210_),
    .B1(net977),
    .B2(_08200_),
    .X(_08211_));
 sky130_fd_sc_hd__a21o_1 _13528_ (.A1(net1111),
    .A2(_08211_),
    .B1(_08199_),
    .X(_08212_));
 sky130_fd_sc_hd__o21ai_1 _13529_ (.A1(net1108),
    .A2(_08199_),
    .B1(net1106),
    .Y(_08213_));
 sky130_fd_sc_hd__a32o_1 _13530_ (.A1(net1124),
    .A2(_08212_),
    .A3(_08213_),
    .B1(_06663_),
    .B2(net1153),
    .X(_08214_));
 sky130_fd_sc_hd__nand2_1 _13531_ (.A(_06663_),
    .B(net1060),
    .Y(_08215_));
 sky130_fd_sc_hd__a21boi_2 _13532_ (.A1(_06128_),
    .A2(_07333_),
    .B1_N(_07334_),
    .Y(_08216_));
 sky130_fd_sc_hd__xnor2_1 _13533_ (.A(_06051_),
    .B(_08216_),
    .Y(_08217_));
 sky130_fd_sc_hd__a21oi_1 _13534_ (.A1(net1064),
    .A2(_08217_),
    .B1(net1177),
    .Y(_08218_));
 sky130_fd_sc_hd__mux2_1 _13535_ (.A0(net1199),
    .A1(_07458_),
    .S(_06047_),
    .X(_08219_));
 sky130_fd_sc_hd__a21o_1 _13536_ (.A1(net1203),
    .A2(_08219_),
    .B1(_06049_),
    .X(_08220_));
 sky130_fd_sc_hd__o221a_1 _13537_ (.A1(net1217),
    .A2(_08042_),
    .B1(_08045_),
    .B2(net1211),
    .C1(_08220_),
    .X(_08221_));
 sky130_fd_sc_hd__a22o_1 _13538_ (.A1(_08215_),
    .A2(_08218_),
    .B1(_08221_),
    .B2(net1233),
    .X(_08222_));
 sky130_fd_sc_hd__a2bb2o_1 _13539_ (.A1_N(_08013_),
    .A2_N(_08214_),
    .B1(_08222_),
    .B2(net1119),
    .X(_08223_));
 sky130_fd_sc_hd__and2_2 _13540_ (.A(net459),
    .B(_08164_),
    .X(_08224_));
 sky130_fd_sc_hd__nor2_1 _13541_ (.A(net459),
    .B(_08164_),
    .Y(_08225_));
 sky130_fd_sc_hd__or2_1 _13542_ (.A(_08224_),
    .B(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__a22o_1 _13543_ (.A1(net1222),
    .A2(_08223_),
    .B1(_08226_),
    .B2(net1132),
    .X(_08227_));
 sky130_fd_sc_hd__nand2_1 _13544_ (.A(net1254),
    .B(_08227_),
    .Y(_08228_));
 sky130_fd_sc_hd__or2_1 _13545_ (.A(net1255),
    .B(_06663_),
    .X(_08229_));
 sky130_fd_sc_hd__a221o_4 _13546_ (.A1(\core.pipe0_currentInstruction[18] ),
    .A2(net1219),
    .B1(_08228_),
    .B2(_08229_),
    .C1(net982),
    .X(_08230_));
 sky130_fd_sc_hd__o211a_1 _13547_ (.A1(\core.pipe1_resultRegister[18] ),
    .A2(net987),
    .B1(_08230_),
    .C1(net1842),
    .X(_00180_));
 sky130_fd_sc_hd__or2_2 _13548_ (.A(_05967_),
    .B(net1116),
    .X(_08231_));
 sky130_fd_sc_hd__a22o_1 _13549_ (.A1(\core.csr.cycleTimer.currentValue[19] ),
    .A2(net724),
    .B1(net720),
    .B2(\core.csr.cycleTimer.currentValue[51] ),
    .X(_08232_));
 sky130_fd_sc_hd__a22o_2 _13550_ (.A1(\core.csr.instretTimer.currentValue[19] ),
    .A2(net702),
    .B1(net698),
    .B2(\core.csr.instretTimer.currentValue[51] ),
    .X(_08233_));
 sky130_fd_sc_hd__nor2_1 _13551_ (.A(\core.csr.cycleTimer.currentValue[19] ),
    .B(net705),
    .Y(_08234_));
 sky130_fd_sc_hd__a22o_1 _13552_ (.A1(\core.csr.cycleTimer.currentValue[51] ),
    .A2(net713),
    .B1(_08233_),
    .B2(net973),
    .X(_08235_));
 sky130_fd_sc_hd__or2_1 _13553_ (.A(\core.csr.traps.mip.csrReadData[19] ),
    .B(net654),
    .X(_08236_));
 sky130_fd_sc_hd__o211a_1 _13554_ (.A1(\core.csr.traps.mtval.csrReadData[19] ),
    .A2(net661),
    .B1(net658),
    .C1(_08236_),
    .X(_08237_));
 sky130_fd_sc_hd__a21o_1 _13555_ (.A1(\core.csr.traps.mcause.csrReadData[19] ),
    .A2(net664),
    .B1(net688),
    .X(_08238_));
 sky130_fd_sc_hd__o221a_1 _13556_ (.A1(\core.csr.trapReturnVector[19] ),
    .A2(net685),
    .B1(_08237_),
    .B2(_08238_),
    .C1(net691),
    .X(_08239_));
 sky130_fd_sc_hd__a221o_1 _13557_ (.A1(\core.csr.traps.mscratch.currentValue[19] ),
    .A2(net694),
    .B1(net676),
    .B2(\core.csr.traps.mtvec.csrReadData[19] ),
    .C1(net682),
    .X(_08240_));
 sky130_fd_sc_hd__o221a_4 _13558_ (.A1(\core.csr.traps.mie.currentValue[19] ),
    .A2(net679),
    .B1(_08239_),
    .B2(_08240_),
    .C1(net607),
    .X(_08241_));
 sky130_fd_sc_hd__a2111oi_2 _13559_ (.A1(\core.csr.mconfigptr.currentValue[19] ),
    .A2(net717),
    .B1(net709),
    .C1(_08235_),
    .D1(_08241_),
    .Y(_08242_));
 sky130_fd_sc_hd__o2bb2a_4 _13560_ (.A1_N(net973),
    .A2_N(_08232_),
    .B1(_08234_),
    .B2(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__inv_2 _13561_ (.A(_08243_),
    .Y(_08244_));
 sky130_fd_sc_hd__o21ai_1 _13562_ (.A1(net1112),
    .A2(_08243_),
    .B1(_08231_),
    .Y(_08245_));
 sky130_fd_sc_hd__a21o_1 _13563_ (.A1(net1109),
    .A2(_08231_),
    .B1(net1105),
    .X(_08246_));
 sky130_fd_sc_hd__a311o_2 _13564_ (.A1(net1122),
    .A2(_08245_),
    .A3(_08246_),
    .B1(_07147_),
    .C1(net1185),
    .X(_08247_));
 sky130_fd_sc_hd__a21oi_1 _13565_ (.A1(net1153),
    .A2(_06662_),
    .B1(_08247_),
    .Y(_08248_));
 sky130_fd_sc_hd__nand2_1 _13566_ (.A(_06662_),
    .B(net1060),
    .Y(_08249_));
 sky130_fd_sc_hd__o21ai_2 _13567_ (.A1(_06050_),
    .A2(_08216_),
    .B1(_07296_),
    .Y(_08250_));
 sky130_fd_sc_hd__xnor2_2 _13568_ (.A(_06661_),
    .B(_08250_),
    .Y(_08251_));
 sky130_fd_sc_hd__a21oi_1 _13569_ (.A1(net1063),
    .A2(_08251_),
    .B1(net1177),
    .Y(_08252_));
 sky130_fd_sc_hd__a221o_1 _13570_ (.A1(_05973_),
    .A2(net1205),
    .B1(net1201),
    .B2(_05971_),
    .C1(net1274),
    .X(_08253_));
 sky130_fd_sc_hd__a21oi_1 _13571_ (.A1(_06644_),
    .A2(_06661_),
    .B1(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__o22a_1 _13572_ (.A1(net1217),
    .A2(_08003_),
    .B1(_08005_),
    .B2(net1210),
    .X(_08255_));
 sky130_fd_sc_hd__a22o_1 _13573_ (.A1(_08249_),
    .A2(_08252_),
    .B1(_08254_),
    .B2(_08255_),
    .X(_08256_));
 sky130_fd_sc_hd__a21o_1 _13574_ (.A1(net1119),
    .A2(_08256_),
    .B1(_08248_),
    .X(_08257_));
 sky130_fd_sc_hd__xnor2_2 _13575_ (.A(net460),
    .B(_08224_),
    .Y(_08258_));
 sky130_fd_sc_hd__inv_2 _13576_ (.A(_08258_),
    .Y(_08259_));
 sky130_fd_sc_hd__a22o_1 _13577_ (.A1(net1222),
    .A2(_08257_),
    .B1(_08258_),
    .B2(net1135),
    .X(_08260_));
 sky130_fd_sc_hd__a22o_1 _13578_ (.A1(net1264),
    .A2(_06662_),
    .B1(net1219),
    .B2(net1780),
    .X(_08261_));
 sky130_fd_sc_hd__or3b_4 _13579_ (.A(net982),
    .B(_08261_),
    .C_N(_08260_),
    .X(_08262_));
 sky130_fd_sc_hd__o211a_1 _13580_ (.A1(\core.pipe1_resultRegister[19] ),
    .A2(net986),
    .B1(_08262_),
    .C1(net1839),
    .X(_00181_));
 sky130_fd_sc_hd__or2_1 _13581_ (.A(_05891_),
    .B(net1116),
    .X(_08263_));
 sky130_fd_sc_hd__a22o_1 _13582_ (.A1(\core.csr.cycleTimer.currentValue[20] ),
    .A2(net724),
    .B1(net720),
    .B2(\core.csr.cycleTimer.currentValue[52] ),
    .X(_08264_));
 sky130_fd_sc_hd__o21ai_1 _13583_ (.A1(\core.csr.cycleTimer.currentValue[20] ),
    .A2(net705),
    .B1(_07250_),
    .Y(_08265_));
 sky130_fd_sc_hd__a22o_2 _13584_ (.A1(\core.csr.instretTimer.currentValue[20] ),
    .A2(net702),
    .B1(net698),
    .B2(\core.csr.instretTimer.currentValue[52] ),
    .X(_08266_));
 sky130_fd_sc_hd__a22o_1 _13585_ (.A1(\core.csr.cycleTimer.currentValue[52] ),
    .A2(net713),
    .B1(_08266_),
    .B2(net973),
    .X(_08267_));
 sky130_fd_sc_hd__or2_1 _13586_ (.A(\core.csr.traps.mip.csrReadData[20] ),
    .B(net654),
    .X(_08268_));
 sky130_fd_sc_hd__o211a_1 _13587_ (.A1(\core.csr.traps.mtval.csrReadData[20] ),
    .A2(net661),
    .B1(net658),
    .C1(_08268_),
    .X(_08269_));
 sky130_fd_sc_hd__a21o_1 _13588_ (.A1(\core.csr.traps.mcause.csrReadData[20] ),
    .A2(net664),
    .B1(net688),
    .X(_08270_));
 sky130_fd_sc_hd__o221a_1 _13589_ (.A1(\core.csr.trapReturnVector[20] ),
    .A2(net685),
    .B1(_08269_),
    .B2(_08270_),
    .C1(net691),
    .X(_08271_));
 sky130_fd_sc_hd__a221o_1 _13590_ (.A1(\core.csr.traps.mscratch.currentValue[20] ),
    .A2(net694),
    .B1(net676),
    .B2(\core.csr.traps.mtvec.csrReadData[20] ),
    .C1(net682),
    .X(_08272_));
 sky130_fd_sc_hd__o221a_4 _13591_ (.A1(\core.csr.traps.mie.currentValue[20] ),
    .A2(net679),
    .B1(_08271_),
    .B2(_08272_),
    .C1(net607),
    .X(_08273_));
 sky130_fd_sc_hd__a2111oi_2 _13592_ (.A1(\core.csr.mconfigptr.currentValue[20] ),
    .A2(net718),
    .B1(net709),
    .C1(_08267_),
    .D1(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__o2bb2a_4 _13593_ (.A1_N(net973),
    .A2_N(_08264_),
    .B1(_08265_),
    .B2(_08274_),
    .X(_08275_));
 sky130_fd_sc_hd__inv_2 _13594_ (.A(_08275_),
    .Y(_08276_));
 sky130_fd_sc_hd__o21ai_1 _13595_ (.A1(net1113),
    .A2(_08275_),
    .B1(_08263_),
    .Y(_08277_));
 sky130_fd_sc_hd__a21o_1 _13596_ (.A1(net1110),
    .A2(_08263_),
    .B1(net1104),
    .X(_08278_));
 sky130_fd_sc_hd__xnor2_1 _13597_ (.A(_05897_),
    .B(_07338_),
    .Y(_08279_));
 sky130_fd_sc_hd__a21o_1 _13598_ (.A1(net1063),
    .A2(_08279_),
    .B1(net1177),
    .X(_08280_));
 sky130_fd_sc_hd__a21oi_1 _13599_ (.A1(_06660_),
    .A2(net1060),
    .B1(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__mux2_1 _13600_ (.A0(net1199),
    .A1(_07458_),
    .S(_05895_),
    .X(_08282_));
 sky130_fd_sc_hd__a21o_1 _13601_ (.A1(net1203),
    .A2(_08282_),
    .B1(_05896_),
    .X(_08283_));
 sky130_fd_sc_hd__o2bb2a_1 _13602_ (.A1_N(net1213),
    .A2_N(_07956_),
    .B1(_07957_),
    .B2(net1217),
    .X(_08284_));
 sky130_fd_sc_hd__a31o_1 _13603_ (.A1(net1233),
    .A2(_08283_),
    .A3(_08284_),
    .B1(_08281_),
    .X(_08285_));
 sky130_fd_sc_hd__a32o_1 _13604_ (.A1(net1124),
    .A2(_08277_),
    .A3(_08278_),
    .B1(_06660_),
    .B2(net1153),
    .X(_08286_));
 sky130_fd_sc_hd__o2bb2a_1 _13605_ (.A1_N(net1118),
    .A2_N(_08285_),
    .B1(_08286_),
    .B2(_08013_),
    .X(_08287_));
 sky130_fd_sc_hd__and3_1 _13606_ (.A(net462),
    .B(net460),
    .C(_08224_),
    .X(_08288_));
 sky130_fd_sc_hd__a21oi_1 _13607_ (.A1(net460),
    .A2(_08224_),
    .B1(net462),
    .Y(_08289_));
 sky130_fd_sc_hd__or2_1 _13608_ (.A(_08288_),
    .B(_08289_),
    .X(_08290_));
 sky130_fd_sc_hd__a2bb2o_1 _13609_ (.A1_N(net1228),
    .A2_N(_08287_),
    .B1(_08290_),
    .B2(net1132),
    .X(_08291_));
 sky130_fd_sc_hd__nand2_1 _13610_ (.A(net1254),
    .B(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__or2_1 _13611_ (.A(net1254),
    .B(_06660_),
    .X(_08293_));
 sky130_fd_sc_hd__a221o_4 _13612_ (.A1(net1776),
    .A2(net1219),
    .B1(_08292_),
    .B2(_08293_),
    .C1(net982),
    .X(_08294_));
 sky130_fd_sc_hd__o211a_1 _13613_ (.A1(\core.pipe1_resultRegister[20] ),
    .A2(net986),
    .B1(_08294_),
    .C1(net1839),
    .X(_00182_));
 sky130_fd_sc_hd__nand2_1 _13614_ (.A(_06659_),
    .B(net1060),
    .Y(_08295_));
 sky130_fd_sc_hd__nand2_1 _13615_ (.A(_07339_),
    .B(_07343_),
    .Y(_08296_));
 sky130_fd_sc_hd__xnor2_1 _13616_ (.A(_06525_),
    .B(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__a21oi_1 _13617_ (.A1(net1062),
    .A2(_08297_),
    .B1(net1177),
    .Y(_08298_));
 sky130_fd_sc_hd__a221o_1 _13618_ (.A1(_05818_),
    .A2(net1205),
    .B1(net1201),
    .B2(_05820_),
    .C1(net1274),
    .X(_08299_));
 sky130_fd_sc_hd__a21oi_1 _13619_ (.A1(_06525_),
    .A2(_06644_),
    .B1(_08299_),
    .Y(_08300_));
 sky130_fd_sc_hd__o22a_1 _13620_ (.A1(net1207),
    .A2(_07921_),
    .B1(_07924_),
    .B2(net1216),
    .X(_08301_));
 sky130_fd_sc_hd__a22o_1 _13621_ (.A1(_08295_),
    .A2(_08298_),
    .B1(_08300_),
    .B2(_08301_),
    .X(_08302_));
 sky130_fd_sc_hd__nand2_1 _13622_ (.A(net1153),
    .B(_06659_),
    .Y(_08303_));
 sky130_fd_sc_hd__or2_1 _13623_ (.A(_05815_),
    .B(net1116),
    .X(_08304_));
 sky130_fd_sc_hd__a22o_1 _13624_ (.A1(\core.csr.cycleTimer.currentValue[21] ),
    .A2(net724),
    .B1(net720),
    .B2(\core.csr.cycleTimer.currentValue[53] ),
    .X(_08305_));
 sky130_fd_sc_hd__a22o_2 _13625_ (.A1(\core.csr.instretTimer.currentValue[21] ),
    .A2(net702),
    .B1(net698),
    .B2(\core.csr.instretTimer.currentValue[53] ),
    .X(_08306_));
 sky130_fd_sc_hd__nor2_1 _13626_ (.A(\core.csr.cycleTimer.currentValue[21] ),
    .B(net705),
    .Y(_08307_));
 sky130_fd_sc_hd__a22o_1 _13627_ (.A1(\core.csr.cycleTimer.currentValue[53] ),
    .A2(net713),
    .B1(_08306_),
    .B2(net973),
    .X(_08308_));
 sky130_fd_sc_hd__or2_1 _13628_ (.A(\core.csr.traps.mip.csrReadData[21] ),
    .B(net655),
    .X(_08309_));
 sky130_fd_sc_hd__o211a_1 _13629_ (.A1(\core.csr.traps.mtval.csrReadData[21] ),
    .A2(net662),
    .B1(net659),
    .C1(_08309_),
    .X(_08310_));
 sky130_fd_sc_hd__a21o_1 _13630_ (.A1(\core.csr.traps.mcause.csrReadData[21] ),
    .A2(net665),
    .B1(net689),
    .X(_08311_));
 sky130_fd_sc_hd__o221a_1 _13631_ (.A1(\core.csr.trapReturnVector[21] ),
    .A2(net686),
    .B1(_08310_),
    .B2(_08311_),
    .C1(net692),
    .X(_08312_));
 sky130_fd_sc_hd__a221o_1 _13632_ (.A1(\core.csr.traps.mscratch.currentValue[21] ),
    .A2(net695),
    .B1(net677),
    .B2(\core.csr.traps.mtvec.csrReadData[21] ),
    .C1(net683),
    .X(_08313_));
 sky130_fd_sc_hd__o221a_4 _13633_ (.A1(\core.csr.traps.mie.currentValue[21] ),
    .A2(net680),
    .B1(_08312_),
    .B2(_08313_),
    .C1(net608),
    .X(_08314_));
 sky130_fd_sc_hd__a2111oi_2 _13634_ (.A1(\core.csr.mconfigptr.currentValue[21] ),
    .A2(net717),
    .B1(net709),
    .C1(_08308_),
    .D1(_08314_),
    .Y(_08315_));
 sky130_fd_sc_hd__o2bb2a_4 _13635_ (.A1_N(net973),
    .A2_N(_08305_),
    .B1(_08307_),
    .B2(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__inv_2 _13636_ (.A(_08316_),
    .Y(_08317_));
 sky130_fd_sc_hd__or2_4 _13637_ (.A(net1113),
    .B(_08316_),
    .X(_08318_));
 sky130_fd_sc_hd__nand2_1 _13638_ (.A(net1110),
    .B(_08304_),
    .Y(_08319_));
 sky130_fd_sc_hd__a221o_1 _13639_ (.A1(_08304_),
    .A2(_08318_),
    .B1(_08319_),
    .B2(net1106),
    .C1(net1120),
    .X(_08320_));
 sky130_fd_sc_hd__a32o_2 _13640_ (.A1(net1059),
    .A2(_08303_),
    .A3(_08320_),
    .B1(_08302_),
    .B2(net1118),
    .X(_08321_));
 sky130_fd_sc_hd__and2_2 _13641_ (.A(net463),
    .B(_08288_),
    .X(_08322_));
 sky130_fd_sc_hd__nor2_1 _13642_ (.A(net463),
    .B(_08288_),
    .Y(_08323_));
 sky130_fd_sc_hd__or2_2 _13643_ (.A(_08322_),
    .B(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__a22oi_4 _13644_ (.A1(net1221),
    .A2(_08321_),
    .B1(_08324_),
    .B2(net1132),
    .Y(_08325_));
 sky130_fd_sc_hd__a221o_1 _13645_ (.A1(net1264),
    .A2(_06659_),
    .B1(net1219),
    .B2(net1771),
    .C1(net982),
    .X(_08326_));
 sky130_fd_sc_hd__o221a_1 _13646_ (.A1(\core.pipe1_resultRegister[21] ),
    .A2(net988),
    .B1(_08325_),
    .B2(_08326_),
    .C1(net1824),
    .X(_00183_));
 sky130_fd_sc_hd__nor2_1 _13647_ (.A(_05737_),
    .B(net1116),
    .Y(_08327_));
 sky130_fd_sc_hd__a22o_1 _13648_ (.A1(\core.csr.cycleTimer.currentValue[22] ),
    .A2(net724),
    .B1(net720),
    .B2(\core.csr.cycleTimer.currentValue[54] ),
    .X(_08328_));
 sky130_fd_sc_hd__o21ai_1 _13649_ (.A1(\core.csr.cycleTimer.currentValue[22] ),
    .A2(net705),
    .B1(_07250_),
    .Y(_08329_));
 sky130_fd_sc_hd__a22o_2 _13650_ (.A1(\core.csr.instretTimer.currentValue[22] ),
    .A2(net701),
    .B1(net697),
    .B2(\core.csr.instretTimer.currentValue[54] ),
    .X(_08330_));
 sky130_fd_sc_hd__a22o_1 _13651_ (.A1(\core.csr.cycleTimer.currentValue[54] ),
    .A2(net713),
    .B1(_08330_),
    .B2(net973),
    .X(_08331_));
 sky130_fd_sc_hd__or2_1 _13652_ (.A(\core.csr.traps.mip.csrReadData[22] ),
    .B(net655),
    .X(_08332_));
 sky130_fd_sc_hd__o211a_1 _13653_ (.A1(\core.csr.traps.mtval.csrReadData[22] ),
    .A2(net661),
    .B1(net659),
    .C1(_08332_),
    .X(_08333_));
 sky130_fd_sc_hd__a21o_1 _13654_ (.A1(\core.csr.traps.mcause.csrReadData[22] ),
    .A2(net665),
    .B1(net689),
    .X(_08334_));
 sky130_fd_sc_hd__o221a_1 _13655_ (.A1(\core.csr.trapReturnVector[22] ),
    .A2(net686),
    .B1(_08333_),
    .B2(_08334_),
    .C1(net692),
    .X(_08335_));
 sky130_fd_sc_hd__a221o_1 _13656_ (.A1(\core.csr.traps.mscratch.currentValue[22] ),
    .A2(net695),
    .B1(net677),
    .B2(\core.csr.traps.mtvec.csrReadData[22] ),
    .C1(net683),
    .X(_08336_));
 sky130_fd_sc_hd__o221a_4 _13657_ (.A1(\core.csr.traps.mie.currentValue[22] ),
    .A2(net680),
    .B1(_08335_),
    .B2(_08336_),
    .C1(net608),
    .X(_08337_));
 sky130_fd_sc_hd__a2111oi_2 _13658_ (.A1(\core.csr.mconfigptr.currentValue[22] ),
    .A2(net717),
    .B1(net709),
    .C1(_08331_),
    .D1(_08337_),
    .Y(_08338_));
 sky130_fd_sc_hd__a2bb2o_4 _13659_ (.A1_N(_08329_),
    .A2_N(_08338_),
    .B1(net973),
    .B2(_08328_),
    .X(_08339_));
 sky130_fd_sc_hd__a21oi_1 _13660_ (.A1(net1111),
    .A2(_08339_),
    .B1(_08327_),
    .Y(_08340_));
 sky130_fd_sc_hd__o21a_1 _13661_ (.A1(net1108),
    .A2(_08327_),
    .B1(net1106),
    .X(_08341_));
 sky130_fd_sc_hd__o32a_1 _13662_ (.A1(net1120),
    .A2(_08340_),
    .A3(_08341_),
    .B1(_06657_),
    .B2(net1150),
    .X(_08342_));
 sky130_fd_sc_hd__or2_1 _13663_ (.A(_06657_),
    .B(net1062),
    .X(_08343_));
 sky130_fd_sc_hd__o21ba_2 _13664_ (.A1(_06525_),
    .A2(_07339_),
    .B1_N(_07344_),
    .X(_08344_));
 sky130_fd_sc_hd__xnor2_2 _13665_ (.A(_05743_),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__nand2_1 _13666_ (.A(net1062),
    .B(_08345_),
    .Y(_08346_));
 sky130_fd_sc_hd__a21oi_1 _13667_ (.A1(_05740_),
    .A2(net1201),
    .B1(net1205),
    .Y(_08347_));
 sky130_fd_sc_hd__o22a_1 _13668_ (.A1(_05743_),
    .A2(net1199),
    .B1(_08347_),
    .B2(_05741_),
    .X(_08348_));
 sky130_fd_sc_hd__o211a_1 _13669_ (.A1(net1215),
    .A2(_07890_),
    .B1(_08348_),
    .C1(net1233),
    .X(_08349_));
 sky130_fd_sc_hd__o21a_1 _13670_ (.A1(net1209),
    .A2(_07887_),
    .B1(_08349_),
    .X(_08350_));
 sky130_fd_sc_hd__a31o_1 _13671_ (.A1(_07950_),
    .A2(_08343_),
    .A3(_08346_),
    .B1(_08350_),
    .X(_08351_));
 sky130_fd_sc_hd__a22o_1 _13672_ (.A1(net1059),
    .A2(_08342_),
    .B1(_08351_),
    .B2(net1118),
    .X(_08352_));
 sky130_fd_sc_hd__xnor2_1 _13673_ (.A(net464),
    .B(_08322_),
    .Y(_08353_));
 sky130_fd_sc_hd__a22o_1 _13674_ (.A1(net1221),
    .A2(_08352_),
    .B1(_08353_),
    .B2(net1132),
    .X(_08354_));
 sky130_fd_sc_hd__nand2_2 _13675_ (.A(net1251),
    .B(_08354_),
    .Y(_08355_));
 sky130_fd_sc_hd__nand2_1 _13676_ (.A(net1264),
    .B(_06657_),
    .Y(_08356_));
 sky130_fd_sc_hd__a221o_4 _13677_ (.A1(net1764),
    .A2(net1219),
    .B1(_08355_),
    .B2(_08356_),
    .C1(net982),
    .X(_08357_));
 sky130_fd_sc_hd__o211a_1 _13678_ (.A1(\core.pipe1_resultRegister[22] ),
    .A2(net988),
    .B1(_08357_),
    .C1(net1837),
    .X(_00184_));
 sky130_fd_sc_hd__nor2_1 _13679_ (.A(_05661_),
    .B(net1116),
    .Y(_08358_));
 sky130_fd_sc_hd__a22o_1 _13680_ (.A1(\core.csr.cycleTimer.currentValue[23] ),
    .A2(net724),
    .B1(net720),
    .B2(\core.csr.cycleTimer.currentValue[55] ),
    .X(_08359_));
 sky130_fd_sc_hd__a22o_2 _13681_ (.A1(\core.csr.instretTimer.currentValue[23] ),
    .A2(net701),
    .B1(net697),
    .B2(\core.csr.instretTimer.currentValue[55] ),
    .X(_08360_));
 sky130_fd_sc_hd__a22o_1 _13682_ (.A1(\core.csr.cycleTimer.currentValue[55] ),
    .A2(net713),
    .B1(_08360_),
    .B2(net973),
    .X(_08361_));
 sky130_fd_sc_hd__a211o_1 _13683_ (.A1(\core.csr.mconfigptr.currentValue[23] ),
    .A2(net717),
    .B1(net709),
    .C1(_08361_),
    .X(_08362_));
 sky130_fd_sc_hd__or2_1 _13684_ (.A(\core.csr.traps.mip.csrReadData[23] ),
    .B(net654),
    .X(_08363_));
 sky130_fd_sc_hd__o211a_1 _13685_ (.A1(\core.csr.traps.mtval.csrReadData[23] ),
    .A2(net661),
    .B1(net658),
    .C1(_08363_),
    .X(_08364_));
 sky130_fd_sc_hd__a21o_1 _13686_ (.A1(\core.csr.traps.mcause.csrReadData[23] ),
    .A2(net664),
    .B1(net688),
    .X(_08365_));
 sky130_fd_sc_hd__o221a_1 _13687_ (.A1(\core.csr.trapReturnVector[23] ),
    .A2(net685),
    .B1(_08364_),
    .B2(_08365_),
    .C1(net691),
    .X(_08366_));
 sky130_fd_sc_hd__a221o_1 _13688_ (.A1(\core.csr.traps.mscratch.currentValue[23] ),
    .A2(net694),
    .B1(net676),
    .B2(\core.csr.traps.mtvec.csrReadData[23] ),
    .C1(net682),
    .X(_08367_));
 sky130_fd_sc_hd__o221a_4 _13689_ (.A1(\core.csr.traps.mie.currentValue[23] ),
    .A2(net679),
    .B1(_08366_),
    .B2(_08367_),
    .C1(net607),
    .X(_08368_));
 sky130_fd_sc_hd__o22a_1 _13690_ (.A1(\core.csr.cycleTimer.currentValue[23] ),
    .A2(net705),
    .B1(_08362_),
    .B2(_08368_),
    .X(_08369_));
 sky130_fd_sc_hd__a21o_4 _13691_ (.A1(net974),
    .A2(_08359_),
    .B1(_08369_),
    .X(_08370_));
 sky130_fd_sc_hd__a21oi_1 _13692_ (.A1(net1111),
    .A2(_08370_),
    .B1(_08358_),
    .Y(_08371_));
 sky130_fd_sc_hd__o21a_1 _13693_ (.A1(net1108),
    .A2(_08358_),
    .B1(net1106),
    .X(_08372_));
 sky130_fd_sc_hd__o32a_1 _13694_ (.A1(net1120),
    .A2(_08371_),
    .A3(_08372_),
    .B1(_06655_),
    .B2(net1150),
    .X(_08373_));
 sky130_fd_sc_hd__or2_1 _13695_ (.A(_06655_),
    .B(net1062),
    .X(_08374_));
 sky130_fd_sc_hd__o21ai_4 _13696_ (.A1(_05742_),
    .A2(_08344_),
    .B1(_07341_),
    .Y(_08375_));
 sky130_fd_sc_hd__xnor2_4 _13697_ (.A(_06529_),
    .B(_08375_),
    .Y(_08376_));
 sky130_fd_sc_hd__nand2_1 _13698_ (.A(net1062),
    .B(_08376_),
    .Y(_08377_));
 sky130_fd_sc_hd__a221oi_2 _13699_ (.A1(_05664_),
    .A2(net1201),
    .B1(_07537_),
    .B2(_06529_),
    .C1(net1274),
    .Y(_08378_));
 sky130_fd_sc_hd__o221a_1 _13700_ (.A1(_05665_),
    .A2(net1203),
    .B1(_07847_),
    .B2(net1207),
    .C1(_08378_),
    .X(_08379_));
 sky130_fd_sc_hd__o21a_1 _13701_ (.A1(net1215),
    .A2(_07850_),
    .B1(_08379_),
    .X(_08380_));
 sky130_fd_sc_hd__a31o_1 _13702_ (.A1(_07950_),
    .A2(_08374_),
    .A3(_08377_),
    .B1(_08380_),
    .X(_08381_));
 sky130_fd_sc_hd__a22o_1 _13703_ (.A1(net1059),
    .A2(_08373_),
    .B1(_08381_),
    .B2(net1118),
    .X(_08382_));
 sky130_fd_sc_hd__and3_1 _13704_ (.A(net465),
    .B(net464),
    .C(_08322_),
    .X(_08383_));
 sky130_fd_sc_hd__a21oi_1 _13705_ (.A1(net464),
    .A2(_08322_),
    .B1(net465),
    .Y(_08384_));
 sky130_fd_sc_hd__or2_1 _13706_ (.A(_08383_),
    .B(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__a22o_1 _13707_ (.A1(net1221),
    .A2(_08382_),
    .B1(_08385_),
    .B2(net1132),
    .X(_08386_));
 sky130_fd_sc_hd__o21ai_4 _13708_ (.A1(net1251),
    .A2(_06655_),
    .B1(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__a211o_4 _13709_ (.A1(net1762),
    .A2(_07141_),
    .B1(net985),
    .C1(_08387_),
    .X(_08388_));
 sky130_fd_sc_hd__o211a_1 _13710_ (.A1(\core.pipe1_resultRegister[23] ),
    .A2(net986),
    .B1(_08388_),
    .C1(net1837),
    .X(_00185_));
 sky130_fd_sc_hd__nor2_1 _13711_ (.A(_05586_),
    .B(net1116),
    .Y(_08389_));
 sky130_fd_sc_hd__a22o_1 _13712_ (.A1(\core.csr.cycleTimer.currentValue[24] ),
    .A2(net724),
    .B1(net720),
    .B2(\core.csr.cycleTimer.currentValue[56] ),
    .X(_08390_));
 sky130_fd_sc_hd__o21ai_1 _13713_ (.A1(\core.csr.cycleTimer.currentValue[24] ),
    .A2(net705),
    .B1(_07250_),
    .Y(_08391_));
 sky130_fd_sc_hd__a22o_1 _13714_ (.A1(\core.csr.instretTimer.currentValue[24] ),
    .A2(net701),
    .B1(net697),
    .B2(\core.csr.instretTimer.currentValue[56] ),
    .X(_08392_));
 sky130_fd_sc_hd__a22o_1 _13715_ (.A1(\core.csr.cycleTimer.currentValue[56] ),
    .A2(net713),
    .B1(_08392_),
    .B2(net974),
    .X(_08393_));
 sky130_fd_sc_hd__or2_1 _13716_ (.A(\core.csr.traps.mip.csrReadData[24] ),
    .B(net655),
    .X(_08394_));
 sky130_fd_sc_hd__o211a_1 _13717_ (.A1(\core.csr.traps.mtval.csrReadData[24] ),
    .A2(net661),
    .B1(net659),
    .C1(_08394_),
    .X(_08395_));
 sky130_fd_sc_hd__a21o_1 _13718_ (.A1(\core.csr.traps.mcause.csrReadData[24] ),
    .A2(net664),
    .B1(net688),
    .X(_08396_));
 sky130_fd_sc_hd__o221a_2 _13719_ (.A1(\core.csr.trapReturnVector[24] ),
    .A2(net685),
    .B1(_08395_),
    .B2(_08396_),
    .C1(net691),
    .X(_08397_));
 sky130_fd_sc_hd__a221o_1 _13720_ (.A1(\core.csr.traps.mscratch.currentValue[24] ),
    .A2(net694),
    .B1(net676),
    .B2(\core.csr.traps.mtvec.csrReadData[24] ),
    .C1(net682),
    .X(_08398_));
 sky130_fd_sc_hd__o221a_4 _13721_ (.A1(\core.csr.traps.mie.currentValue[24] ),
    .A2(net679),
    .B1(_08397_),
    .B2(_08398_),
    .C1(net607),
    .X(_08399_));
 sky130_fd_sc_hd__a2111oi_2 _13722_ (.A1(\core.csr.mconfigptr.currentValue[24] ),
    .A2(net718),
    .B1(net709),
    .C1(_08393_),
    .D1(_08399_),
    .Y(_08400_));
 sky130_fd_sc_hd__a2bb2o_4 _13723_ (.A1_N(_08391_),
    .A2_N(_08400_),
    .B1(net974),
    .B2(_08390_),
    .X(_08401_));
 sky130_fd_sc_hd__a21oi_1 _13724_ (.A1(net1111),
    .A2(_08401_),
    .B1(_08389_),
    .Y(_08402_));
 sky130_fd_sc_hd__o21a_1 _13725_ (.A1(net1108),
    .A2(_08389_),
    .B1(net1106),
    .X(_08403_));
 sky130_fd_sc_hd__o32a_1 _13726_ (.A1(net1120),
    .A2(_08402_),
    .A3(_08403_),
    .B1(_06630_),
    .B2(net1150),
    .X(_08404_));
 sky130_fd_sc_hd__xnor2_2 _13727_ (.A(_05591_),
    .B(_07348_),
    .Y(_08405_));
 sky130_fd_sc_hd__a21oi_1 _13728_ (.A1(net1062),
    .A2(_08405_),
    .B1(net1177),
    .Y(_08406_));
 sky130_fd_sc_hd__o21a_1 _13729_ (.A1(_06630_),
    .A2(net1062),
    .B1(_08406_),
    .X(_08407_));
 sky130_fd_sc_hd__a21oi_1 _13730_ (.A1(_05589_),
    .A2(net1201),
    .B1(net1205),
    .Y(_08408_));
 sky130_fd_sc_hd__o22a_1 _13731_ (.A1(_05592_),
    .A2(net1199),
    .B1(_08408_),
    .B2(_05590_),
    .X(_08409_));
 sky130_fd_sc_hd__o22a_1 _13732_ (.A1(net1207),
    .A2(_07832_),
    .B1(_07835_),
    .B2(net1215),
    .X(_08410_));
 sky130_fd_sc_hd__a31o_1 _13733_ (.A1(net1233),
    .A2(_08409_),
    .A3(_08410_),
    .B1(_08407_),
    .X(_08411_));
 sky130_fd_sc_hd__a22o_1 _13734_ (.A1(net1059),
    .A2(_08404_),
    .B1(_08411_),
    .B2(net1118),
    .X(_08412_));
 sky130_fd_sc_hd__and2_1 _13735_ (.A(net466),
    .B(_08383_),
    .X(_08413_));
 sky130_fd_sc_hd__nor2_1 _13736_ (.A(net466),
    .B(_08383_),
    .Y(_08414_));
 sky130_fd_sc_hd__or2_1 _13737_ (.A(_08413_),
    .B(_08414_),
    .X(_08415_));
 sky130_fd_sc_hd__a22o_1 _13738_ (.A1(net1221),
    .A2(_08412_),
    .B1(_08415_),
    .B2(net1132),
    .X(_08416_));
 sky130_fd_sc_hd__nand2_2 _13739_ (.A(net1251),
    .B(_08416_),
    .Y(_08417_));
 sky130_fd_sc_hd__nand2_1 _13740_ (.A(net1264),
    .B(_06630_),
    .Y(_08418_));
 sky130_fd_sc_hd__a221o_4 _13741_ (.A1(net1754),
    .A2(net1219),
    .B1(_08417_),
    .B2(_08418_),
    .C1(net982),
    .X(_08419_));
 sky130_fd_sc_hd__o211a_1 _13742_ (.A1(\core.pipe1_resultRegister[24] ),
    .A2(net986),
    .B1(_08419_),
    .C1(net1840),
    .X(_00186_));
 sky130_fd_sc_hd__or2_1 _13743_ (.A(_05511_),
    .B(net1116),
    .X(_08420_));
 sky130_fd_sc_hd__a22o_1 _13744_ (.A1(\core.csr.cycleTimer.currentValue[25] ),
    .A2(net724),
    .B1(net720),
    .B2(\core.csr.cycleTimer.currentValue[57] ),
    .X(_08421_));
 sky130_fd_sc_hd__a22o_1 _13745_ (.A1(\core.csr.instretTimer.currentValue[25] ),
    .A2(net701),
    .B1(net697),
    .B2(\core.csr.instretTimer.currentValue[57] ),
    .X(_08422_));
 sky130_fd_sc_hd__nor2_1 _13746_ (.A(\core.csr.cycleTimer.currentValue[25] ),
    .B(net706),
    .Y(_08423_));
 sky130_fd_sc_hd__a221o_1 _13747_ (.A1(\core.csr.cycleTimer.currentValue[57] ),
    .A2(net713),
    .B1(_08422_),
    .B2(net974),
    .C1(net710),
    .X(_08424_));
 sky130_fd_sc_hd__or2_1 _13748_ (.A(\core.csr.traps.mip.csrReadData[25] ),
    .B(net654),
    .X(_08425_));
 sky130_fd_sc_hd__o211a_1 _13749_ (.A1(\core.csr.traps.mtval.csrReadData[25] ),
    .A2(net661),
    .B1(net658),
    .C1(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__a21o_1 _13750_ (.A1(\core.csr.traps.mcause.csrReadData[25] ),
    .A2(net664),
    .B1(net688),
    .X(_08427_));
 sky130_fd_sc_hd__o221a_1 _13751_ (.A1(\core.csr.trapReturnVector[25] ),
    .A2(net685),
    .B1(_08426_),
    .B2(_08427_),
    .C1(net691),
    .X(_08428_));
 sky130_fd_sc_hd__a221o_1 _13752_ (.A1(\core.csr.traps.mscratch.currentValue[25] ),
    .A2(net694),
    .B1(net676),
    .B2(\core.csr.traps.mtvec.csrReadData[25] ),
    .C1(net682),
    .X(_08429_));
 sky130_fd_sc_hd__o221a_4 _13753_ (.A1(\core.csr.traps.mie.currentValue[25] ),
    .A2(net679),
    .B1(_08428_),
    .B2(_08429_),
    .C1(net607),
    .X(_08430_));
 sky130_fd_sc_hd__a211oi_2 _13754_ (.A1(\core.csr.mconfigptr.currentValue[25] ),
    .A2(net718),
    .B1(_08424_),
    .C1(_08430_),
    .Y(_08431_));
 sky130_fd_sc_hd__o2bb2a_4 _13755_ (.A1_N(net974),
    .A2_N(_08421_),
    .B1(_08423_),
    .B2(_08431_),
    .X(_08432_));
 sky130_fd_sc_hd__inv_2 _13756_ (.A(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__or2_4 _13757_ (.A(net1112),
    .B(_08432_),
    .X(_08434_));
 sky130_fd_sc_hd__nand2_1 _13758_ (.A(net1110),
    .B(_08420_),
    .Y(_08435_));
 sky130_fd_sc_hd__a221o_1 _13759_ (.A1(_08420_),
    .A2(_08434_),
    .B1(_08435_),
    .B2(net1106),
    .C1(net1120),
    .X(_08436_));
 sky130_fd_sc_hd__o211a_1 _13760_ (.A1(net1150),
    .A2(_06628_),
    .B1(net1059),
    .C1(_08436_),
    .X(_08437_));
 sky130_fd_sc_hd__or2_1 _13761_ (.A(_06628_),
    .B(net1062),
    .X(_08438_));
 sky130_fd_sc_hd__a21oi_2 _13762_ (.A1(_05592_),
    .A2(_07348_),
    .B1(_07352_),
    .Y(_08439_));
 sky130_fd_sc_hd__xnor2_2 _13763_ (.A(_06534_),
    .B(_08439_),
    .Y(_08440_));
 sky130_fd_sc_hd__a21oi_1 _13764_ (.A1(net1062),
    .A2(_08440_),
    .B1(net1177),
    .Y(_08441_));
 sky130_fd_sc_hd__a21oi_1 _13765_ (.A1(_05515_),
    .A2(net1201),
    .B1(net1274),
    .Y(_08442_));
 sky130_fd_sc_hd__o221a_1 _13766_ (.A1(_06534_),
    .A2(_06645_),
    .B1(net1203),
    .B2(_05514_),
    .C1(_08442_),
    .X(_08443_));
 sky130_fd_sc_hd__o22a_1 _13767_ (.A1(net1207),
    .A2(_07788_),
    .B1(_07790_),
    .B2(net1215),
    .X(_08444_));
 sky130_fd_sc_hd__a22o_1 _13768_ (.A1(_08438_),
    .A2(_08441_),
    .B1(_08443_),
    .B2(_08444_),
    .X(_08445_));
 sky130_fd_sc_hd__a21o_1 _13769_ (.A1(net1118),
    .A2(_08445_),
    .B1(_08437_),
    .X(_08446_));
 sky130_fd_sc_hd__xnor2_1 _13770_ (.A(net467),
    .B(_08413_),
    .Y(_08447_));
 sky130_fd_sc_hd__a22o_1 _13771_ (.A1(net1221),
    .A2(_08446_),
    .B1(_08447_),
    .B2(net1132),
    .X(_08448_));
 sky130_fd_sc_hd__o21ai_4 _13772_ (.A1(net1251),
    .A2(_06628_),
    .B1(_08448_),
    .Y(_08449_));
 sky130_fd_sc_hd__a211o_4 _13773_ (.A1(\core.pipe0_currentInstruction[25] ),
    .A2(net1220),
    .B1(net983),
    .C1(_08449_),
    .X(_08450_));
 sky130_fd_sc_hd__o211a_1 _13774_ (.A1(\core.pipe1_resultRegister[25] ),
    .A2(net987),
    .B1(_08450_),
    .C1(net1840),
    .X(_00187_));
 sky130_fd_sc_hd__or2_1 _13775_ (.A(_05437_),
    .B(net1116),
    .X(_08451_));
 sky130_fd_sc_hd__a22o_1 _13776_ (.A1(\core.csr.cycleTimer.currentValue[26] ),
    .A2(net725),
    .B1(net721),
    .B2(\core.csr.cycleTimer.currentValue[58] ),
    .X(_08452_));
 sky130_fd_sc_hd__a22o_1 _13777_ (.A1(\core.csr.instretTimer.currentValue[26] ),
    .A2(net701),
    .B1(net697),
    .B2(\core.csr.instretTimer.currentValue[58] ),
    .X(_08453_));
 sky130_fd_sc_hd__nor2_1 _13778_ (.A(\core.csr.cycleTimer.currentValue[26] ),
    .B(net706),
    .Y(_08454_));
 sky130_fd_sc_hd__a221o_1 _13779_ (.A1(\core.csr.cycleTimer.currentValue[58] ),
    .A2(net714),
    .B1(_08453_),
    .B2(net975),
    .C1(net710),
    .X(_08455_));
 sky130_fd_sc_hd__or2_1 _13780_ (.A(\core.csr.traps.mip.csrReadData[26] ),
    .B(net655),
    .X(_08456_));
 sky130_fd_sc_hd__o211a_1 _13781_ (.A1(\core.csr.traps.mtval.csrReadData[26] ),
    .A2(net662),
    .B1(net659),
    .C1(_08456_),
    .X(_08457_));
 sky130_fd_sc_hd__a21o_1 _13782_ (.A1(\core.csr.traps.mcause.csrReadData[26] ),
    .A2(net664),
    .B1(net688),
    .X(_08458_));
 sky130_fd_sc_hd__o221a_1 _13783_ (.A1(\core.csr.trapReturnVector[26] ),
    .A2(net685),
    .B1(_08457_),
    .B2(_08458_),
    .C1(net691),
    .X(_08459_));
 sky130_fd_sc_hd__a221o_1 _13784_ (.A1(\core.csr.traps.mscratch.currentValue[26] ),
    .A2(net694),
    .B1(net676),
    .B2(\core.csr.traps.mtvec.csrReadData[26] ),
    .C1(net682),
    .X(_08460_));
 sky130_fd_sc_hd__o221a_4 _13785_ (.A1(\core.csr.traps.mie.currentValue[26] ),
    .A2(net679),
    .B1(_08459_),
    .B2(_08460_),
    .C1(net607),
    .X(_08461_));
 sky130_fd_sc_hd__a211oi_2 _13786_ (.A1(\core.csr.mconfigptr.currentValue[26] ),
    .A2(net717),
    .B1(_08455_),
    .C1(_08461_),
    .Y(_08462_));
 sky130_fd_sc_hd__o2bb2a_4 _13787_ (.A1_N(net975),
    .A2_N(_08452_),
    .B1(_08454_),
    .B2(_08462_),
    .X(_08463_));
 sky130_fd_sc_hd__inv_2 _13788_ (.A(_08463_),
    .Y(_08464_));
 sky130_fd_sc_hd__o21ai_1 _13789_ (.A1(net1113),
    .A2(_08463_),
    .B1(_08451_),
    .Y(_08465_));
 sky130_fd_sc_hd__a21o_1 _13790_ (.A1(net1110),
    .A2(_08451_),
    .B1(net1104),
    .X(_08466_));
 sky130_fd_sc_hd__and3_1 _13791_ (.A(net1124),
    .B(_08465_),
    .C(_08466_),
    .X(_08467_));
 sky130_fd_sc_hd__a211o_1 _13792_ (.A1(net1153),
    .A2(_06627_),
    .B1(_08013_),
    .C1(_08467_),
    .X(_08468_));
 sky130_fd_sc_hd__a31o_4 _13793_ (.A1(_05592_),
    .A2(_06534_),
    .A3(_07348_),
    .B1(_07353_),
    .X(_08469_));
 sky130_fd_sc_hd__xnor2_4 _13794_ (.A(_05443_),
    .B(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__a21o_1 _13795_ (.A1(net1062),
    .A2(_08470_),
    .B1(net1177),
    .X(_08471_));
 sky130_fd_sc_hd__a21oi_1 _13796_ (.A1(_06627_),
    .A2(net1060),
    .B1(_08471_),
    .Y(_08472_));
 sky130_fd_sc_hd__mux2_1 _13797_ (.A0(net1199),
    .A1(_07458_),
    .S(_05440_),
    .X(_08473_));
 sky130_fd_sc_hd__a21o_1 _13798_ (.A1(net1203),
    .A2(_08473_),
    .B1(_05441_),
    .X(_08474_));
 sky130_fd_sc_hd__o221a_1 _13799_ (.A1(net1208),
    .A2(_07740_),
    .B1(_07745_),
    .B2(net1216),
    .C1(_08474_),
    .X(_08475_));
 sky130_fd_sc_hd__a21oi_1 _13800_ (.A1(net1233),
    .A2(_08475_),
    .B1(_08472_),
    .Y(_08476_));
 sky130_fd_sc_hd__o21ai_1 _13801_ (.A1(_07146_),
    .A2(_08476_),
    .B1(_08468_),
    .Y(_08477_));
 sky130_fd_sc_hd__and3_1 _13802_ (.A(net468),
    .B(net467),
    .C(_08413_),
    .X(_08478_));
 sky130_fd_sc_hd__a21oi_1 _13803_ (.A1(net467),
    .A2(_08413_),
    .B1(net468),
    .Y(_08479_));
 sky130_fd_sc_hd__or2_2 _13804_ (.A(_08478_),
    .B(_08479_),
    .X(_08480_));
 sky130_fd_sc_hd__a22o_1 _13805_ (.A1(net1221),
    .A2(_08477_),
    .B1(_08480_),
    .B2(net1132),
    .X(_08481_));
 sky130_fd_sc_hd__nand2_2 _13806_ (.A(net1254),
    .B(_08481_),
    .Y(_08482_));
 sky130_fd_sc_hd__or2_1 _13807_ (.A(_03879_),
    .B(_06627_),
    .X(_08483_));
 sky130_fd_sc_hd__a221o_4 _13808_ (.A1(\core.pipe0_currentInstruction[26] ),
    .A2(_07141_),
    .B1(_08482_),
    .B2(_08483_),
    .C1(net985),
    .X(_08484_));
 sky130_fd_sc_hd__o211a_1 _13809_ (.A1(\core.pipe1_resultRegister[26] ),
    .A2(net987),
    .B1(_08484_),
    .C1(net1841),
    .X(_00188_));
 sky130_fd_sc_hd__or2_1 _13810_ (.A(_06626_),
    .B(net1063),
    .X(_08485_));
 sky130_fd_sc_hd__a21o_2 _13811_ (.A1(_05442_),
    .A2(_08469_),
    .B1(_07350_),
    .X(_08486_));
 sky130_fd_sc_hd__xnor2_4 _13812_ (.A(_06538_),
    .B(_08486_),
    .Y(_08487_));
 sky130_fd_sc_hd__a21oi_1 _13813_ (.A1(net1063),
    .A2(_08487_),
    .B1(net1177),
    .Y(_08488_));
 sky130_fd_sc_hd__a221o_1 _13814_ (.A1(_05368_),
    .A2(net1205),
    .B1(net1201),
    .B2(_05369_),
    .C1(net1274),
    .X(_08489_));
 sky130_fd_sc_hd__a21oi_1 _13815_ (.A1(_06538_),
    .A2(_06644_),
    .B1(_08489_),
    .Y(_08490_));
 sky130_fd_sc_hd__o22a_1 _13816_ (.A1(net1210),
    .A2(_07696_),
    .B1(_07700_),
    .B2(net1216),
    .X(_08491_));
 sky130_fd_sc_hd__a22o_1 _13817_ (.A1(_08485_),
    .A2(_08488_),
    .B1(_08490_),
    .B2(_08491_),
    .X(_08492_));
 sky130_fd_sc_hd__or2_1 _13818_ (.A(_05364_),
    .B(net1116),
    .X(_08493_));
 sky130_fd_sc_hd__a22o_1 _13819_ (.A1(\core.csr.cycleTimer.currentValue[27] ),
    .A2(net725),
    .B1(net721),
    .B2(\core.csr.cycleTimer.currentValue[59] ),
    .X(_08494_));
 sky130_fd_sc_hd__a22o_1 _13820_ (.A1(\core.csr.instretTimer.currentValue[27] ),
    .A2(net701),
    .B1(net697),
    .B2(\core.csr.instretTimer.currentValue[59] ),
    .X(_08495_));
 sky130_fd_sc_hd__nor2_1 _13821_ (.A(\core.csr.cycleTimer.currentValue[27] ),
    .B(net706),
    .Y(_08496_));
 sky130_fd_sc_hd__a22o_1 _13822_ (.A1(\core.csr.cycleTimer.currentValue[59] ),
    .A2(net714),
    .B1(_08495_),
    .B2(net976),
    .X(_08497_));
 sky130_fd_sc_hd__or2_1 _13823_ (.A(\core.csr.traps.mip.csrReadData[27] ),
    .B(net654),
    .X(_08498_));
 sky130_fd_sc_hd__o211a_1 _13824_ (.A1(\core.csr.traps.mtval.csrReadData[27] ),
    .A2(net661),
    .B1(net658),
    .C1(_08498_),
    .X(_08499_));
 sky130_fd_sc_hd__a21o_1 _13825_ (.A1(\core.csr.traps.mcause.csrReadData[27] ),
    .A2(net664),
    .B1(net688),
    .X(_08500_));
 sky130_fd_sc_hd__o221a_2 _13826_ (.A1(\core.csr.trapReturnVector[27] ),
    .A2(net685),
    .B1(_08499_),
    .B2(_08500_),
    .C1(net691),
    .X(_08501_));
 sky130_fd_sc_hd__a221o_1 _13827_ (.A1(\core.csr.traps.mscratch.currentValue[27] ),
    .A2(net694),
    .B1(net676),
    .B2(\core.csr.traps.mtvec.csrReadData[27] ),
    .C1(net682),
    .X(_08502_));
 sky130_fd_sc_hd__o221a_4 _13828_ (.A1(\core.csr.traps.mie.currentValue[27] ),
    .A2(net679),
    .B1(_08501_),
    .B2(_08502_),
    .C1(net607),
    .X(_08503_));
 sky130_fd_sc_hd__a2111oi_2 _13829_ (.A1(\core.csr.mconfigptr.currentValue[27] ),
    .A2(net719),
    .B1(net710),
    .C1(_08497_),
    .D1(_08503_),
    .Y(_08504_));
 sky130_fd_sc_hd__o2bb2a_4 _13830_ (.A1_N(net975),
    .A2_N(_08494_),
    .B1(_08496_),
    .B2(_08504_),
    .X(_08505_));
 sky130_fd_sc_hd__inv_2 _13831_ (.A(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__o21a_1 _13832_ (.A1(net1113),
    .A2(_08505_),
    .B1(_08493_),
    .X(_08507_));
 sky130_fd_sc_hd__a21oi_1 _13833_ (.A1(net1110),
    .A2(_08493_),
    .B1(net1104),
    .Y(_08508_));
 sky130_fd_sc_hd__o32a_1 _13834_ (.A1(net1120),
    .A2(_08507_),
    .A3(_08508_),
    .B1(_06626_),
    .B2(net1150),
    .X(_08509_));
 sky130_fd_sc_hd__a22o_1 _13835_ (.A1(net1118),
    .A2(_08492_),
    .B1(_08509_),
    .B2(net1059),
    .X(_08510_));
 sky130_fd_sc_hd__and2_2 _13836_ (.A(net469),
    .B(_08478_),
    .X(_08511_));
 sky130_fd_sc_hd__nor2_1 _13837_ (.A(net469),
    .B(_08478_),
    .Y(_08512_));
 sky130_fd_sc_hd__or2_1 _13838_ (.A(_08511_),
    .B(_08512_),
    .X(_08513_));
 sky130_fd_sc_hd__a22o_1 _13839_ (.A1(net1223),
    .A2(_08510_),
    .B1(_08513_),
    .B2(net1132),
    .X(_08514_));
 sky130_fd_sc_hd__o21ai_4 _13840_ (.A1(net1256),
    .A2(_06626_),
    .B1(_08514_),
    .Y(_08515_));
 sky130_fd_sc_hd__a211o_4 _13841_ (.A1(\core.pipe0_currentInstruction[27] ),
    .A2(net1220),
    .B1(net983),
    .C1(_08515_),
    .X(_08516_));
 sky130_fd_sc_hd__o211a_1 _13842_ (.A1(\core.pipe1_resultRegister[27] ),
    .A2(net987),
    .B1(_08516_),
    .C1(net1842),
    .X(_00189_));
 sky130_fd_sc_hd__nand2_1 _13843_ (.A(_05292_),
    .B(net1115),
    .Y(_08517_));
 sky130_fd_sc_hd__a22o_1 _13844_ (.A1(\core.csr.cycleTimer.currentValue[28] ),
    .A2(net725),
    .B1(net721),
    .B2(\core.csr.cycleTimer.currentValue[60] ),
    .X(_08518_));
 sky130_fd_sc_hd__a22o_1 _13845_ (.A1(\core.csr.instretTimer.currentValue[28] ),
    .A2(net701),
    .B1(net697),
    .B2(\core.csr.instretTimer.currentValue[60] ),
    .X(_08519_));
 sky130_fd_sc_hd__nor2_1 _13846_ (.A(\core.csr.cycleTimer.currentValue[28] ),
    .B(net705),
    .Y(_08520_));
 sky130_fd_sc_hd__a22o_1 _13847_ (.A1(\core.csr.cycleTimer.currentValue[60] ),
    .A2(net714),
    .B1(_08519_),
    .B2(net975),
    .X(_08521_));
 sky130_fd_sc_hd__or2_1 _13848_ (.A(\core.csr.traps.mip.csrReadData[28] ),
    .B(net654),
    .X(_08522_));
 sky130_fd_sc_hd__o211a_1 _13849_ (.A1(\core.csr.traps.mtval.csrReadData[28] ),
    .A2(net661),
    .B1(net658),
    .C1(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__a21o_1 _13850_ (.A1(\core.csr.traps.mcause.csrReadData[28] ),
    .A2(net664),
    .B1(net688),
    .X(_08524_));
 sky130_fd_sc_hd__o221a_1 _13851_ (.A1(\core.csr.trapReturnVector[28] ),
    .A2(net685),
    .B1(_08523_),
    .B2(_08524_),
    .C1(net691),
    .X(_08525_));
 sky130_fd_sc_hd__a221o_1 _13852_ (.A1(\core.csr.traps.mscratch.currentValue[28] ),
    .A2(net694),
    .B1(net676),
    .B2(\core.csr.traps.mtvec.csrReadData[28] ),
    .C1(net682),
    .X(_08526_));
 sky130_fd_sc_hd__o221a_4 _13853_ (.A1(\core.csr.traps.mie.currentValue[28] ),
    .A2(net679),
    .B1(_08525_),
    .B2(_08526_),
    .C1(net607),
    .X(_08527_));
 sky130_fd_sc_hd__a2111oi_2 _13854_ (.A1(\core.csr.mconfigptr.currentValue[28] ),
    .A2(net719),
    .B1(net710),
    .C1(_08521_),
    .D1(_08527_),
    .Y(_08528_));
 sky130_fd_sc_hd__o2bb2a_4 _13855_ (.A1_N(net975),
    .A2_N(_08518_),
    .B1(_08520_),
    .B2(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__inv_2 _13856_ (.A(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__o21a_1 _13857_ (.A1(net1113),
    .A2(_08529_),
    .B1(_08517_),
    .X(_08531_));
 sky130_fd_sc_hd__a21oi_1 _13858_ (.A1(net1110),
    .A2(_08517_),
    .B1(net1104),
    .Y(_08532_));
 sky130_fd_sc_hd__or2_1 _13859_ (.A(_06625_),
    .B(net1063),
    .X(_08533_));
 sky130_fd_sc_hd__xor2_2 _13860_ (.A(_06624_),
    .B(_07357_),
    .X(_08534_));
 sky130_fd_sc_hd__nand2_1 _13861_ (.A(net1063),
    .B(_08534_),
    .Y(_08535_));
 sky130_fd_sc_hd__a221oi_1 _13862_ (.A1(_05294_),
    .A2(net1205),
    .B1(net1201),
    .B2(_05295_),
    .C1(net1274),
    .Y(_08536_));
 sky130_fd_sc_hd__o22a_1 _13863_ (.A1(net1210),
    .A2(_07646_),
    .B1(_07652_),
    .B2(net1216),
    .X(_08537_));
 sky130_fd_sc_hd__o211a_1 _13864_ (.A1(_06624_),
    .A2(_06645_),
    .B1(_08536_),
    .C1(_08537_),
    .X(_08538_));
 sky130_fd_sc_hd__a31o_1 _13865_ (.A1(_07950_),
    .A2(_08533_),
    .A3(_08535_),
    .B1(_08538_),
    .X(_08539_));
 sky130_fd_sc_hd__o32a_1 _13866_ (.A1(net1121),
    .A2(_08531_),
    .A3(_08532_),
    .B1(_06625_),
    .B2(net1150),
    .X(_08540_));
 sky130_fd_sc_hd__a22o_1 _13867_ (.A1(net1118),
    .A2(_08539_),
    .B1(_08540_),
    .B2(net1059),
    .X(_08541_));
 sky130_fd_sc_hd__xnor2_1 _13868_ (.A(net470),
    .B(_08511_),
    .Y(_08542_));
 sky130_fd_sc_hd__a22o_1 _13869_ (.A1(net1221),
    .A2(_08541_),
    .B1(_08542_),
    .B2(net1132),
    .X(_08543_));
 sky130_fd_sc_hd__nand2_1 _13870_ (.A(net1254),
    .B(_08543_),
    .Y(_08544_));
 sky130_fd_sc_hd__nand2_1 _13871_ (.A(net1264),
    .B(_06625_),
    .Y(_08545_));
 sky130_fd_sc_hd__a221o_4 _13872_ (.A1(\core.pipe0_currentInstruction[28] ),
    .A2(net1219),
    .B1(_08544_),
    .B2(_08545_),
    .C1(net982),
    .X(_08546_));
 sky130_fd_sc_hd__o211a_1 _13873_ (.A1(\core.pipe1_resultRegister[28] ),
    .A2(net987),
    .B1(_08546_),
    .C1(net1841),
    .X(_00190_));
 sky130_fd_sc_hd__and2_1 _13874_ (.A(_05217_),
    .B(net1115),
    .X(_08547_));
 sky130_fd_sc_hd__a22o_1 _13875_ (.A1(\core.csr.cycleTimer.currentValue[29] ),
    .A2(net726),
    .B1(net722),
    .B2(\core.csr.cycleTimer.currentValue[61] ),
    .X(_08548_));
 sky130_fd_sc_hd__o21ai_1 _13876_ (.A1(\core.csr.cycleTimer.currentValue[29] ),
    .A2(net707),
    .B1(_07250_),
    .Y(_08549_));
 sky130_fd_sc_hd__a22o_1 _13877_ (.A1(\core.csr.instretTimer.currentValue[29] ),
    .A2(net701),
    .B1(net697),
    .B2(\core.csr.instretTimer.currentValue[61] ),
    .X(_08550_));
 sky130_fd_sc_hd__a22o_1 _13878_ (.A1(\core.csr.cycleTimer.currentValue[61] ),
    .A2(net715),
    .B1(_08550_),
    .B2(net976),
    .X(_08551_));
 sky130_fd_sc_hd__or2_1 _13879_ (.A(\core.csr.traps.mip.csrReadData[29] ),
    .B(net654),
    .X(_08552_));
 sky130_fd_sc_hd__o211a_1 _13880_ (.A1(\core.csr.traps.mtval.csrReadData[29] ),
    .A2(net661),
    .B1(net658),
    .C1(_08552_),
    .X(_08553_));
 sky130_fd_sc_hd__a21o_1 _13881_ (.A1(\core.csr.traps.mcause.csrReadData[29] ),
    .A2(net664),
    .B1(net688),
    .X(_08554_));
 sky130_fd_sc_hd__o221a_1 _13882_ (.A1(\core.csr.trapReturnVector[29] ),
    .A2(net685),
    .B1(_08553_),
    .B2(_08554_),
    .C1(net691),
    .X(_08555_));
 sky130_fd_sc_hd__a221o_1 _13883_ (.A1(\core.csr.traps.mscratch.currentValue[29] ),
    .A2(net694),
    .B1(net676),
    .B2(\core.csr.traps.mtvec.csrReadData[29] ),
    .C1(net682),
    .X(_08556_));
 sky130_fd_sc_hd__o221a_4 _13884_ (.A1(\core.csr.traps.mie.currentValue[29] ),
    .A2(net679),
    .B1(_08555_),
    .B2(_08556_),
    .C1(net607),
    .X(_08557_));
 sky130_fd_sc_hd__a2111oi_2 _13885_ (.A1(\core.csr.mconfigptr.currentValue[29] ),
    .A2(net719),
    .B1(net711),
    .C1(_08551_),
    .D1(_08557_),
    .Y(_08558_));
 sky130_fd_sc_hd__a2bb2o_4 _13886_ (.A1_N(_08549_),
    .A2_N(_08558_),
    .B1(net976),
    .B2(_08548_),
    .X(_08559_));
 sky130_fd_sc_hd__a21oi_1 _13887_ (.A1(net1111),
    .A2(_08559_),
    .B1(_08547_),
    .Y(_08560_));
 sky130_fd_sc_hd__o21a_1 _13888_ (.A1(net1108),
    .A2(_08547_),
    .B1(net1106),
    .X(_08561_));
 sky130_fd_sc_hd__o32a_1 _13889_ (.A1(net1121),
    .A2(_08560_),
    .A3(_08561_),
    .B1(_06623_),
    .B2(net1150),
    .X(_08562_));
 sky130_fd_sc_hd__a21boi_4 _13890_ (.A1(_06624_),
    .A2(_07357_),
    .B1_N(_07360_),
    .Y(_08563_));
 sky130_fd_sc_hd__xnor2_4 _13891_ (.A(_06622_),
    .B(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__a21oi_1 _13892_ (.A1(net1064),
    .A2(_08564_),
    .B1(net1177),
    .Y(_08565_));
 sky130_fd_sc_hd__o21a_1 _13893_ (.A1(_06623_),
    .A2(net1064),
    .B1(_08565_),
    .X(_08566_));
 sky130_fd_sc_hd__a21oi_1 _13894_ (.A1(_05221_),
    .A2(net1201),
    .B1(net1274),
    .Y(_08567_));
 sky130_fd_sc_hd__o221a_1 _13895_ (.A1(_06622_),
    .A2(_06645_),
    .B1(net1203),
    .B2(_05219_),
    .C1(_08567_),
    .X(_08568_));
 sky130_fd_sc_hd__o22a_1 _13896_ (.A1(net1208),
    .A2(_07591_),
    .B1(_07597_),
    .B2(net1215),
    .X(_08569_));
 sky130_fd_sc_hd__a21oi_1 _13897_ (.A1(_08568_),
    .A2(_08569_),
    .B1(_08566_),
    .Y(_08570_));
 sky130_fd_sc_hd__a2bb2o_1 _13898_ (.A1_N(_07146_),
    .A2_N(_08570_),
    .B1(_08562_),
    .B2(_08012_),
    .X(_08571_));
 sky130_fd_sc_hd__nand2_1 _13899_ (.A(net1223),
    .B(_08571_),
    .Y(_08572_));
 sky130_fd_sc_hd__and3_2 _13900_ (.A(net471),
    .B(net470),
    .C(_08511_),
    .X(_08573_));
 sky130_fd_sc_hd__a21oi_1 _13901_ (.A1(net470),
    .A2(_08511_),
    .B1(net471),
    .Y(_08574_));
 sky130_fd_sc_hd__nor2_2 _13902_ (.A(_08573_),
    .B(_08574_),
    .Y(_08575_));
 sky130_fd_sc_hd__or2_1 _13903_ (.A(net1136),
    .B(_08575_),
    .X(_08576_));
 sky130_fd_sc_hd__nor2_1 _13904_ (.A(net1254),
    .B(_06623_),
    .Y(_08577_));
 sky130_fd_sc_hd__a221o_1 _13905_ (.A1(\core.pipe0_currentInstruction[29] ),
    .A2(net1219),
    .B1(_08572_),
    .B2(_08576_),
    .C1(net982),
    .X(_08578_));
 sky130_fd_sc_hd__o221a_1 _13906_ (.A1(\core.pipe1_resultRegister[29] ),
    .A2(net988),
    .B1(_08577_),
    .B2(_08578_),
    .C1(net1824),
    .X(_00191_));
 sky130_fd_sc_hd__a31o_4 _13907_ (.A1(_06622_),
    .A2(_06624_),
    .A3(_07357_),
    .B1(_07361_),
    .X(_08579_));
 sky130_fd_sc_hd__xnor2_4 _13908_ (.A(_05149_),
    .B(_08579_),
    .Y(_08580_));
 sky130_fd_sc_hd__a21oi_1 _13909_ (.A1(net1064),
    .A2(_08580_),
    .B1(net1178),
    .Y(_08581_));
 sky130_fd_sc_hd__o21a_1 _13910_ (.A1(_06543_),
    .A2(net1064),
    .B1(_08581_),
    .X(_08582_));
 sky130_fd_sc_hd__nand2_1 _13911_ (.A(net1213),
    .B(_07530_),
    .Y(_08583_));
 sky130_fd_sc_hd__a21oi_1 _13912_ (.A1(_05146_),
    .A2(net1201),
    .B1(net1205),
    .Y(_08584_));
 sky130_fd_sc_hd__or2_1 _13913_ (.A(_05147_),
    .B(_08584_),
    .X(_08585_));
 sky130_fd_sc_hd__o221a_1 _13914_ (.A1(net1218),
    .A2(_07535_),
    .B1(net1198),
    .B2(_05148_),
    .C1(_08585_),
    .X(_08586_));
 sky130_fd_sc_hd__a31o_1 _13915_ (.A1(net1233),
    .A2(_08583_),
    .A3(_08586_),
    .B1(_08582_),
    .X(_08587_));
 sky130_fd_sc_hd__or2_1 _13916_ (.A(_04068_),
    .B(_06543_),
    .X(_08588_));
 sky130_fd_sc_hd__nor2_1 _13917_ (.A(_05143_),
    .B(net1117),
    .Y(_08589_));
 sky130_fd_sc_hd__a22o_1 _13918_ (.A1(\core.csr.cycleTimer.currentValue[30] ),
    .A2(net726),
    .B1(net722),
    .B2(\core.csr.cycleTimer.currentValue[62] ),
    .X(_08590_));
 sky130_fd_sc_hd__a22o_1 _13919_ (.A1(\core.csr.instretTimer.currentValue[30] ),
    .A2(net701),
    .B1(net697),
    .B2(\core.csr.instretTimer.currentValue[62] ),
    .X(_08591_));
 sky130_fd_sc_hd__a221o_1 _13920_ (.A1(\core.csr.cycleTimer.currentValue[62] ),
    .A2(net715),
    .B1(_08591_),
    .B2(net976),
    .C1(net711),
    .X(_08592_));
 sky130_fd_sc_hd__mux2_1 _13921_ (.A0(\core.csr.traps.mip.csrReadData[30] ),
    .A1(\core.csr.traps.mtval.csrReadData[30] ),
    .S(net655),
    .X(_08593_));
 sky130_fd_sc_hd__a221o_1 _13922_ (.A1(\core.csr.traps.mcause.csrReadData[30] ),
    .A2(_07281_),
    .B1(_07472_),
    .B2(_08593_),
    .C1(_07283_),
    .X(_08594_));
 sky130_fd_sc_hd__o21a_2 _13923_ (.A1(\core.csr.trapReturnVector[30] ),
    .A2(_07284_),
    .B1(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__a221o_1 _13924_ (.A1(\core.csr.traps.mtvec.csrReadData[30] ),
    .A2(_07231_),
    .B1(_07280_),
    .B2(\core.csr.traps.mscratch.currentValue[30] ),
    .C1(_08595_),
    .X(_08596_));
 sky130_fd_sc_hd__mux2_1 _13925_ (.A0(\core.csr.traps.mie.currentValue[30] ),
    .A1(_08596_),
    .S(_07219_),
    .X(_08597_));
 sky130_fd_sc_hd__o32a_2 _13926_ (.A1(\core.csr.mconfigptr.currentValue[30] ),
    .A2(_07230_),
    .A3(_07274_),
    .B1(_07875_),
    .B2(_08597_),
    .X(_08598_));
 sky130_fd_sc_hd__o22a_1 _13927_ (.A1(\core.csr.cycleTimer.currentValue[30] ),
    .A2(net707),
    .B1(_08592_),
    .B2(_08598_),
    .X(_08599_));
 sky130_fd_sc_hd__a21o_4 _13928_ (.A1(net975),
    .A2(_08590_),
    .B1(_08599_),
    .X(_08600_));
 sky130_fd_sc_hd__a21oi_1 _13929_ (.A1(net1111),
    .A2(_08600_),
    .B1(_08589_),
    .Y(_08601_));
 sky130_fd_sc_hd__o21a_1 _13930_ (.A1(net1108),
    .A2(_08589_),
    .B1(net1106),
    .X(_08602_));
 sky130_fd_sc_hd__or3_1 _13931_ (.A(net1120),
    .B(_08601_),
    .C(_08602_),
    .X(_08603_));
 sky130_fd_sc_hd__a32o_1 _13932_ (.A1(_08012_),
    .A2(_08588_),
    .A3(_08603_),
    .B1(_08587_),
    .B2(net1119),
    .X(_08604_));
 sky130_fd_sc_hd__nand2_2 _13933_ (.A(net473),
    .B(_08573_),
    .Y(_08605_));
 sky130_fd_sc_hd__or2_1 _13934_ (.A(net473),
    .B(_08573_),
    .X(_08606_));
 sky130_fd_sc_hd__nand2_2 _13935_ (.A(_08605_),
    .B(_08606_),
    .Y(_08607_));
 sky130_fd_sc_hd__a22o_1 _13936_ (.A1(net1225),
    .A2(_08604_),
    .B1(_08607_),
    .B2(net1134),
    .X(_08608_));
 sky130_fd_sc_hd__nand2_1 _13937_ (.A(net1259),
    .B(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__nand2_1 _13938_ (.A(net1264),
    .B(_06543_),
    .Y(_08610_));
 sky130_fd_sc_hd__a221o_4 _13939_ (.A1(net1752),
    .A2(net1220),
    .B1(_08609_),
    .B2(_08610_),
    .C1(net983),
    .X(_08611_));
 sky130_fd_sc_hd__o211a_1 _13940_ (.A1(\core.pipe1_resultRegister[30] ),
    .A2(net987),
    .B1(_08611_),
    .C1(net1841),
    .X(_00192_));
 sky130_fd_sc_hd__or2_1 _13941_ (.A(_06612_),
    .B(net1117),
    .X(_08612_));
 sky130_fd_sc_hd__a22o_1 _13942_ (.A1(\core.csr.cycleTimer.currentValue[31] ),
    .A2(net726),
    .B1(net722),
    .B2(\core.csr.cycleTimer.currentValue[63] ),
    .X(_08613_));
 sky130_fd_sc_hd__a22o_1 _13943_ (.A1(\core.csr.instretTimer.currentValue[31] ),
    .A2(net701),
    .B1(net697),
    .B2(\core.csr.instretTimer.currentValue[63] ),
    .X(_08614_));
 sky130_fd_sc_hd__nor2_1 _13944_ (.A(\core.csr.cycleTimer.currentValue[31] ),
    .B(net707),
    .Y(_08615_));
 sky130_fd_sc_hd__a22o_1 _13945_ (.A1(\core.csr.cycleTimer.currentValue[63] ),
    .A2(net715),
    .B1(_08614_),
    .B2(net978),
    .X(_08616_));
 sky130_fd_sc_hd__or2_1 _13946_ (.A(\core.csr.traps.mip.csrReadData[31] ),
    .B(net654),
    .X(_08617_));
 sky130_fd_sc_hd__o211a_1 _13947_ (.A1(\core.csr.traps.mtval.csrReadData[31] ),
    .A2(net661),
    .B1(net658),
    .C1(_08617_),
    .X(_08618_));
 sky130_fd_sc_hd__a21o_1 _13948_ (.A1(\core.csr.traps.mcause.csrReadData[31] ),
    .A2(net664),
    .B1(net688),
    .X(_08619_));
 sky130_fd_sc_hd__o221a_1 _13949_ (.A1(\core.csr.trapReturnVector[31] ),
    .A2(net685),
    .B1(_08618_),
    .B2(_08619_),
    .C1(net691),
    .X(_08620_));
 sky130_fd_sc_hd__a221o_1 _13950_ (.A1(\core.csr.traps.mscratch.currentValue[31] ),
    .A2(net695),
    .B1(net677),
    .B2(\core.csr.traps.mtvec.csrReadData[31] ),
    .C1(net683),
    .X(_08621_));
 sky130_fd_sc_hd__o221a_4 _13951_ (.A1(\core.csr.traps.mie.currentValue[31] ),
    .A2(net680),
    .B1(_08620_),
    .B2(_08621_),
    .C1(net608),
    .X(_08622_));
 sky130_fd_sc_hd__a2111oi_2 _13952_ (.A1(\core.csr.mconfigptr.currentValue[31] ),
    .A2(net719),
    .B1(net711),
    .C1(_08616_),
    .D1(_08622_),
    .Y(_08623_));
 sky130_fd_sc_hd__o2bb2a_4 _13953_ (.A1_N(net978),
    .A2_N(_08613_),
    .B1(_08615_),
    .B2(_08623_),
    .X(_08624_));
 sky130_fd_sc_hd__inv_2 _13954_ (.A(_08624_),
    .Y(_08625_));
 sky130_fd_sc_hd__o21a_1 _13955_ (.A1(net1113),
    .A2(_08624_),
    .B1(_08612_),
    .X(_08626_));
 sky130_fd_sc_hd__a21oi_1 _13956_ (.A1(net1110),
    .A2(_08612_),
    .B1(net1104),
    .Y(_08627_));
 sky130_fd_sc_hd__o32a_1 _13957_ (.A1(net1120),
    .A2(_08626_),
    .A3(_08627_),
    .B1(_06619_),
    .B2(net1150),
    .X(_08628_));
 sky130_fd_sc_hd__or2_1 _13958_ (.A(_06619_),
    .B(net1064),
    .X(_08629_));
 sky130_fd_sc_hd__a211o_1 _13959_ (.A1(_05148_),
    .A2(_08579_),
    .B1(_07362_),
    .C1(_06617_),
    .X(_08630_));
 sky130_fd_sc_hd__o21ai_4 _13960_ (.A1(_06615_),
    .A2(_07364_),
    .B1(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__or2_1 _13961_ (.A(net1060),
    .B(_08631_),
    .X(_08632_));
 sky130_fd_sc_hd__nor2_1 _13962_ (.A(_06613_),
    .B(net1203),
    .Y(_08633_));
 sky130_fd_sc_hd__o21ai_1 _13963_ (.A1(_06613_),
    .A2(_07458_),
    .B1(net1203),
    .Y(_08634_));
 sky130_fd_sc_hd__o21ai_1 _13964_ (.A1(_06580_),
    .A2(_08633_),
    .B1(_08634_),
    .Y(_08635_));
 sky130_fd_sc_hd__o221a_1 _13965_ (.A1(_06617_),
    .A2(_06645_),
    .B1(net1212),
    .B2(_07441_),
    .C1(_08635_),
    .X(_08636_));
 sky130_fd_sc_hd__o211a_1 _13966_ (.A1(net1218),
    .A2(_07454_),
    .B1(_08636_),
    .C1(net1233),
    .X(_08637_));
 sky130_fd_sc_hd__a31o_1 _13967_ (.A1(_07950_),
    .A2(_08629_),
    .A3(_08632_),
    .B1(_08637_),
    .X(_08638_));
 sky130_fd_sc_hd__a22o_1 _13968_ (.A1(net1059),
    .A2(_08628_),
    .B1(_08638_),
    .B2(net1119),
    .X(_08639_));
 sky130_fd_sc_hd__xnor2_2 _13969_ (.A(_03823_),
    .B(_08605_),
    .Y(_08640_));
 sky130_fd_sc_hd__a22o_1 _13970_ (.A1(net1222),
    .A2(_08639_),
    .B1(_08640_),
    .B2(net1135),
    .X(_08641_));
 sky130_fd_sc_hd__a21o_1 _13971_ (.A1(net1751),
    .A2(net1219),
    .B1(net982),
    .X(_08642_));
 sky130_fd_sc_hd__o21ai_1 _13972_ (.A1(net1255),
    .A2(_06619_),
    .B1(_08641_),
    .Y(_08643_));
 sky130_fd_sc_hd__o221a_1 _13973_ (.A1(\core.pipe1_resultRegister[31] ),
    .A2(net988),
    .B1(_08642_),
    .B2(_08643_),
    .C1(net1805),
    .X(_00193_));
 sky130_fd_sc_hd__or2_1 _13974_ (.A(\core.pipe1_csrData[0] ),
    .B(net1072),
    .X(_08644_));
 sky130_fd_sc_hd__o211a_1 _13975_ (.A1(net1068),
    .A2(_07252_),
    .B1(_08644_),
    .C1(net1838),
    .X(_00194_));
 sky130_fd_sc_hd__nand2_1 _13976_ (.A(net1074),
    .B(_07484_),
    .Y(_08645_));
 sky130_fd_sc_hd__o211a_1 _13977_ (.A1(\core.pipe1_csrData[1] ),
    .A2(net1074),
    .B1(_08645_),
    .C1(net1858),
    .X(_00195_));
 sky130_fd_sc_hd__nand2_1 _13978_ (.A(net1071),
    .B(_07564_),
    .Y(_08646_));
 sky130_fd_sc_hd__o211a_1 _13979_ (.A1(\core.pipe1_csrData[2] ),
    .A2(net1071),
    .B1(_08646_),
    .C1(net1836),
    .X(_00196_));
 sky130_fd_sc_hd__nand2_1 _13980_ (.A(net1071),
    .B(_07620_),
    .Y(_08647_));
 sky130_fd_sc_hd__o211a_1 _13981_ (.A1(\core.pipe1_csrData[3] ),
    .A2(net1071),
    .B1(_08647_),
    .C1(net1836),
    .X(_00197_));
 sky130_fd_sc_hd__or2_1 _13982_ (.A(\core.pipe1_csrData[4] ),
    .B(net1069),
    .X(_08648_));
 sky130_fd_sc_hd__o211a_1 _13983_ (.A1(net1068),
    .A2(_07676_),
    .B1(_08648_),
    .C1(net1838),
    .X(_00198_));
 sky130_fd_sc_hd__or2_1 _13984_ (.A(\core.pipe1_csrData[5] ),
    .B(net1071),
    .X(_08649_));
 sky130_fd_sc_hd__o211a_1 _13985_ (.A1(net1068),
    .A2(_07721_),
    .B1(_08649_),
    .C1(net1837),
    .X(_00199_));
 sky130_fd_sc_hd__nand2_1 _13986_ (.A(net1071),
    .B(_07771_),
    .Y(_08650_));
 sky130_fd_sc_hd__o211a_1 _13987_ (.A1(\core.pipe1_csrData[6] ),
    .A2(net1071),
    .B1(_08650_),
    .C1(net1855),
    .X(_00200_));
 sky130_fd_sc_hd__nand2_1 _13988_ (.A(net1069),
    .B(_07812_),
    .Y(_08651_));
 sky130_fd_sc_hd__o211a_1 _13989_ (.A1(\core.pipe1_csrData[7] ),
    .A2(net1069),
    .B1(_08651_),
    .C1(net1838),
    .X(_00201_));
 sky130_fd_sc_hd__nand2_1 _13990_ (.A(net1073),
    .B(_07873_),
    .Y(_08652_));
 sky130_fd_sc_hd__o211a_1 _13991_ (.A1(\core.pipe1_csrData[8] ),
    .A2(net1074),
    .B1(_08652_),
    .C1(net1858),
    .X(_00202_));
 sky130_fd_sc_hd__or2_1 _13992_ (.A(\core.pipe1_csrData[9] ),
    .B(net1072),
    .X(_08653_));
 sky130_fd_sc_hd__o211a_1 _13993_ (.A1(net1068),
    .A2(_07910_),
    .B1(_08653_),
    .C1(net1841),
    .X(_00203_));
 sky130_fd_sc_hd__or2_1 _13994_ (.A(\core.pipe1_csrData[10] ),
    .B(net1073),
    .X(_08654_));
 sky130_fd_sc_hd__o211a_1 _13995_ (.A1(net1068),
    .A2(_07943_),
    .B1(_08654_),
    .C1(net1856),
    .X(_00204_));
 sky130_fd_sc_hd__nand2_1 _13996_ (.A(net1073),
    .B(_07977_),
    .Y(_08655_));
 sky130_fd_sc_hd__o211a_1 _13997_ (.A1(\core.pipe1_csrData[11] ),
    .A2(net1073),
    .B1(_08655_),
    .C1(net1856),
    .X(_00205_));
 sky130_fd_sc_hd__nand2_1 _13998_ (.A(net1073),
    .B(_07997_),
    .Y(_08656_));
 sky130_fd_sc_hd__o211a_1 _13999_ (.A1(\core.pipe1_csrData[12] ),
    .A2(net1073),
    .B1(_08656_),
    .C1(net1841),
    .X(_00206_));
 sky130_fd_sc_hd__nand2_1 _14000_ (.A(net1073),
    .B(_08034_),
    .Y(_08657_));
 sky130_fd_sc_hd__o211a_1 _14001_ (.A1(\core.pipe1_csrData[13] ),
    .A2(net1074),
    .B1(_08657_),
    .C1(net1858),
    .X(_00207_));
 sky130_fd_sc_hd__nand2_1 _14002_ (.A(net1072),
    .B(_08069_),
    .Y(_08658_));
 sky130_fd_sc_hd__o211a_1 _14003_ (.A1(\core.pipe1_csrData[14] ),
    .A2(net1072),
    .B1(_08658_),
    .C1(net1842),
    .X(_00208_));
 sky130_fd_sc_hd__nand2_1 _14004_ (.A(net1071),
    .B(_08122_),
    .Y(_08659_));
 sky130_fd_sc_hd__o211a_1 _14005_ (.A1(\core.pipe1_csrData[15] ),
    .A2(net1070),
    .B1(_08659_),
    .C1(net1838),
    .X(_00209_));
 sky130_fd_sc_hd__nand2_1 _14006_ (.A(net1070),
    .B(_08144_),
    .Y(_08660_));
 sky130_fd_sc_hd__o211a_1 _14007_ (.A1(\core.pipe1_csrData[16] ),
    .A2(net1070),
    .B1(_08660_),
    .C1(net1838),
    .X(_00210_));
 sky130_fd_sc_hd__nand2_1 _14008_ (.A(net1070),
    .B(_08189_),
    .Y(_08661_));
 sky130_fd_sc_hd__o211a_1 _14009_ (.A1(\core.pipe1_csrData[17] ),
    .A2(net1070),
    .B1(_08661_),
    .C1(net1838),
    .X(_00211_));
 sky130_fd_sc_hd__or2_1 _14010_ (.A(\core.pipe1_csrData[18] ),
    .B(net1072),
    .X(_08662_));
 sky130_fd_sc_hd__o211a_1 _14011_ (.A1(net1068),
    .A2(_08211_),
    .B1(_08662_),
    .C1(net1841),
    .X(_00212_));
 sky130_fd_sc_hd__nand2_1 _14012_ (.A(net1069),
    .B(_08243_),
    .Y(_08663_));
 sky130_fd_sc_hd__o211a_1 _14013_ (.A1(\core.pipe1_csrData[19] ),
    .A2(net1069),
    .B1(_08663_),
    .C1(net1838),
    .X(_00213_));
 sky130_fd_sc_hd__nand2_1 _14014_ (.A(net1069),
    .B(_08275_),
    .Y(_08664_));
 sky130_fd_sc_hd__o211a_1 _14015_ (.A1(\core.pipe1_csrData[20] ),
    .A2(net1070),
    .B1(_08664_),
    .C1(net1838),
    .X(_00214_));
 sky130_fd_sc_hd__nand2_1 _14016_ (.A(net1070),
    .B(_08316_),
    .Y(_08665_));
 sky130_fd_sc_hd__o211a_1 _14017_ (.A1(\core.pipe1_csrData[21] ),
    .A2(net1069),
    .B1(_08665_),
    .C1(net1838),
    .X(_00215_));
 sky130_fd_sc_hd__or2_1 _14018_ (.A(\core.pipe1_csrData[22] ),
    .B(net1069),
    .X(_08666_));
 sky130_fd_sc_hd__o211a_1 _14019_ (.A1(net1068),
    .A2(_08339_),
    .B1(_08666_),
    .C1(net1837),
    .X(_00216_));
 sky130_fd_sc_hd__or2_1 _14020_ (.A(\core.pipe1_csrData[23] ),
    .B(net1069),
    .X(_08667_));
 sky130_fd_sc_hd__o211a_1 _14021_ (.A1(net1068),
    .A2(_08370_),
    .B1(_08667_),
    .C1(net1837),
    .X(_00217_));
 sky130_fd_sc_hd__or2_1 _14022_ (.A(\core.pipe1_csrData[24] ),
    .B(net1070),
    .X(_08668_));
 sky130_fd_sc_hd__o211a_1 _14023_ (.A1(net1068),
    .A2(_08401_),
    .B1(_08668_),
    .C1(net1840),
    .X(_00218_));
 sky130_fd_sc_hd__nand2_1 _14024_ (.A(net1072),
    .B(_08432_),
    .Y(_08669_));
 sky130_fd_sc_hd__o211a_1 _14025_ (.A1(\core.pipe1_csrData[25] ),
    .A2(net1072),
    .B1(_08669_),
    .C1(net1841),
    .X(_00219_));
 sky130_fd_sc_hd__nand2_1 _14026_ (.A(net1072),
    .B(_08463_),
    .Y(_08670_));
 sky130_fd_sc_hd__o211a_1 _14027_ (.A1(\core.pipe1_csrData[26] ),
    .A2(net1075),
    .B1(_08670_),
    .C1(net1841),
    .X(_00220_));
 sky130_fd_sc_hd__nand2_1 _14028_ (.A(net1072),
    .B(_08505_),
    .Y(_08671_));
 sky130_fd_sc_hd__o211a_1 _14029_ (.A1(\core.pipe1_csrData[27] ),
    .A2(net1072),
    .B1(_08671_),
    .C1(net1841),
    .X(_00221_));
 sky130_fd_sc_hd__nand2_1 _14030_ (.A(net1073),
    .B(_08529_),
    .Y(_08672_));
 sky130_fd_sc_hd__o211a_1 _14031_ (.A1(\core.pipe1_csrData[28] ),
    .A2(net1073),
    .B1(_08672_),
    .C1(net1856),
    .X(_00222_));
 sky130_fd_sc_hd__or2_1 _14032_ (.A(\core.pipe1_csrData[29] ),
    .B(net1073),
    .X(_08673_));
 sky130_fd_sc_hd__o211a_1 _14033_ (.A1(net1068),
    .A2(_08559_),
    .B1(_08673_),
    .C1(net1856),
    .X(_00223_));
 sky130_fd_sc_hd__or2_1 _14034_ (.A(\core.pipe1_csrData[30] ),
    .B(net1074),
    .X(_08674_));
 sky130_fd_sc_hd__o211a_1 _14035_ (.A1(_07163_),
    .A2(_08600_),
    .B1(_08674_),
    .C1(net1856),
    .X(_00224_));
 sky130_fd_sc_hd__nand2_1 _14036_ (.A(net1070),
    .B(_08624_),
    .Y(_08675_));
 sky130_fd_sc_hd__o211a_1 _14037_ (.A1(\core.pipe1_csrData[31] ),
    .A2(net1069),
    .B1(_08675_),
    .C1(net1838),
    .X(_00225_));
 sky130_fd_sc_hd__and3b_4 _14038_ (.A_N(\core.csr.currentInstruction[10] ),
    .B(net1801),
    .C(_03904_),
    .X(_08676_));
 sky130_fd_sc_hd__nor3_4 _14039_ (.A(\core.csr.currentInstruction[8] ),
    .B(_03910_),
    .C(_06849_),
    .Y(_08677_));
 sky130_fd_sc_hd__or3_2 _14040_ (.A(\core.csr.currentInstruction[8] ),
    .B(_03910_),
    .C(_06849_),
    .X(_08678_));
 sky130_fd_sc_hd__nand2_8 _14041_ (.A(_08676_),
    .B(_08677_),
    .Y(_08679_));
 sky130_fd_sc_hd__mux2_1 _14042_ (.A0(net1078),
    .A1(\core.registers[21][0] ),
    .S(net970),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _14043_ (.A0(net1082),
    .A1(\core.registers[21][1] ),
    .S(net972),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _14044_ (.A0(net1085),
    .A1(\core.registers[21][2] ),
    .S(net970),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _14045_ (.A0(net1090),
    .A1(\core.registers[21][3] ),
    .S(net969),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _14046_ (.A0(net1027),
    .A1(\core.registers[21][4] ),
    .S(net972),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _14047_ (.A0(net1032),
    .A1(\core.registers[21][5] ),
    .S(net972),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _14048_ (.A0(net1036),
    .A1(\core.registers[21][6] ),
    .S(net972),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _14049_ (.A0(net1138),
    .A1(\core.registers[21][7] ),
    .S(net972),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _14050_ (.A0(net899),
    .A1(\core.registers[21][8] ),
    .S(net971),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _14051_ (.A0(net902),
    .A1(\core.registers[21][9] ),
    .S(net971),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _14052_ (.A0(net759),
    .A1(\core.registers[21][10] ),
    .S(net971),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _14053_ (.A0(net761),
    .A1(\core.registers[21][11] ),
    .S(net971),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _14054_ (.A0(net729),
    .A1(\core.registers[21][12] ),
    .S(net971),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _14055_ (.A0(net733),
    .A1(\core.registers[21][13] ),
    .S(net972),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _14056_ (.A0(net738),
    .A1(\core.registers[21][14] ),
    .S(net969),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _14057_ (.A0(net741),
    .A1(\core.registers[21][15] ),
    .S(net970),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _14058_ (.A0(net830),
    .A1(\core.registers[21][16] ),
    .S(net970),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _14059_ (.A0(net836),
    .A1(\core.registers[21][17] ),
    .S(net969),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _14060_ (.A0(net838),
    .A1(\core.registers[21][18] ),
    .S(net971),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _14061_ (.A0(net843),
    .A1(\core.registers[21][19] ),
    .S(net969),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _14062_ (.A0(net847),
    .A1(\core.registers[21][20] ),
    .S(net969),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _14063_ (.A0(net852),
    .A1(\core.registers[21][21] ),
    .S(net969),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _14064_ (.A0(net858),
    .A1(\core.registers[21][22] ),
    .S(net970),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _14065_ (.A0(net862),
    .A1(\core.registers[21][23] ),
    .S(net969),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _14066_ (.A0(net994),
    .A1(\core.registers[21][24] ),
    .S(net969),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _14067_ (.A0(net998),
    .A1(\core.registers[21][25] ),
    .S(net969),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _14068_ (.A0(net1002),
    .A1(\core.registers[21][26] ),
    .S(net971),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _14069_ (.A0(net866),
    .A1(\core.registers[21][27] ),
    .S(net971),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _14070_ (.A0(net871),
    .A1(\core.registers[21][28] ),
    .S(net972),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _14071_ (.A0(net874),
    .A1(\core.registers[21][29] ),
    .S(net971),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _14072_ (.A0(net878),
    .A1(\core.registers[21][30] ),
    .S(net971),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _14073_ (.A0(net1023),
    .A1(\core.registers[21][31] ),
    .S(net969),
    .X(_00257_));
 sky130_fd_sc_hd__and3b_4 _14074_ (.A_N(_06849_),
    .B(_03911_),
    .C(_03910_),
    .X(_08680_));
 sky130_fd_sc_hd__nand2_8 _14075_ (.A(_08676_),
    .B(_08680_),
    .Y(_08681_));
 sky130_fd_sc_hd__mux2_1 _14076_ (.A0(net1079),
    .A1(\core.registers[20][0] ),
    .S(net966),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _14077_ (.A0(net1082),
    .A1(\core.registers[20][1] ),
    .S(net968),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _14078_ (.A0(net1085),
    .A1(\core.registers[20][2] ),
    .S(net966),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _14079_ (.A0(net1090),
    .A1(\core.registers[20][3] ),
    .S(net965),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _14080_ (.A0(net1027),
    .A1(\core.registers[20][4] ),
    .S(net968),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _14081_ (.A0(net1032),
    .A1(\core.registers[20][5] ),
    .S(net968),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _14082_ (.A0(net1035),
    .A1(\core.registers[20][6] ),
    .S(net968),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _14083_ (.A0(net1139),
    .A1(\core.registers[20][7] ),
    .S(net968),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _14084_ (.A0(net899),
    .A1(\core.registers[20][8] ),
    .S(net967),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _14085_ (.A0(net903),
    .A1(\core.registers[20][9] ),
    .S(net967),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _14086_ (.A0(net759),
    .A1(\core.registers[20][10] ),
    .S(net967),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _14087_ (.A0(net761),
    .A1(\core.registers[20][11] ),
    .S(net967),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _14088_ (.A0(net729),
    .A1(\core.registers[20][12] ),
    .S(net967),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _14089_ (.A0(net733),
    .A1(\core.registers[20][13] ),
    .S(net968),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _14090_ (.A0(net738),
    .A1(\core.registers[20][14] ),
    .S(net965),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _14091_ (.A0(net740),
    .A1(\core.registers[20][15] ),
    .S(net966),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _14092_ (.A0(net830),
    .A1(\core.registers[20][16] ),
    .S(net966),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _14093_ (.A0(net836),
    .A1(\core.registers[20][17] ),
    .S(net965),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _14094_ (.A0(net838),
    .A1(\core.registers[20][18] ),
    .S(net967),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _14095_ (.A0(net843),
    .A1(\core.registers[20][19] ),
    .S(net965),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _14096_ (.A0(net847),
    .A1(\core.registers[20][20] ),
    .S(net965),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _14097_ (.A0(net852),
    .A1(\core.registers[20][21] ),
    .S(net965),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _14098_ (.A0(net858),
    .A1(\core.registers[20][22] ),
    .S(net966),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _14099_ (.A0(net862),
    .A1(\core.registers[20][23] ),
    .S(net965),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _14100_ (.A0(net994),
    .A1(\core.registers[20][24] ),
    .S(net965),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _14101_ (.A0(net998),
    .A1(\core.registers[20][25] ),
    .S(net965),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _14102_ (.A0(net1002),
    .A1(\core.registers[20][26] ),
    .S(net967),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _14103_ (.A0(net866),
    .A1(\core.registers[20][27] ),
    .S(net967),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _14104_ (.A0(net870),
    .A1(\core.registers[20][28] ),
    .S(net968),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _14105_ (.A0(net874),
    .A1(\core.registers[20][29] ),
    .S(net967),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _14106_ (.A0(net878),
    .A1(\core.registers[20][30] ),
    .S(net967),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _14107_ (.A0(net1023),
    .A1(\core.registers[20][31] ),
    .S(net965),
    .X(_00289_));
 sky130_fd_sc_hd__nand2_8 _14108_ (.A(_03908_),
    .B(_08677_),
    .Y(_08682_));
 sky130_fd_sc_hd__mux2_1 _14109_ (.A0(net1078),
    .A1(\core.registers[1][0] ),
    .S(net962),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _14110_ (.A0(net1081),
    .A1(\core.registers[1][1] ),
    .S(net964),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _14111_ (.A0(net1088),
    .A1(\core.registers[1][2] ),
    .S(net962),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _14112_ (.A0(net1092),
    .A1(\core.registers[1][3] ),
    .S(net961),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _14113_ (.A0(net1028),
    .A1(\core.registers[1][4] ),
    .S(net962),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _14114_ (.A0(net1034),
    .A1(\core.registers[1][5] ),
    .S(net962),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _14115_ (.A0(net1035),
    .A1(\core.registers[1][6] ),
    .S(net962),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _14116_ (.A0(net1139),
    .A1(\core.registers[1][7] ),
    .S(net964),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _14117_ (.A0(net898),
    .A1(\core.registers[1][8] ),
    .S(net963),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _14118_ (.A0(net902),
    .A1(\core.registers[1][9] ),
    .S(net963),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _14119_ (.A0(net760),
    .A1(\core.registers[1][10] ),
    .S(net963),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _14120_ (.A0(net763),
    .A1(\core.registers[1][11] ),
    .S(net963),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _14121_ (.A0(net728),
    .A1(\core.registers[1][12] ),
    .S(net963),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _14122_ (.A0(net734),
    .A1(\core.registers[1][13] ),
    .S(net963),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _14123_ (.A0(net738),
    .A1(\core.registers[1][14] ),
    .S(net961),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _14124_ (.A0(net742),
    .A1(\core.registers[1][15] ),
    .S(net962),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _14125_ (.A0(net833),
    .A1(\core.registers[1][16] ),
    .S(net962),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _14126_ (.A0(net837),
    .A1(\core.registers[1][17] ),
    .S(net961),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _14127_ (.A0(net838),
    .A1(\core.registers[1][18] ),
    .S(net963),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _14128_ (.A0(net844),
    .A1(\core.registers[1][19] ),
    .S(net961),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _14129_ (.A0(net849),
    .A1(\core.registers[1][20] ),
    .S(net961),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _14130_ (.A0(net853),
    .A1(\core.registers[1][21] ),
    .S(net961),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _14131_ (.A0(net857),
    .A1(\core.registers[1][22] ),
    .S(net962),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _14132_ (.A0(net863),
    .A1(\core.registers[1][23] ),
    .S(net961),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _14133_ (.A0(net995),
    .A1(\core.registers[1][24] ),
    .S(net961),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _14134_ (.A0(net999),
    .A1(\core.registers[1][25] ),
    .S(net961),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _14135_ (.A0(net1003),
    .A1(\core.registers[1][26] ),
    .S(net964),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _14136_ (.A0(net866),
    .A1(\core.registers[1][27] ),
    .S(net963),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _14137_ (.A0(net871),
    .A1(\core.registers[1][28] ),
    .S(net964),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _14138_ (.A0(net875),
    .A1(\core.registers[1][29] ),
    .S(net963),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _14139_ (.A0(net880),
    .A1(\core.registers[1][30] ),
    .S(net963),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _14140_ (.A0(net1023),
    .A1(\core.registers[1][31] ),
    .S(net961),
    .X(_00321_));
 sky130_fd_sc_hd__nor4_1 _14141_ (.A(_04971_),
    .B(net670),
    .C(_07600_),
    .D(_07656_),
    .Y(_08683_));
 sky130_fd_sc_hd__or4b_1 _14142_ (.A(_07683_),
    .B(_07731_),
    .C(_07780_),
    .D_N(_08683_),
    .X(_08684_));
 sky130_fd_sc_hd__or4b_2 _14143_ (.A(_07822_),
    .B(_08684_),
    .C(_07882_),
    .D_N(_07843_),
    .X(_08685_));
 sky130_fd_sc_hd__or4bb_1 _14144_ (.A(_08685_),
    .B(_08001_),
    .C_N(_07952_),
    .D_N(_07918_),
    .X(_08686_));
 sky130_fd_sc_hd__or3_1 _14145_ (.A(_08040_),
    .B(_08152_),
    .C(_08686_),
    .X(_08687_));
 sky130_fd_sc_hd__or3_1 _14146_ (.A(_08075_),
    .B(_08170_),
    .C(_08687_),
    .X(_08688_));
 sky130_fd_sc_hd__or4_2 _14147_ (.A(_08098_),
    .B(_08217_),
    .C(_08279_),
    .D(_08688_),
    .X(_08689_));
 sky130_fd_sc_hd__or2_1 _14148_ (.A(_08251_),
    .B(_08405_),
    .X(_08690_));
 sky130_fd_sc_hd__or4_2 _14149_ (.A(_08297_),
    .B(_08345_),
    .C(_08689_),
    .D(_08690_),
    .X(_08691_));
 sky130_fd_sc_hd__or2_2 _14150_ (.A(_08440_),
    .B(_08534_),
    .X(_08692_));
 sky130_fd_sc_hd__nor4_4 _14151_ (.A(_08376_),
    .B(_08470_),
    .C(_08691_),
    .D(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__nor3_4 _14152_ (.A(_08487_),
    .B(_08564_),
    .C(_08580_),
    .Y(_08694_));
 sky130_fd_sc_hd__and4_2 _14153_ (.A(net1274),
    .B(_08631_),
    .C(_08693_),
    .D(_08694_),
    .X(_08695_));
 sky130_fd_sc_hd__a31oi_4 _14154_ (.A1(_08631_),
    .A2(_08693_),
    .A3(_08694_),
    .B1(net1212),
    .Y(_08696_));
 sky130_fd_sc_hd__nor2_1 _14155_ (.A(_07366_),
    .B(net1198),
    .Y(_08697_));
 sky130_fd_sc_hd__mux2_1 _14156_ (.A0(net1206),
    .A1(net1200),
    .S(_07365_),
    .X(_08698_));
 sky130_fd_sc_hd__a211o_2 _14157_ (.A1(_07142_),
    .A2(_07366_),
    .B1(_08697_),
    .C1(_08698_),
    .X(_08699_));
 sky130_fd_sc_hd__or3_4 _14158_ (.A(_08695_),
    .B(_08696_),
    .C(_08699_),
    .X(_08700_));
 sky130_fd_sc_hd__o21ai_2 _14159_ (.A1(_06997_),
    .A2(_08700_),
    .B1(net1719),
    .Y(_08701_));
 sky130_fd_sc_hd__o211a_1 _14160_ (.A1(\core.cancelStall ),
    .A2(net1719),
    .B1(net1823),
    .C1(_08701_),
    .X(_00322_));
 sky130_fd_sc_hd__or4b_4 _14161_ (.A(\jtag.state[2] ),
    .B(net1720),
    .C(net1721),
    .D_N(\jtag.state[3] ),
    .X(_08702_));
 sky130_fd_sc_hd__nand2_2 _14162_ (.A(\jtag.tckRisingEdge ),
    .B(_06844_),
    .Y(_08703_));
 sky130_fd_sc_hd__nor2_1 _14163_ (.A(_08702_),
    .B(_08703_),
    .Y(_08704_));
 sky130_fd_sc_hd__or3_1 _14164_ (.A(\jtag.dataBSRRegister.data[26] ),
    .B(_08702_),
    .C(_08703_),
    .X(_08705_));
 sky130_fd_sc_hd__or3_4 _14165_ (.A(\jtag.managementState[0] ),
    .B(net1611),
    .C(_08705_),
    .X(_08706_));
 sky130_fd_sc_hd__mux2_1 _14166_ (.A0(\jtag.dataBSRRegister.data[0] ),
    .A1(\jtag.managementAddress[0] ),
    .S(net1176),
    .X(_08707_));
 sky130_fd_sc_hd__and2_1 _14167_ (.A(net1852),
    .B(_08707_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _14168_ (.A0(\jtag.dataBSRRegister.data[1] ),
    .A1(\jtag.managementAddress[1] ),
    .S(net1175),
    .X(_08708_));
 sky130_fd_sc_hd__and2_1 _14169_ (.A(net1852),
    .B(_08708_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _14170_ (.A0(\jtag.dataBSRRegister.data[2] ),
    .A1(\jtag.managementAddress[2] ),
    .S(net1175),
    .X(_08709_));
 sky130_fd_sc_hd__and2_1 _14171_ (.A(net1852),
    .B(_08709_),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _14172_ (.A0(\jtag.dataBSRRegister.data[3] ),
    .A1(\jtag.managementAddress[3] ),
    .S(net1175),
    .X(_08710_));
 sky130_fd_sc_hd__and2_1 _14173_ (.A(net1850),
    .B(_08710_),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _14174_ (.A0(\jtag.dataBSRRegister.data[4] ),
    .A1(\jtag.managementAddress[4] ),
    .S(net1175),
    .X(_08711_));
 sky130_fd_sc_hd__and2_1 _14175_ (.A(net1850),
    .B(_08711_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _14176_ (.A0(\jtag.dataBSRRegister.data[5] ),
    .A1(\jtag.managementAddress[5] ),
    .S(net1175),
    .X(_08712_));
 sky130_fd_sc_hd__and2_1 _14177_ (.A(net1839),
    .B(_08712_),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _14178_ (.A0(\jtag.dataBSRRegister.data[6] ),
    .A1(\jtag.managementAddress[6] ),
    .S(net1175),
    .X(_08713_));
 sky130_fd_sc_hd__and2_1 _14179_ (.A(net1840),
    .B(_08713_),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _14180_ (.A0(\jtag.dataBSRRegister.data[7] ),
    .A1(\jtag.managementAddress[7] ),
    .S(net1175),
    .X(_08714_));
 sky130_fd_sc_hd__and2_1 _14181_ (.A(net1842),
    .B(_08714_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _14182_ (.A0(\jtag.dataBSRRegister.data[8] ),
    .A1(\jtag.managementAddress[8] ),
    .S(net1176),
    .X(_08715_));
 sky130_fd_sc_hd__and2_1 _14183_ (.A(net1856),
    .B(_08715_),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _14184_ (.A0(\jtag.dataBSRRegister.data[9] ),
    .A1(\jtag.managementAddress[9] ),
    .S(net1175),
    .X(_08716_));
 sky130_fd_sc_hd__and2_1 _14185_ (.A(net1864),
    .B(_08716_),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _14186_ (.A0(\jtag.dataBSRRegister.data[10] ),
    .A1(\jtag.managementAddress[10] ),
    .S(net1175),
    .X(_08717_));
 sky130_fd_sc_hd__and2_1 _14187_ (.A(net1864),
    .B(_08717_),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _14188_ (.A0(\jtag.dataBSRRegister.data[11] ),
    .A1(\jtag.managementAddress[11] ),
    .S(net1176),
    .X(_08718_));
 sky130_fd_sc_hd__and2_1 _14189_ (.A(net1864),
    .B(_08718_),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _14190_ (.A0(\jtag.dataBSRRegister.data[12] ),
    .A1(\jtag.managementAddress[12] ),
    .S(net1176),
    .X(_08719_));
 sky130_fd_sc_hd__and2_1 _14191_ (.A(net1865),
    .B(_08719_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _14192_ (.A0(\jtag.dataBSRRegister.data[13] ),
    .A1(\jtag.managementAddress[13] ),
    .S(net1176),
    .X(_08720_));
 sky130_fd_sc_hd__and2_1 _14193_ (.A(net1865),
    .B(_08720_),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _14194_ (.A0(\jtag.dataBSRRegister.data[14] ),
    .A1(\jtag.managementAddress[14] ),
    .S(net1176),
    .X(_08721_));
 sky130_fd_sc_hd__and2_1 _14195_ (.A(net1857),
    .B(_08721_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _14196_ (.A0(\jtag.dataBSRRegister.data[15] ),
    .A1(\jtag.managementAddress[15] ),
    .S(net1176),
    .X(_08722_));
 sky130_fd_sc_hd__and2_1 _14197_ (.A(net1857),
    .B(_08722_),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _14198_ (.A0(\jtag.dataBSRRegister.data[16] ),
    .A1(\jtag.managementAddress[16] ),
    .S(net1176),
    .X(_08723_));
 sky130_fd_sc_hd__and2_1 _14199_ (.A(net1860),
    .B(_08723_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _14200_ (.A0(\jtag.dataBSRRegister.data[17] ),
    .A1(\jtag.managementAddress[17] ),
    .S(net1176),
    .X(_08724_));
 sky130_fd_sc_hd__and2_1 _14201_ (.A(net1860),
    .B(_08724_),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _14202_ (.A0(\jtag.dataBSRRegister.data[18] ),
    .A1(\jtag.managementAddress[18] ),
    .S(_08706_),
    .X(_08725_));
 sky130_fd_sc_hd__and2_1 _14203_ (.A(net1860),
    .B(_08725_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _14204_ (.A0(\jtag.dataBSRRegister.data[19] ),
    .A1(\jtag.managementAddress[19] ),
    .S(_08706_),
    .X(_08726_));
 sky130_fd_sc_hd__and2_1 _14205_ (.A(net1859),
    .B(_08726_),
    .X(_00342_));
 sky130_fd_sc_hd__or2_1 _14206_ (.A(net450),
    .B(net599),
    .X(_08727_));
 sky130_fd_sc_hd__o211a_1 _14207_ (.A1(\core.pipe0_fetch.lastProgramCounter[0] ),
    .A2(net594),
    .B1(_08727_),
    .C1(net1820),
    .X(_00343_));
 sky130_fd_sc_hd__or2_1 _14208_ (.A(net461),
    .B(net599),
    .X(_08728_));
 sky130_fd_sc_hd__o211a_1 _14209_ (.A1(\core.pipe0_fetch.lastProgramCounter[1] ),
    .A2(net592),
    .B1(_08728_),
    .C1(net1806),
    .X(_00344_));
 sky130_fd_sc_hd__nand2_1 _14210_ (.A(_03827_),
    .B(net595),
    .Y(_08729_));
 sky130_fd_sc_hd__o211a_1 _14211_ (.A1(\core.pipe0_fetch.lastProgramCounter[2] ),
    .A2(net595),
    .B1(_08729_),
    .C1(net1802),
    .X(_00345_));
 sky130_fd_sc_hd__or2_1 _14212_ (.A(net475),
    .B(net601),
    .X(_08730_));
 sky130_fd_sc_hd__o211a_1 _14213_ (.A1(\core.pipe0_fetch.lastProgramCounter[3] ),
    .A2(net595),
    .B1(_08730_),
    .C1(net1802),
    .X(_00346_));
 sky130_fd_sc_hd__or2_1 _14214_ (.A(net1748),
    .B(net601),
    .X(_08731_));
 sky130_fd_sc_hd__o211a_1 _14215_ (.A1(\core.pipe0_fetch.lastProgramCounter[4] ),
    .A2(net595),
    .B1(_08731_),
    .C1(net1802),
    .X(_00347_));
 sky130_fd_sc_hd__or2_1 _14216_ (.A(net477),
    .B(net601),
    .X(_08732_));
 sky130_fd_sc_hd__o211a_1 _14217_ (.A1(\core.pipe0_fetch.lastProgramCounter[5] ),
    .A2(net595),
    .B1(_08732_),
    .C1(net1802),
    .X(_00348_));
 sky130_fd_sc_hd__or2_1 _14218_ (.A(net478),
    .B(net601),
    .X(_08733_));
 sky130_fd_sc_hd__o211a_1 _14219_ (.A1(\core.pipe0_fetch.lastProgramCounter[6] ),
    .A2(net592),
    .B1(_08733_),
    .C1(net1803),
    .X(_00349_));
 sky130_fd_sc_hd__nand2_1 _14220_ (.A(_03826_),
    .B(net596),
    .Y(_08734_));
 sky130_fd_sc_hd__o211a_1 _14221_ (.A1(\core.pipe0_fetch.lastProgramCounter[7] ),
    .A2(net596),
    .B1(_08734_),
    .C1(net1830),
    .X(_00350_));
 sky130_fd_sc_hd__or2_1 _14222_ (.A(net480),
    .B(net600),
    .X(_08735_));
 sky130_fd_sc_hd__o211a_1 _14223_ (.A1(\core.pipe0_fetch.lastProgramCounter[8] ),
    .A2(net593),
    .B1(_08735_),
    .C1(net1812),
    .X(_00351_));
 sky130_fd_sc_hd__nand2_1 _14224_ (.A(_03825_),
    .B(net596),
    .Y(_08736_));
 sky130_fd_sc_hd__o211a_1 _14225_ (.A1(\core.pipe0_fetch.lastProgramCounter[9] ),
    .A2(net596),
    .B1(_08736_),
    .C1(net1825),
    .X(_00352_));
 sky130_fd_sc_hd__or2_1 _14226_ (.A(net451),
    .B(net601),
    .X(_08737_));
 sky130_fd_sc_hd__o211a_1 _14227_ (.A1(\core.pipe0_fetch.lastProgramCounter[10] ),
    .A2(net592),
    .B1(_08737_),
    .C1(net1806),
    .X(_00353_));
 sky130_fd_sc_hd__or2_1 _14228_ (.A(net452),
    .B(net599),
    .X(_08738_));
 sky130_fd_sc_hd__o211a_1 _14229_ (.A1(\core.pipe0_fetch.lastProgramCounter[11] ),
    .A2(net594),
    .B1(_08738_),
    .C1(net1811),
    .X(_00354_));
 sky130_fd_sc_hd__or2_1 _14230_ (.A(net453),
    .B(net600),
    .X(_08739_));
 sky130_fd_sc_hd__o211a_1 _14231_ (.A1(\core.pipe0_fetch.lastProgramCounter[12] ),
    .A2(net594),
    .B1(_08739_),
    .C1(net1812),
    .X(_00355_));
 sky130_fd_sc_hd__or2_1 _14232_ (.A(net454),
    .B(net600),
    .X(_08740_));
 sky130_fd_sc_hd__o211a_1 _14233_ (.A1(\core.pipe0_fetch.lastProgramCounter[13] ),
    .A2(net593),
    .B1(_08740_),
    .C1(net1811),
    .X(_00356_));
 sky130_fd_sc_hd__or2_1 _14234_ (.A(net455),
    .B(net600),
    .X(_08741_));
 sky130_fd_sc_hd__o211a_1 _14235_ (.A1(\core.pipe0_fetch.lastProgramCounter[14] ),
    .A2(net593),
    .B1(_08741_),
    .C1(net1807),
    .X(_00357_));
 sky130_fd_sc_hd__or2_1 _14236_ (.A(net456),
    .B(net599),
    .X(_08742_));
 sky130_fd_sc_hd__o211a_1 _14237_ (.A1(\core.pipe0_fetch.lastProgramCounter[15] ),
    .A2(net593),
    .B1(_08742_),
    .C1(net1807),
    .X(_00358_));
 sky130_fd_sc_hd__or2_1 _14238_ (.A(net1747),
    .B(net599),
    .X(_08743_));
 sky130_fd_sc_hd__o211a_1 _14239_ (.A1(\core.pipe0_fetch.lastProgramCounter[16] ),
    .A2(net592),
    .B1(_08743_),
    .C1(net1806),
    .X(_00359_));
 sky130_fd_sc_hd__or2_1 _14240_ (.A(net458),
    .B(net601),
    .X(_08744_));
 sky130_fd_sc_hd__o211a_1 _14241_ (.A1(\core.pipe0_fetch.lastProgramCounter[17] ),
    .A2(net592),
    .B1(_08744_),
    .C1(net1806),
    .X(_00360_));
 sky130_fd_sc_hd__or2_1 _14242_ (.A(net459),
    .B(net601),
    .X(_08745_));
 sky130_fd_sc_hd__o211a_1 _14243_ (.A1(\core.pipe0_fetch.lastProgramCounter[18] ),
    .A2(net592),
    .B1(_08745_),
    .C1(net1806),
    .X(_00361_));
 sky130_fd_sc_hd__or2_1 _14244_ (.A(net460),
    .B(net601),
    .X(_08746_));
 sky130_fd_sc_hd__o211a_1 _14245_ (.A1(\core.pipe0_fetch.lastProgramCounter[19] ),
    .A2(net592),
    .B1(_08746_),
    .C1(net1809),
    .X(_00362_));
 sky130_fd_sc_hd__or2_1 _14246_ (.A(net462),
    .B(net599),
    .X(_08747_));
 sky130_fd_sc_hd__o211a_1 _14247_ (.A1(\core.pipe0_fetch.lastProgramCounter[20] ),
    .A2(net594),
    .B1(_08747_),
    .C1(net1809),
    .X(_00363_));
 sky130_fd_sc_hd__or2_1 _14248_ (.A(net463),
    .B(net599),
    .X(_08748_));
 sky130_fd_sc_hd__o211a_1 _14249_ (.A1(\core.pipe0_fetch.lastProgramCounter[21] ),
    .A2(net593),
    .B1(_08748_),
    .C1(net1807),
    .X(_00364_));
 sky130_fd_sc_hd__or2_1 _14250_ (.A(net464),
    .B(net600),
    .X(_08749_));
 sky130_fd_sc_hd__o211a_1 _14251_ (.A1(\core.pipe0_fetch.lastProgramCounter[22] ),
    .A2(net593),
    .B1(_08749_),
    .C1(net1808),
    .X(_00365_));
 sky130_fd_sc_hd__nand2_1 _14252_ (.A(_03824_),
    .B(net595),
    .Y(_08750_));
 sky130_fd_sc_hd__o211a_1 _14253_ (.A1(\core.pipe0_fetch.lastProgramCounter[23] ),
    .A2(net595),
    .B1(_08750_),
    .C1(net1810),
    .X(_00366_));
 sky130_fd_sc_hd__or2_1 _14254_ (.A(net466),
    .B(net600),
    .X(_08751_));
 sky130_fd_sc_hd__o211a_1 _14255_ (.A1(\core.pipe0_fetch.lastProgramCounter[24] ),
    .A2(net593),
    .B1(_08751_),
    .C1(net1811),
    .X(_00367_));
 sky130_fd_sc_hd__or2_1 _14256_ (.A(net467),
    .B(net600),
    .X(_08752_));
 sky130_fd_sc_hd__o211a_1 _14257_ (.A1(\core.pipe0_fetch.lastProgramCounter[25] ),
    .A2(net593),
    .B1(_08752_),
    .C1(net1811),
    .X(_00368_));
 sky130_fd_sc_hd__or2_1 _14258_ (.A(net468),
    .B(net600),
    .X(_08753_));
 sky130_fd_sc_hd__o211a_1 _14259_ (.A1(\core.pipe0_fetch.lastProgramCounter[26] ),
    .A2(net593),
    .B1(_08753_),
    .C1(net1807),
    .X(_00369_));
 sky130_fd_sc_hd__or2_1 _14260_ (.A(net469),
    .B(net600),
    .X(_08754_));
 sky130_fd_sc_hd__o211a_1 _14261_ (.A1(\core.pipe0_fetch.lastProgramCounter[27] ),
    .A2(net593),
    .B1(_08754_),
    .C1(net1811),
    .X(_00370_));
 sky130_fd_sc_hd__or2_1 _14262_ (.A(net470),
    .B(net599),
    .X(_08755_));
 sky130_fd_sc_hd__o211a_1 _14263_ (.A1(\core.pipe0_fetch.lastProgramCounter[28] ),
    .A2(net592),
    .B1(_08755_),
    .C1(net1807),
    .X(_00371_));
 sky130_fd_sc_hd__or2_1 _14264_ (.A(net471),
    .B(net599),
    .X(_08756_));
 sky130_fd_sc_hd__o211a_1 _14265_ (.A1(\core.pipe0_fetch.lastProgramCounter[29] ),
    .A2(net592),
    .B1(_08756_),
    .C1(net1807),
    .X(_00372_));
 sky130_fd_sc_hd__or2_1 _14266_ (.A(net473),
    .B(net599),
    .X(_08757_));
 sky130_fd_sc_hd__o211a_1 _14267_ (.A1(\core.pipe0_fetch.lastProgramCounter[30] ),
    .A2(net592),
    .B1(_08757_),
    .C1(net1809),
    .X(_00373_));
 sky130_fd_sc_hd__nand2_1 _14268_ (.A(_03823_),
    .B(net598),
    .Y(_08758_));
 sky130_fd_sc_hd__o211a_1 _14269_ (.A1(\core.pipe0_fetch.lastProgramCounter[31] ),
    .A2(net598),
    .B1(_08758_),
    .C1(net1814),
    .X(_00374_));
 sky130_fd_sc_hd__and3b_2 _14270_ (.A_N(net1801),
    .B(_03904_),
    .C(\core.csr.currentInstruction[10] ),
    .X(_08759_));
 sky130_fd_sc_hd__or2_4 _14271_ (.A(\core.csr.currentInstruction[7] ),
    .B(_06850_),
    .X(_08760_));
 sky130_fd_sc_hd__nor2_8 _14272_ (.A(_03909_),
    .B(_06850_),
    .Y(_08761_));
 sky130_fd_sc_hd__nand2_2 _14273_ (.A(_08759_),
    .B(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__mux2_1 _14274_ (.A0(net1077),
    .A1(\core.registers[26][0] ),
    .S(net824),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _14275_ (.A0(net1080),
    .A1(\core.registers[26][1] ),
    .S(net824),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _14276_ (.A0(net1088),
    .A1(\core.registers[26][2] ),
    .S(net823),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _14277_ (.A0(net1089),
    .A1(\core.registers[26][3] ),
    .S(net824),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _14278_ (.A0(net1029),
    .A1(\core.registers[26][4] ),
    .S(net822),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _14279_ (.A0(net1032),
    .A1(\core.registers[26][5] ),
    .S(net823),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _14280_ (.A0(net1038),
    .A1(\core.registers[26][6] ),
    .S(net823),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _14281_ (.A0(net1137),
    .A1(\core.registers[26][7] ),
    .S(net822),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _14282_ (.A0(net897),
    .A1(\core.registers[26][8] ),
    .S(net823),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _14283_ (.A0(net900),
    .A1(\core.registers[26][9] ),
    .S(net822),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _14284_ (.A0(net757),
    .A1(\core.registers[26][10] ),
    .S(net822),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _14285_ (.A0(net764),
    .A1(\core.registers[26][11] ),
    .S(net822),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _14286_ (.A0(net731),
    .A1(\core.registers[26][12] ),
    .S(net822),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _14287_ (.A0(net735),
    .A1(\core.registers[26][13] ),
    .S(net823),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _14288_ (.A0(net737),
    .A1(\core.registers[26][14] ),
    .S(net821),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _14289_ (.A0(net741),
    .A1(\core.registers[26][15] ),
    .S(net823),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _14290_ (.A0(net831),
    .A1(\core.registers[26][16] ),
    .S(net823),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _14291_ (.A0(net834),
    .A1(\core.registers[26][17] ),
    .S(net821),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _14292_ (.A0(net841),
    .A1(\core.registers[26][18] ),
    .S(net822),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _14293_ (.A0(net842),
    .A1(\core.registers[26][19] ),
    .S(net821),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _14294_ (.A0(net846),
    .A1(\core.registers[26][20] ),
    .S(net821),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _14295_ (.A0(net850),
    .A1(\core.registers[26][21] ),
    .S(net821),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _14296_ (.A0(net855),
    .A1(\core.registers[26][22] ),
    .S(net823),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _14297_ (.A0(net860),
    .A1(\core.registers[26][23] ),
    .S(net821),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _14298_ (.A0(net992),
    .A1(\core.registers[26][24] ),
    .S(net821),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _14299_ (.A0(net997),
    .A1(\core.registers[26][25] ),
    .S(net821),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _14300_ (.A0(net1000),
    .A1(\core.registers[26][26] ),
    .S(net821),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _14301_ (.A0(net864),
    .A1(\core.registers[26][27] ),
    .S(net823),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _14302_ (.A0(net870),
    .A1(\core.registers[26][28] ),
    .S(net822),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _14303_ (.A0(net873),
    .A1(\core.registers[26][29] ),
    .S(net822),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _14304_ (.A0(net877),
    .A1(\core.registers[26][30] ),
    .S(net822),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _14305_ (.A0(net1026),
    .A1(\core.registers[26][31] ),
    .S(net821),
    .X(_00406_));
 sky130_fd_sc_hd__or3_4 _14306_ (.A(\core.csr.currentInstruction[11] ),
    .B(net1801),
    .C(_03907_),
    .X(_08763_));
 sky130_fd_sc_hd__nor2_2 _14307_ (.A(_06852_),
    .B(_08763_),
    .Y(_08764_));
 sky130_fd_sc_hd__mux2_1 _14308_ (.A0(\core.registers[11][0] ),
    .A1(net1077),
    .S(net820),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _14309_ (.A0(\core.registers[11][1] ),
    .A1(net1080),
    .S(net818),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _14310_ (.A0(\core.registers[11][2] ),
    .A1(net1085),
    .S(net817),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _14311_ (.A0(\core.registers[11][3] ),
    .A1(net1090),
    .S(net820),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _14312_ (.A0(\core.registers[11][4] ),
    .A1(net1029),
    .S(net818),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _14313_ (.A0(\core.registers[11][5] ),
    .A1(net1031),
    .S(net818),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _14314_ (.A0(\core.registers[11][6] ),
    .A1(net1036),
    .S(net818),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _14315_ (.A0(\core.registers[11][7] ),
    .A1(net1139),
    .S(net818),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _14316_ (.A0(\core.registers[11][8] ),
    .A1(net896),
    .S(net818),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _14317_ (.A0(\core.registers[11][9] ),
    .A1(net900),
    .S(net819),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _14318_ (.A0(\core.registers[11][10] ),
    .A1(net757),
    .S(net818),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _14319_ (.A0(\core.registers[11][11] ),
    .A1(net761),
    .S(net819),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _14320_ (.A0(\core.registers[11][12] ),
    .A1(net728),
    .S(net819),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _14321_ (.A0(\core.registers[11][13] ),
    .A1(net732),
    .S(net819),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _14322_ (.A0(\core.registers[11][14] ),
    .A1(net736),
    .S(net817),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _14323_ (.A0(\core.registers[11][15] ),
    .A1(net740),
    .S(net820),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _14324_ (.A0(\core.registers[11][16] ),
    .A1(net832),
    .S(net818),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _14325_ (.A0(\core.registers[11][17] ),
    .A1(net835),
    .S(net820),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _14326_ (.A0(\core.registers[11][18] ),
    .A1(net840),
    .S(net819),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _14327_ (.A0(\core.registers[11][19] ),
    .A1(net843),
    .S(net817),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _14328_ (.A0(\core.registers[11][20] ),
    .A1(net847),
    .S(net817),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _14329_ (.A0(\core.registers[11][21] ),
    .A1(net850),
    .S(net817),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _14330_ (.A0(\core.registers[11][22] ),
    .A1(net855),
    .S(net818),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _14331_ (.A0(\core.registers[11][23] ),
    .A1(net860),
    .S(net817),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _14332_ (.A0(\core.registers[11][24] ),
    .A1(net992),
    .S(net817),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _14333_ (.A0(\core.registers[11][25] ),
    .A1(net996),
    .S(net817),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _14334_ (.A0(\core.registers[11][26] ),
    .A1(net1000),
    .S(net817),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _14335_ (.A0(\core.registers[11][27] ),
    .A1(net865),
    .S(net818),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _14336_ (.A0(\core.registers[11][28] ),
    .A1(net869),
    .S(net819),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _14337_ (.A0(\core.registers[11][29] ),
    .A1(net873),
    .S(net819),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _14338_ (.A0(\core.registers[11][30] ),
    .A1(net880),
    .S(net819),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _14339_ (.A0(\core.registers[11][31] ),
    .A1(net1026),
    .S(net817),
    .X(_00438_));
 sky130_fd_sc_hd__nand2_1 _14340_ (.A(net1823),
    .B(_06691_),
    .Y(_08765_));
 sky130_fd_sc_hd__inv_2 _14341_ (.A(_08765_),
    .Y(_00510_));
 sky130_fd_sc_hd__and3_4 _14342_ (.A(net1824),
    .B(_06691_),
    .C(_06830_),
    .X(_00439_));
 sky130_fd_sc_hd__and3_4 _14343_ (.A(net1805),
    .B(_06691_),
    .C(_06831_),
    .X(_00440_));
 sky130_fd_sc_hd__and3_4 _14344_ (.A(net1805),
    .B(_06691_),
    .C(_06832_),
    .X(_00441_));
 sky130_fd_sc_hd__and3_4 _14345_ (.A(net1805),
    .B(_06691_),
    .C(_06833_),
    .X(_00442_));
 sky130_fd_sc_hd__nor2_1 _14346_ (.A(net1906),
    .B(_03876_),
    .Y(_00443_));
 sky130_fd_sc_hd__nor2_4 _14347_ (.A(net1879),
    .B(_06654_),
    .Y(_00444_));
 sky130_fd_sc_hd__nor2_1 _14348_ (.A(_03821_),
    .B(net1871),
    .Y(_00545_));
 sky130_fd_sc_hd__and2_2 _14349_ (.A(net1830),
    .B(net1313),
    .X(_00445_));
 sky130_fd_sc_hd__or3_4 _14350_ (.A(_03903_),
    .B(_03904_),
    .C(_03906_),
    .X(_08766_));
 sky130_fd_sc_hd__nor2_8 _14351_ (.A(_06852_),
    .B(_08766_),
    .Y(_08767_));
 sky130_fd_sc_hd__mux2_1 _14352_ (.A0(\core.registers[7][0] ),
    .A1(net1078),
    .S(net813),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _14353_ (.A0(\core.registers[7][1] ),
    .A1(net1081),
    .S(net816),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _14354_ (.A0(\core.registers[7][2] ),
    .A1(net1086),
    .S(net814),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _14355_ (.A0(\core.registers[7][3] ),
    .A1(net1092),
    .S(net813),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _14356_ (.A0(\core.registers[7][4] ),
    .A1(net1028),
    .S(net816),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _14357_ (.A0(\core.registers[7][5] ),
    .A1(net1033),
    .S(net814),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _14358_ (.A0(\core.registers[7][6] ),
    .A1(net1035),
    .S(net814),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _14359_ (.A0(\core.registers[7][7] ),
    .A1(net1140),
    .S(net816),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _14360_ (.A0(\core.registers[7][8] ),
    .A1(net898),
    .S(net815),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _14361_ (.A0(\core.registers[7][9] ),
    .A1(net902),
    .S(net815),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _14362_ (.A0(\core.registers[7][10] ),
    .A1(net759),
    .S(net815),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _14363_ (.A0(\core.registers[7][11] ),
    .A1(net762),
    .S(net815),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _14364_ (.A0(\core.registers[7][12] ),
    .A1(net729),
    .S(net815),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _14365_ (.A0(\core.registers[7][13] ),
    .A1(net733),
    .S(net815),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _14366_ (.A0(\core.registers[7][14] ),
    .A1(net738),
    .S(net813),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _14367_ (.A0(\core.registers[7][15] ),
    .A1(net742),
    .S(net814),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _14368_ (.A0(\core.registers[7][16] ),
    .A1(net832),
    .S(net814),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _14369_ (.A0(\core.registers[7][17] ),
    .A1(net837),
    .S(net813),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _14370_ (.A0(\core.registers[7][18] ),
    .A1(net839),
    .S(net816),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _14371_ (.A0(\core.registers[7][19] ),
    .A1(net844),
    .S(net813),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _14372_ (.A0(\core.registers[7][20] ),
    .A1(net848),
    .S(net813),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _14373_ (.A0(\core.registers[7][21] ),
    .A1(net852),
    .S(net813),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _14374_ (.A0(\core.registers[7][22] ),
    .A1(net857),
    .S(net814),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _14375_ (.A0(\core.registers[7][23] ),
    .A1(net863),
    .S(net813),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _14376_ (.A0(\core.registers[7][24] ),
    .A1(net995),
    .S(net813),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _14377_ (.A0(\core.registers[7][25] ),
    .A1(net998),
    .S(net814),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _14378_ (.A0(\core.registers[7][26] ),
    .A1(net1002),
    .S(net815),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _14379_ (.A0(\core.registers[7][27] ),
    .A1(net866),
    .S(net815),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _14380_ (.A0(\core.registers[7][28] ),
    .A1(net871),
    .S(net816),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _14381_ (.A0(\core.registers[7][29] ),
    .A1(net875),
    .S(net815),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _14382_ (.A0(\core.registers[7][30] ),
    .A1(net879),
    .S(net815),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _14383_ (.A0(\core.registers[7][31] ),
    .A1(net1024),
    .S(net813),
    .X(_00477_));
 sky130_fd_sc_hd__or4b_4 _14384_ (.A(_03909_),
    .B(_06849_),
    .C(_08763_),
    .D_N(_03911_),
    .X(_08768_));
 sky130_fd_sc_hd__mux2_1 _14385_ (.A0(net1076),
    .A1(\core.registers[8][0] ),
    .S(net1018),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _14386_ (.A0(net1080),
    .A1(\core.registers[8][1] ),
    .S(net1017),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _14387_ (.A0(net1086),
    .A1(\core.registers[8][2] ),
    .S(net1018),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _14388_ (.A0(net1089),
    .A1(\core.registers[8][3] ),
    .S(net1015),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _14389_ (.A0(net1029),
    .A1(\core.registers[8][4] ),
    .S(net1017),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _14390_ (.A0(net1031),
    .A1(\core.registers[8][5] ),
    .S(net1017),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _14391_ (.A0(net1038),
    .A1(\core.registers[8][6] ),
    .S(net1017),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _14392_ (.A0(net1137),
    .A1(\core.registers[8][7] ),
    .S(net1017),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _14393_ (.A0(net896),
    .A1(\core.registers[8][8] ),
    .S(net1016),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _14394_ (.A0(net903),
    .A1(\core.registers[8][9] ),
    .S(net1016),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _14395_ (.A0(net760),
    .A1(\core.registers[8][10] ),
    .S(net1016),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _14396_ (.A0(net763),
    .A1(\core.registers[8][11] ),
    .S(net1016),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _14397_ (.A0(net728),
    .A1(\core.registers[8][12] ),
    .S(net1016),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _14398_ (.A0(net732),
    .A1(\core.registers[8][13] ),
    .S(net1016),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _14399_ (.A0(net736),
    .A1(\core.registers[8][14] ),
    .S(net1015),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _14400_ (.A0(net740),
    .A1(\core.registers[8][15] ),
    .S(net1018),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _14401_ (.A0(net832),
    .A1(\core.registers[8][16] ),
    .S(net1017),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _14402_ (.A0(net834),
    .A1(\core.registers[8][17] ),
    .S(net1018),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _14403_ (.A0(net840),
    .A1(\core.registers[8][18] ),
    .S(net1016),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _14404_ (.A0(net843),
    .A1(\core.registers[8][19] ),
    .S(net1015),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _14405_ (.A0(net847),
    .A1(\core.registers[8][20] ),
    .S(net1015),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _14406_ (.A0(net850),
    .A1(\core.registers[8][21] ),
    .S(net1015),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _14407_ (.A0(net856),
    .A1(\core.registers[8][22] ),
    .S(net1017),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _14408_ (.A0(net860),
    .A1(\core.registers[8][23] ),
    .S(net1015),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _14409_ (.A0(net992),
    .A1(\core.registers[8][24] ),
    .S(net1015),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _14410_ (.A0(net996),
    .A1(\core.registers[8][25] ),
    .S(net1015),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _14411_ (.A0(net1000),
    .A1(\core.registers[8][26] ),
    .S(net1015),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _14412_ (.A0(net864),
    .A1(\core.registers[8][27] ),
    .S(net1017),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _14413_ (.A0(net870),
    .A1(\core.registers[8][28] ),
    .S(net1016),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _14414_ (.A0(net876),
    .A1(\core.registers[8][29] ),
    .S(net1016),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _14415_ (.A0(net877),
    .A1(\core.registers[8][30] ),
    .S(net1016),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _14416_ (.A0(net1026),
    .A1(\core.registers[8][31] ),
    .S(net1015),
    .X(_00509_));
 sky130_fd_sc_hd__and3_4 _14417_ (.A(net1837),
    .B(_06701_),
    .C(_06703_),
    .X(_00516_));
 sky130_fd_sc_hd__and3_1 _14418_ (.A(\wbSRAMInterface.currentByteSelect[0] ),
    .B(net1614),
    .C(_00516_),
    .X(_00511_));
 sky130_fd_sc_hd__and3_1 _14419_ (.A(\wbSRAMInterface.currentByteSelect[1] ),
    .B(net1614),
    .C(_00516_),
    .X(_00512_));
 sky130_fd_sc_hd__and3_1 _14420_ (.A(\wbSRAMInterface.currentByteSelect[2] ),
    .B(net1614),
    .C(_00516_),
    .X(_00513_));
 sky130_fd_sc_hd__and3_1 _14421_ (.A(\wbSRAMInterface.currentByteSelect[3] ),
    .B(net1614),
    .C(_00516_),
    .X(_00514_));
 sky130_fd_sc_hd__and2b_1 _14422_ (.A_N(_06706_),
    .B(_00516_),
    .X(_00515_));
 sky130_fd_sc_hd__nor2_4 _14423_ (.A(_03815_),
    .B(net1879),
    .Y(_00517_));
 sky130_fd_sc_hd__nor2_4 _14424_ (.A(_03814_),
    .B(net1875),
    .Y(_00518_));
 sky130_fd_sc_hd__and2_1 _14425_ (.A(\core.fetchProgramCounter[2] ),
    .B(net1804),
    .X(_00519_));
 sky130_fd_sc_hd__and2_1 _14426_ (.A(\core.fetchProgramCounter[3] ),
    .B(net1802),
    .X(_00520_));
 sky130_fd_sc_hd__and2_1 _14427_ (.A(\core.fetchProgramCounter[4] ),
    .B(net1804),
    .X(_00521_));
 sky130_fd_sc_hd__and2_1 _14428_ (.A(\core.fetchProgramCounter[5] ),
    .B(net1802),
    .X(_00522_));
 sky130_fd_sc_hd__and2_1 _14429_ (.A(\core.fetchProgramCounter[6] ),
    .B(net1803),
    .X(_00523_));
 sky130_fd_sc_hd__and2_1 _14430_ (.A(\core.fetchProgramCounter[7] ),
    .B(net1830),
    .X(_00524_));
 sky130_fd_sc_hd__and2_1 _14431_ (.A(\core.fetchProgramCounter[8] ),
    .B(net1811),
    .X(_00525_));
 sky130_fd_sc_hd__and2_1 _14432_ (.A(\core.fetchProgramCounter[9] ),
    .B(net1825),
    .X(_00526_));
 sky130_fd_sc_hd__and2_1 _14433_ (.A(\core.fetchProgramCounter[10] ),
    .B(net1803),
    .X(_00527_));
 sky130_fd_sc_hd__and2_1 _14434_ (.A(\core.fetchProgramCounter[11] ),
    .B(net1807),
    .X(_00528_));
 sky130_fd_sc_hd__and2_2 _14435_ (.A(\core.fetchProgramCounter[12] ),
    .B(net1828),
    .X(_00529_));
 sky130_fd_sc_hd__and2_1 _14436_ (.A(\core.fetchProgramCounter[13] ),
    .B(net1811),
    .X(_00530_));
 sky130_fd_sc_hd__and2_1 _14437_ (.A(\core.fetchProgramCounter[14] ),
    .B(net1807),
    .X(_00531_));
 sky130_fd_sc_hd__and2_1 _14438_ (.A(\core.fetchProgramCounter[15] ),
    .B(net1807),
    .X(_00532_));
 sky130_fd_sc_hd__and2_2 _14439_ (.A(\core.fetchProgramCounter[16] ),
    .B(net1815),
    .X(_00533_));
 sky130_fd_sc_hd__and2_1 _14440_ (.A(\core.fetchProgramCounter[17] ),
    .B(net1806),
    .X(_00534_));
 sky130_fd_sc_hd__and2_1 _14441_ (.A(\core.fetchProgramCounter[18] ),
    .B(net1806),
    .X(_00535_));
 sky130_fd_sc_hd__and2_1 _14442_ (.A(\core.fetchProgramCounter[19] ),
    .B(net1809),
    .X(_00536_));
 sky130_fd_sc_hd__and2_1 _14443_ (.A(\core.fetchProgramCounter[20] ),
    .B(net1806),
    .X(_00537_));
 sky130_fd_sc_hd__and2_1 _14444_ (.A(\core.fetchProgramCounter[21] ),
    .B(net1806),
    .X(_00538_));
 sky130_fd_sc_hd__and2_1 _14445_ (.A(\core.fetchProgramCounter[22] ),
    .B(net1808),
    .X(_00539_));
 sky130_fd_sc_hd__and2_1 _14446_ (.A(\core.fetchProgramCounter[23] ),
    .B(net1810),
    .X(_00540_));
 sky130_fd_sc_hd__and2_1 _14447_ (.A(\core.fetchProgramCounter[24] ),
    .B(net1811),
    .X(_00541_));
 sky130_fd_sc_hd__and2_1 _14448_ (.A(\core.fetchProgramCounter[25] ),
    .B(net1811),
    .X(_00542_));
 sky130_fd_sc_hd__and2_1 _14449_ (.A(\core.fetchProgramCounter[26] ),
    .B(net1808),
    .X(_00543_));
 sky130_fd_sc_hd__and2_1 _14450_ (.A(\core.fetchProgramCounter[27] ),
    .B(net1811),
    .X(_00544_));
 sky130_fd_sc_hd__and2_1 _14451_ (.A(\core.fetchProgramCounter[29] ),
    .B(net1807),
    .X(_00546_));
 sky130_fd_sc_hd__and2_1 _14452_ (.A(\core.fetchProgramCounter[30] ),
    .B(net1806),
    .X(_00547_));
 sky130_fd_sc_hd__and2_1 _14453_ (.A(\core.fetchProgramCounter[31] ),
    .B(net1814),
    .X(_00548_));
 sky130_fd_sc_hd__nor2_8 _14454_ (.A(_06853_),
    .B(_08760_),
    .Y(_08769_));
 sky130_fd_sc_hd__mux2_1 _14455_ (.A0(\core.registers[18][0] ),
    .A1(net1078),
    .S(net810),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _14456_ (.A0(\core.registers[18][1] ),
    .A1(net1083),
    .S(net812),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _14457_ (.A0(\core.registers[18][2] ),
    .A1(net1085),
    .S(net810),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _14458_ (.A0(\core.registers[18][3] ),
    .A1(net1090),
    .S(net809),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _14459_ (.A0(\core.registers[18][4] ),
    .A1(net1028),
    .S(net812),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _14460_ (.A0(\core.registers[18][5] ),
    .A1(net1033),
    .S(net812),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _14461_ (.A0(\core.registers[18][6] ),
    .A1(net1037),
    .S(net812),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _14462_ (.A0(\core.registers[18][7] ),
    .A1(net1138),
    .S(net812),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _14463_ (.A0(\core.registers[18][8] ),
    .A1(net898),
    .S(net811),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _14464_ (.A0(\core.registers[18][9] ),
    .A1(net900),
    .S(net811),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _14465_ (.A0(\core.registers[18][10] ),
    .A1(net760),
    .S(net811),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _14466_ (.A0(\core.registers[18][11] ),
    .A1(net761),
    .S(net811),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _14467_ (.A0(\core.registers[18][12] ),
    .A1(net729),
    .S(net812),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _14468_ (.A0(\core.registers[18][13] ),
    .A1(net733),
    .S(net811),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _14469_ (.A0(\core.registers[18][14] ),
    .A1(net738),
    .S(net809),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _14470_ (.A0(\core.registers[18][15] ),
    .A1(net742),
    .S(net810),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _14471_ (.A0(\core.registers[18][16] ),
    .A1(net830),
    .S(net810),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _14472_ (.A0(\core.registers[18][17] ),
    .A1(net835),
    .S(net809),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _14473_ (.A0(\core.registers[18][18] ),
    .A1(net838),
    .S(net811),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _14474_ (.A0(\core.registers[18][19] ),
    .A1(net842),
    .S(net809),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _14475_ (.A0(\core.registers[18][20] ),
    .A1(net848),
    .S(net809),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _14476_ (.A0(\core.registers[18][21] ),
    .A1(net852),
    .S(net809),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _14477_ (.A0(\core.registers[18][22] ),
    .A1(net858),
    .S(net810),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _14478_ (.A0(\core.registers[18][23] ),
    .A1(net862),
    .S(net809),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _14479_ (.A0(\core.registers[18][24] ),
    .A1(net994),
    .S(net809),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _14480_ (.A0(\core.registers[18][25] ),
    .A1(net998),
    .S(net809),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _14481_ (.A0(\core.registers[18][26] ),
    .A1(net1002),
    .S(net811),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _14482_ (.A0(\core.registers[18][27] ),
    .A1(net867),
    .S(net811),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _14483_ (.A0(\core.registers[18][28] ),
    .A1(net871),
    .S(net812),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _14484_ (.A0(\core.registers[18][29] ),
    .A1(net874),
    .S(net811),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _14485_ (.A0(\core.registers[18][30] ),
    .A1(net878),
    .S(net811),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _14486_ (.A0(\core.registers[18][31] ),
    .A1(net1023),
    .S(net809),
    .X(_00580_));
 sky130_fd_sc_hd__nor2_1 _14487_ (.A(net1906),
    .B(net375),
    .Y(_00581_));
 sky130_fd_sc_hd__and3_4 _14488_ (.A(net1801),
    .B(_03905_),
    .C(_03906_),
    .X(_08770_));
 sky130_fd_sc_hd__nand2_2 _14489_ (.A(_08677_),
    .B(_08770_),
    .Y(_08771_));
 sky130_fd_sc_hd__mux2_1 _14490_ (.A0(net1076),
    .A1(\core.registers[13][0] ),
    .S(net960),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _14491_ (.A0(net1082),
    .A1(\core.registers[13][1] ),
    .S(net958),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _14492_ (.A0(net1086),
    .A1(\core.registers[13][2] ),
    .S(net960),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _14493_ (.A0(net1089),
    .A1(\core.registers[13][3] ),
    .S(net957),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _14494_ (.A0(net1027),
    .A1(\core.registers[13][4] ),
    .S(net959),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _14495_ (.A0(net1031),
    .A1(\core.registers[13][5] ),
    .S(net959),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _14496_ (.A0(net1037),
    .A1(\core.registers[13][6] ),
    .S(net959),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _14497_ (.A0(net1137),
    .A1(\core.registers[13][7] ),
    .S(net959),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _14498_ (.A0(net896),
    .A1(\core.registers[13][8] ),
    .S(net959),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _14499_ (.A0(net900),
    .A1(\core.registers[13][9] ),
    .S(net958),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _14500_ (.A0(net760),
    .A1(\core.registers[13][10] ),
    .S(net958),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _14501_ (.A0(net761),
    .A1(\core.registers[13][11] ),
    .S(net958),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _14502_ (.A0(net728),
    .A1(\core.registers[13][12] ),
    .S(net958),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _14503_ (.A0(net732),
    .A1(\core.registers[13][13] ),
    .S(net958),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _14504_ (.A0(net736),
    .A1(\core.registers[13][14] ),
    .S(net957),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _14505_ (.A0(net740),
    .A1(\core.registers[13][15] ),
    .S(net960),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _14506_ (.A0(net831),
    .A1(\core.registers[13][16] ),
    .S(net959),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _14507_ (.A0(net834),
    .A1(\core.registers[13][17] ),
    .S(net957),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _14508_ (.A0(net840),
    .A1(\core.registers[13][18] ),
    .S(net958),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _14509_ (.A0(net843),
    .A1(\core.registers[13][19] ),
    .S(net957),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _14510_ (.A0(net849),
    .A1(\core.registers[13][20] ),
    .S(net957),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _14511_ (.A0(net850),
    .A1(\core.registers[13][21] ),
    .S(net957),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _14512_ (.A0(net855),
    .A1(\core.registers[13][22] ),
    .S(net959),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _14513_ (.A0(net860),
    .A1(\core.registers[13][23] ),
    .S(net957),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _14514_ (.A0(net992),
    .A1(\core.registers[13][24] ),
    .S(net957),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _14515_ (.A0(net996),
    .A1(\core.registers[13][25] ),
    .S(net957),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _14516_ (.A0(net1001),
    .A1(\core.registers[13][26] ),
    .S(net957),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _14517_ (.A0(net864),
    .A1(\core.registers[13][27] ),
    .S(net959),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _14518_ (.A0(net869),
    .A1(\core.registers[13][28] ),
    .S(net958),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _14519_ (.A0(net876),
    .A1(\core.registers[13][29] ),
    .S(net958),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _14520_ (.A0(net878),
    .A1(\core.registers[13][30] ),
    .S(net958),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _14521_ (.A0(net1025),
    .A1(\core.registers[13][31] ),
    .S(net960),
    .X(_00613_));
 sky130_fd_sc_hd__a21oi_1 _14522_ (.A1(net601),
    .A2(net1311),
    .B1(net525),
    .Y(_08772_));
 sky130_fd_sc_hd__o21ba_1 _14523_ (.A1(\coreWBInterface.state[1] ),
    .A2(_08772_),
    .B1_N(net370),
    .X(_08773_));
 sky130_fd_sc_hd__a21o_1 _14524_ (.A1(net42),
    .A2(net333),
    .B1(net1872),
    .X(_08774_));
 sky130_fd_sc_hd__nor3_1 _14525_ (.A(_06677_),
    .B(_08773_),
    .C(net1295),
    .Y(_00614_));
 sky130_fd_sc_hd__nor2_1 _14526_ (.A(net9),
    .B(_06676_),
    .Y(_08775_));
 sky130_fd_sc_hd__nor2_1 _14527_ (.A(\coreWBInterface.state[0] ),
    .B(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__or2_1 _14528_ (.A(_03852_),
    .B(_06676_),
    .X(_08777_));
 sky130_fd_sc_hd__o22a_1 _14529_ (.A1(\coreWBInterface.readDataBuffered[0] ),
    .A2(net1270),
    .B1(net1293),
    .B2(net10),
    .X(_08778_));
 sky130_fd_sc_hd__or2_1 _14530_ (.A(net1297),
    .B(_08778_),
    .X(_00615_));
 sky130_fd_sc_hd__o22a_1 _14531_ (.A1(\coreWBInterface.readDataBuffered[1] ),
    .A2(net1268),
    .B1(net1291),
    .B2(net21),
    .X(_08779_));
 sky130_fd_sc_hd__or2_1 _14532_ (.A(net1295),
    .B(_08779_),
    .X(_00616_));
 sky130_fd_sc_hd__o22a_1 _14533_ (.A1(\coreWBInterface.readDataBuffered[2] ),
    .A2(net1268),
    .B1(net1291),
    .B2(net32),
    .X(_08780_));
 sky130_fd_sc_hd__or2_1 _14534_ (.A(net1295),
    .B(_08780_),
    .X(_00617_));
 sky130_fd_sc_hd__o22a_1 _14535_ (.A1(\coreWBInterface.readDataBuffered[3] ),
    .A2(net1268),
    .B1(net1291),
    .B2(net35),
    .X(_08781_));
 sky130_fd_sc_hd__or2_1 _14536_ (.A(net1295),
    .B(_08781_),
    .X(_00618_));
 sky130_fd_sc_hd__o22a_1 _14537_ (.A1(\coreWBInterface.readDataBuffered[4] ),
    .A2(net1268),
    .B1(net1291),
    .B2(net36),
    .X(_08782_));
 sky130_fd_sc_hd__or2_1 _14538_ (.A(net1295),
    .B(_08782_),
    .X(_00619_));
 sky130_fd_sc_hd__o22a_1 _14539_ (.A1(\coreWBInterface.readDataBuffered[5] ),
    .A2(net1268),
    .B1(net1291),
    .B2(net37),
    .X(_08783_));
 sky130_fd_sc_hd__or2_1 _14540_ (.A(net1295),
    .B(_08783_),
    .X(_00620_));
 sky130_fd_sc_hd__o22a_1 _14541_ (.A1(\coreWBInterface.readDataBuffered[6] ),
    .A2(net1268),
    .B1(net1291),
    .B2(net38),
    .X(_08784_));
 sky130_fd_sc_hd__or2_1 _14542_ (.A(net1295),
    .B(_08784_),
    .X(_00621_));
 sky130_fd_sc_hd__o22a_1 _14543_ (.A1(\coreWBInterface.readDataBuffered[7] ),
    .A2(net1268),
    .B1(net1291),
    .B2(net39),
    .X(_08785_));
 sky130_fd_sc_hd__or2_1 _14544_ (.A(net1295),
    .B(_08785_),
    .X(_00622_));
 sky130_fd_sc_hd__o22a_1 _14545_ (.A1(\coreWBInterface.readDataBuffered[8] ),
    .A2(net1269),
    .B1(net1292),
    .B2(net40),
    .X(_08786_));
 sky130_fd_sc_hd__or2_1 _14546_ (.A(net1296),
    .B(_08786_),
    .X(_00623_));
 sky130_fd_sc_hd__o22a_1 _14547_ (.A1(\coreWBInterface.readDataBuffered[9] ),
    .A2(net1270),
    .B1(net1293),
    .B2(net41),
    .X(_08787_));
 sky130_fd_sc_hd__or2_1 _14548_ (.A(net1297),
    .B(_08787_),
    .X(_00624_));
 sky130_fd_sc_hd__o22a_1 _14549_ (.A1(\coreWBInterface.readDataBuffered[10] ),
    .A2(net1270),
    .B1(net1293),
    .B2(net11),
    .X(_08788_));
 sky130_fd_sc_hd__or2_1 _14550_ (.A(net1297),
    .B(_08788_),
    .X(_00625_));
 sky130_fd_sc_hd__o22a_1 _14551_ (.A1(\coreWBInterface.readDataBuffered[11] ),
    .A2(net1270),
    .B1(net1293),
    .B2(net12),
    .X(_08789_));
 sky130_fd_sc_hd__or2_1 _14552_ (.A(net1297),
    .B(_08789_),
    .X(_00626_));
 sky130_fd_sc_hd__o22a_1 _14553_ (.A1(\coreWBInterface.readDataBuffered[12] ),
    .A2(net1268),
    .B1(net1291),
    .B2(net13),
    .X(_08790_));
 sky130_fd_sc_hd__or2_1 _14554_ (.A(net1298),
    .B(_08790_),
    .X(_00627_));
 sky130_fd_sc_hd__o22a_1 _14555_ (.A1(\coreWBInterface.readDataBuffered[13] ),
    .A2(net1268),
    .B1(net1291),
    .B2(net14),
    .X(_08791_));
 sky130_fd_sc_hd__or2_1 _14556_ (.A(net1298),
    .B(_08791_),
    .X(_00628_));
 sky130_fd_sc_hd__o22a_1 _14557_ (.A1(\coreWBInterface.readDataBuffered[14] ),
    .A2(net1269),
    .B1(net1292),
    .B2(net15),
    .X(_08792_));
 sky130_fd_sc_hd__or2_1 _14558_ (.A(net1296),
    .B(_08792_),
    .X(_00629_));
 sky130_fd_sc_hd__o22a_1 _14559_ (.A1(\coreWBInterface.readDataBuffered[15] ),
    .A2(net1268),
    .B1(net1291),
    .B2(net16),
    .X(_08793_));
 sky130_fd_sc_hd__or2_1 _14560_ (.A(net1298),
    .B(_08793_),
    .X(_00630_));
 sky130_fd_sc_hd__o22a_1 _14561_ (.A1(\coreWBInterface.readDataBuffered[16] ),
    .A2(net1271),
    .B1(net1294),
    .B2(net17),
    .X(_08794_));
 sky130_fd_sc_hd__or2_1 _14562_ (.A(net1298),
    .B(_08794_),
    .X(_00631_));
 sky130_fd_sc_hd__o22a_1 _14563_ (.A1(\coreWBInterface.readDataBuffered[17] ),
    .A2(net1269),
    .B1(net1292),
    .B2(net18),
    .X(_08795_));
 sky130_fd_sc_hd__or2_1 _14564_ (.A(net1296),
    .B(_08795_),
    .X(_00632_));
 sky130_fd_sc_hd__o22a_1 _14565_ (.A1(\coreWBInterface.readDataBuffered[18] ),
    .A2(net1270),
    .B1(net1293),
    .B2(net19),
    .X(_08796_));
 sky130_fd_sc_hd__or2_1 _14566_ (.A(net1297),
    .B(_08796_),
    .X(_00633_));
 sky130_fd_sc_hd__o22a_1 _14567_ (.A1(\coreWBInterface.readDataBuffered[19] ),
    .A2(net1270),
    .B1(net1293),
    .B2(net20),
    .X(_08797_));
 sky130_fd_sc_hd__or2_1 _14568_ (.A(net1297),
    .B(_08797_),
    .X(_00634_));
 sky130_fd_sc_hd__o22a_1 _14569_ (.A1(\coreWBInterface.readDataBuffered[20] ),
    .A2(net1270),
    .B1(net1293),
    .B2(net22),
    .X(_08798_));
 sky130_fd_sc_hd__or2_1 _14570_ (.A(net1297),
    .B(_08798_),
    .X(_00635_));
 sky130_fd_sc_hd__o22a_1 _14571_ (.A1(\coreWBInterface.readDataBuffered[21] ),
    .A2(net1270),
    .B1(net1293),
    .B2(net23),
    .X(_08799_));
 sky130_fd_sc_hd__or2_1 _14572_ (.A(net1297),
    .B(_08799_),
    .X(_00636_));
 sky130_fd_sc_hd__o22a_1 _14573_ (.A1(\coreWBInterface.readDataBuffered[22] ),
    .A2(net1270),
    .B1(net1293),
    .B2(net24),
    .X(_08800_));
 sky130_fd_sc_hd__or2_1 _14574_ (.A(net1297),
    .B(_08800_),
    .X(_00637_));
 sky130_fd_sc_hd__o22a_1 _14575_ (.A1(\coreWBInterface.readDataBuffered[23] ),
    .A2(net1270),
    .B1(net1293),
    .B2(net25),
    .X(_08801_));
 sky130_fd_sc_hd__or2_1 _14576_ (.A(net1297),
    .B(_08801_),
    .X(_00638_));
 sky130_fd_sc_hd__o22a_1 _14577_ (.A1(\coreWBInterface.readDataBuffered[24] ),
    .A2(net1269),
    .B1(net1292),
    .B2(net26),
    .X(_08802_));
 sky130_fd_sc_hd__or2_1 _14578_ (.A(net1296),
    .B(_08802_),
    .X(_00639_));
 sky130_fd_sc_hd__o22a_1 _14579_ (.A1(\coreWBInterface.readDataBuffered[25] ),
    .A2(net1269),
    .B1(net1292),
    .B2(net27),
    .X(_08803_));
 sky130_fd_sc_hd__or2_1 _14580_ (.A(net1296),
    .B(_08803_),
    .X(_00640_));
 sky130_fd_sc_hd__o22a_1 _14581_ (.A1(\coreWBInterface.readDataBuffered[26] ),
    .A2(net1269),
    .B1(net1292),
    .B2(net28),
    .X(_08804_));
 sky130_fd_sc_hd__or2_1 _14582_ (.A(net1296),
    .B(_08804_),
    .X(_00641_));
 sky130_fd_sc_hd__o22a_1 _14583_ (.A1(\coreWBInterface.readDataBuffered[27] ),
    .A2(net1269),
    .B1(net1292),
    .B2(net29),
    .X(_08805_));
 sky130_fd_sc_hd__or2_1 _14584_ (.A(net1296),
    .B(_08805_),
    .X(_00642_));
 sky130_fd_sc_hd__o22a_1 _14585_ (.A1(\coreWBInterface.readDataBuffered[28] ),
    .A2(net1269),
    .B1(net1292),
    .B2(net30),
    .X(_08806_));
 sky130_fd_sc_hd__or2_1 _14586_ (.A(net1298),
    .B(_08806_),
    .X(_00643_));
 sky130_fd_sc_hd__o22a_1 _14587_ (.A1(\coreWBInterface.readDataBuffered[29] ),
    .A2(net1269),
    .B1(net1292),
    .B2(net31),
    .X(_08807_));
 sky130_fd_sc_hd__or2_1 _14588_ (.A(net1296),
    .B(_08807_),
    .X(_00644_));
 sky130_fd_sc_hd__o22a_1 _14589_ (.A1(\coreWBInterface.readDataBuffered[30] ),
    .A2(net1269),
    .B1(net1292),
    .B2(net33),
    .X(_08808_));
 sky130_fd_sc_hd__or2_1 _14590_ (.A(net1296),
    .B(_08808_),
    .X(_00645_));
 sky130_fd_sc_hd__o22a_1 _14591_ (.A1(\coreWBInterface.readDataBuffered[31] ),
    .A2(net1271),
    .B1(net1294),
    .B2(net34),
    .X(_08809_));
 sky130_fd_sc_hd__or2_1 _14592_ (.A(net1296),
    .B(_08809_),
    .X(_00646_));
 sky130_fd_sc_hd__a21o_1 _14593_ (.A1(_04057_),
    .A2(net525),
    .B1(net333),
    .X(_08810_));
 sky130_fd_sc_hd__a2bb2o_1 _14594_ (.A1_N(_08772_),
    .A2_N(net333),
    .B1(net9),
    .B2(_06677_),
    .X(_08811_));
 sky130_fd_sc_hd__o2bb2a_1 _14595_ (.A1_N(_08810_),
    .A2_N(_08811_),
    .B1(net9),
    .B2(_03854_),
    .X(_08812_));
 sky130_fd_sc_hd__nor2_1 _14596_ (.A(net1295),
    .B(_08812_),
    .Y(_00647_));
 sky130_fd_sc_hd__o31a_1 _14597_ (.A1(net333),
    .A2(_04056_),
    .A3(_06711_),
    .B1(_08811_),
    .X(_08813_));
 sky130_fd_sc_hd__o21ba_1 _14598_ (.A1(_08775_),
    .A2(_08813_),
    .B1_N(net1295),
    .X(_00648_));
 sky130_fd_sc_hd__or2_4 _14599_ (.A(_06853_),
    .B(_08678_),
    .X(_08814_));
 sky130_fd_sc_hd__mux2_1 _14600_ (.A0(net1078),
    .A1(\core.registers[17][0] ),
    .S(net954),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _14601_ (.A0(net1082),
    .A1(\core.registers[17][1] ),
    .S(net955),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _14602_ (.A0(net1085),
    .A1(\core.registers[17][2] ),
    .S(net954),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _14603_ (.A0(net1090),
    .A1(\core.registers[17][3] ),
    .S(net953),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _14604_ (.A0(net1027),
    .A1(\core.registers[17][4] ),
    .S(net956),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _14605_ (.A0(net1033),
    .A1(\core.registers[17][5] ),
    .S(net956),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _14606_ (.A0(net1035),
    .A1(\core.registers[17][6] ),
    .S(net956),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _14607_ (.A0(net1139),
    .A1(\core.registers[17][7] ),
    .S(net956),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _14608_ (.A0(net898),
    .A1(\core.registers[17][8] ),
    .S(net955),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _14609_ (.A0(net902),
    .A1(\core.registers[17][9] ),
    .S(net955),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _14610_ (.A0(net759),
    .A1(\core.registers[17][10] ),
    .S(net955),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _14611_ (.A0(net762),
    .A1(\core.registers[17][11] ),
    .S(net955),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _14612_ (.A0(net729),
    .A1(\core.registers[17][12] ),
    .S(net956),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _14613_ (.A0(net733),
    .A1(\core.registers[17][13] ),
    .S(net955),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _14614_ (.A0(net738),
    .A1(\core.registers[17][14] ),
    .S(net953),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _14615_ (.A0(net741),
    .A1(\core.registers[17][15] ),
    .S(net954),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _14616_ (.A0(net830),
    .A1(\core.registers[17][16] ),
    .S(net954),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _14617_ (.A0(net835),
    .A1(\core.registers[17][17] ),
    .S(net953),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _14618_ (.A0(net838),
    .A1(\core.registers[17][18] ),
    .S(net955),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _14619_ (.A0(net844),
    .A1(\core.registers[17][19] ),
    .S(net953),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _14620_ (.A0(net847),
    .A1(\core.registers[17][20] ),
    .S(net953),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _14621_ (.A0(net852),
    .A1(\core.registers[17][21] ),
    .S(net953),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _14622_ (.A0(net857),
    .A1(\core.registers[17][22] ),
    .S(net954),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _14623_ (.A0(net862),
    .A1(\core.registers[17][23] ),
    .S(net953),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _14624_ (.A0(net994),
    .A1(\core.registers[17][24] ),
    .S(net953),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _14625_ (.A0(net998),
    .A1(\core.registers[17][25] ),
    .S(net953),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _14626_ (.A0(net1003),
    .A1(\core.registers[17][26] ),
    .S(net956),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _14627_ (.A0(net867),
    .A1(\core.registers[17][27] ),
    .S(net955),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _14628_ (.A0(net871),
    .A1(\core.registers[17][28] ),
    .S(net956),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _14629_ (.A0(net874),
    .A1(\core.registers[17][29] ),
    .S(net955),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _14630_ (.A0(net879),
    .A1(\core.registers[17][30] ),
    .S(net955),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _14631_ (.A0(net1023),
    .A1(\core.registers[17][31] ),
    .S(net953),
    .X(_00680_));
 sky130_fd_sc_hd__nand2_2 _14632_ (.A(_08680_),
    .B(_08770_),
    .Y(_01893_));
 sky130_fd_sc_hd__mux2_1 _14633_ (.A0(net1076),
    .A1(\core.registers[12][0] ),
    .S(net952),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _14634_ (.A0(net1082),
    .A1(\core.registers[12][1] ),
    .S(net950),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _14635_ (.A0(net1086),
    .A1(\core.registers[12][2] ),
    .S(net952),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _14636_ (.A0(net1089),
    .A1(\core.registers[12][3] ),
    .S(net952),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _14637_ (.A0(net1027),
    .A1(\core.registers[12][4] ),
    .S(net951),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _14638_ (.A0(net1031),
    .A1(\core.registers[12][5] ),
    .S(net951),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _14639_ (.A0(net1037),
    .A1(\core.registers[12][6] ),
    .S(net951),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _14640_ (.A0(net1137),
    .A1(\core.registers[12][7] ),
    .S(net951),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _14641_ (.A0(net896),
    .A1(\core.registers[12][8] ),
    .S(net951),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _14642_ (.A0(net900),
    .A1(\core.registers[12][9] ),
    .S(net950),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _14643_ (.A0(net760),
    .A1(\core.registers[12][10] ),
    .S(net950),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _14644_ (.A0(net763),
    .A1(\core.registers[12][11] ),
    .S(net950),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _14645_ (.A0(net728),
    .A1(\core.registers[12][12] ),
    .S(net950),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _14646_ (.A0(net732),
    .A1(\core.registers[12][13] ),
    .S(net950),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _14647_ (.A0(net736),
    .A1(\core.registers[12][14] ),
    .S(net949),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _14648_ (.A0(net740),
    .A1(\core.registers[12][15] ),
    .S(net952),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _14649_ (.A0(net831),
    .A1(\core.registers[12][16] ),
    .S(net951),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _14650_ (.A0(net834),
    .A1(\core.registers[12][17] ),
    .S(net949),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _14651_ (.A0(net840),
    .A1(\core.registers[12][18] ),
    .S(net950),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(net844),
    .A1(\core.registers[12][19] ),
    .S(net949),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _14653_ (.A0(net847),
    .A1(\core.registers[12][20] ),
    .S(net949),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _14654_ (.A0(net850),
    .A1(\core.registers[12][21] ),
    .S(net949),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _14655_ (.A0(net855),
    .A1(\core.registers[12][22] ),
    .S(net951),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _14656_ (.A0(net861),
    .A1(\core.registers[12][23] ),
    .S(net949),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _14657_ (.A0(net992),
    .A1(\core.registers[12][24] ),
    .S(net949),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _14658_ (.A0(net996),
    .A1(\core.registers[12][25] ),
    .S(net949),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _14659_ (.A0(net1001),
    .A1(\core.registers[12][26] ),
    .S(net949),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _14660_ (.A0(net864),
    .A1(\core.registers[12][27] ),
    .S(net951),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _14661_ (.A0(net869),
    .A1(\core.registers[12][28] ),
    .S(net950),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _14662_ (.A0(net876),
    .A1(\core.registers[12][29] ),
    .S(net950),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _14663_ (.A0(net878),
    .A1(\core.registers[12][30] ),
    .S(net950),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _14664_ (.A0(net1025),
    .A1(\core.registers[12][31] ),
    .S(net949),
    .X(_00712_));
 sky130_fd_sc_hd__a21bo_1 _14665_ (.A1(_07005_),
    .A2(net1273),
    .B1_N(_06704_),
    .X(_01894_));
 sky130_fd_sc_hd__a21o_2 _14666_ (.A1(net505),
    .A2(_06701_),
    .B1(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__a211o_4 _14667_ (.A1(net505),
    .A2(_06701_),
    .B1(_06702_),
    .C1(_01894_),
    .X(_01896_));
 sky130_fd_sc_hd__nor2_1 _14668_ (.A(_07020_),
    .B(_07158_),
    .Y(_01897_));
 sky130_fd_sc_hd__or2_2 _14669_ (.A(_07020_),
    .B(_07158_),
    .X(_01898_));
 sky130_fd_sc_hd__nor2_2 _14670_ (.A(_07031_),
    .B(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__or2_2 _14671_ (.A(_07031_),
    .B(_01898_),
    .X(_01900_));
 sky130_fd_sc_hd__and4bb_1 _14672_ (.A_N(_07027_),
    .B_N(_07028_),
    .C(_07029_),
    .D(_01897_),
    .X(_01901_));
 sky130_fd_sc_hd__or4b_1 _14673_ (.A(_07027_),
    .B(_07028_),
    .C(_01898_),
    .D_N(_07029_),
    .X(_01902_));
 sky130_fd_sc_hd__or2_1 _14674_ (.A(\core.csr.currentInstruction[0] ),
    .B(net937),
    .X(_01903_));
 sky130_fd_sc_hd__or3_4 _14675_ (.A(_07030_),
    .B(_07032_),
    .C(_07033_),
    .X(_01904_));
 sky130_fd_sc_hd__inv_2 _14676_ (.A(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__and4_2 _14677_ (.A(_07021_),
    .B(_07026_),
    .C(_01897_),
    .D(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__a221o_1 _14678_ (.A1(net1020),
    .A2(_07252_),
    .B1(_01906_),
    .B2(\core.registers[0][0] ),
    .C1(net941),
    .X(_01907_));
 sky130_fd_sc_hd__and4_1 _14679_ (.A(_07021_),
    .B(_07026_),
    .C(_01897_),
    .D(_01905_),
    .X(_01908_));
 sky130_fd_sc_hd__or4b_4 _14680_ (.A(_07027_),
    .B(_07028_),
    .C(_01898_),
    .D_N(_07029_),
    .X(_01909_));
 sky130_fd_sc_hd__and3b_1 _14681_ (.A_N(_07025_),
    .B(_01897_),
    .C(_07021_),
    .X(_01910_));
 sky130_fd_sc_hd__nor2_2 _14682_ (.A(_07024_),
    .B(_01904_),
    .Y(_01911_));
 sky130_fd_sc_hd__and2_2 _14683_ (.A(_01910_),
    .B(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__a21o_1 _14684_ (.A1(_01903_),
    .A2(_01907_),
    .B1(net945),
    .X(_01913_));
 sky130_fd_sc_hd__and2_1 _14685_ (.A(\wbSRAMInterface.currentByteSelect[0] ),
    .B(net1230),
    .X(_01914_));
 sky130_fd_sc_hd__nand2_4 _14686_ (.A(\wbSRAMInterface.currentByteSelect[0] ),
    .B(net1230),
    .Y(_01915_));
 sky130_fd_sc_hd__or2_1 _14687_ (.A(_07039_),
    .B(_07040_),
    .X(_01916_));
 sky130_fd_sc_hd__or4_4 _14688_ (.A(_07020_),
    .B(_07027_),
    .C(_01904_),
    .D(_01916_),
    .X(_01917_));
 sky130_fd_sc_hd__a21oi_1 _14689_ (.A1(_06703_),
    .A2(net1232),
    .B1(_07010_),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2_4 _14690_ (.A(_07041_),
    .B(_01915_),
    .Y(_01919_));
 sky130_fd_sc_hd__o211a_1 _14691_ (.A1(net450),
    .A2(net942),
    .B1(_01913_),
    .C1(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__o21ba_1 _14692_ (.A1(_07010_),
    .A2(net1232),
    .B1_N(_01917_),
    .X(_01921_));
 sky130_fd_sc_hd__o21ai_1 _14693_ (.A1(_06703_),
    .A2(_07010_),
    .B1(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__a21o_1 _14694_ (.A1(_07041_),
    .A2(_01922_),
    .B1(_07006_),
    .X(_01923_));
 sky130_fd_sc_hd__a211o_1 _14695_ (.A1(net1726),
    .A2(_01914_),
    .B1(_01920_),
    .C1(net673),
    .X(_01924_));
 sky130_fd_sc_hd__nand2_8 _14696_ (.A(net1738),
    .B(\localMemoryInterface.lastWBByteSelect[0] ),
    .Y(_01925_));
 sky130_fd_sc_hd__mux2_8 _14697_ (.A0(net43),
    .A1(net68),
    .S(net1741),
    .X(_01926_));
 sky130_fd_sc_hd__nor2_1 _14698_ (.A(_01925_),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__o2bb2a_2 _14699_ (.A1_N(net1277),
    .A2_N(_01924_),
    .B1(_01927_),
    .B2(net1908),
    .X(_01928_));
 sky130_fd_sc_hd__nor2_1 _14700_ (.A(net491),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__a211o_1 _14701_ (.A1(net410),
    .A2(net491),
    .B1(_01929_),
    .C1(net1880),
    .X(_00713_));
 sky130_fd_sc_hd__a2bb2o_1 _14702_ (.A1_N(_07161_),
    .A2_N(_07484_),
    .B1(_01912_),
    .B2(\core.registers[0][1] ),
    .X(_01930_));
 sky130_fd_sc_hd__mux2_1 _14703_ (.A0(\core.csr.currentInstruction[1] ),
    .A1(_01930_),
    .S(_01909_),
    .X(_01931_));
 sky130_fd_sc_hd__or2_1 _14704_ (.A(net461),
    .B(net943),
    .X(_01932_));
 sky130_fd_sc_hd__o211a_1 _14705_ (.A1(net947),
    .A2(_01931_),
    .B1(_01932_),
    .C1(_01919_),
    .X(_01933_));
 sky130_fd_sc_hd__a311o_1 _14706_ (.A1(\coreManagement.control[1] ),
    .A2(_07041_),
    .A3(_01914_),
    .B1(net673),
    .C1(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__mux2_8 _14707_ (.A0(net54),
    .A1(net69),
    .S(net1741),
    .X(_01935_));
 sky130_fd_sc_hd__nor2_1 _14708_ (.A(_01925_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__o2bb2a_2 _14709_ (.A1_N(net1277),
    .A2_N(_01934_),
    .B1(_01936_),
    .B2(net1908),
    .X(_01937_));
 sky130_fd_sc_hd__nor2_1 _14710_ (.A(net491),
    .B(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__a211o_1 _14711_ (.A1(net421),
    .A2(net491),
    .B1(_01938_),
    .C1(net1881),
    .X(_00714_));
 sky130_fd_sc_hd__a32o_1 _14712_ (.A1(\core.registers[0][2] ),
    .A2(_01910_),
    .A3(_01911_),
    .B1(net1020),
    .B2(_07565_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _14713_ (.A0(\core.csr.currentInstruction[2] ),
    .A1(_01939_),
    .S(_01909_),
    .X(_01940_));
 sky130_fd_sc_hd__nand2_1 _14714_ (.A(_03827_),
    .B(net945),
    .Y(_01941_));
 sky130_fd_sc_hd__o211a_1 _14715_ (.A1(net947),
    .A2(_01940_),
    .B1(_01941_),
    .C1(_01919_),
    .X(_01942_));
 sky130_fd_sc_hd__a311o_1 _14716_ (.A1(\core.management_interruptEnable ),
    .A2(_07041_),
    .A3(_01914_),
    .B1(net673),
    .C1(_01942_),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_8 _14717_ (.A0(net65),
    .A1(net70),
    .S(net1741),
    .X(_01944_));
 sky130_fd_sc_hd__nor2_1 _14718_ (.A(_01925_),
    .B(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__o2bb2a_2 _14719_ (.A1_N(net1277),
    .A2_N(_01943_),
    .B1(_01945_),
    .B2(net1908),
    .X(_01946_));
 sky130_fd_sc_hd__nor2_1 _14720_ (.A(net491),
    .B(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__a211o_1 _14721_ (.A1(net432),
    .A2(net491),
    .B1(_01947_),
    .C1(net1881),
    .X(_00715_));
 sky130_fd_sc_hd__a32o_1 _14722_ (.A1(\core.registers[0][3] ),
    .A2(_01910_),
    .A3(_01911_),
    .B1(net1020),
    .B2(_07621_),
    .X(_01948_));
 sky130_fd_sc_hd__mux2_1 _14723_ (.A0(\core.csr.currentInstruction[3] ),
    .A1(_01948_),
    .S(_01909_),
    .X(_01949_));
 sky130_fd_sc_hd__or2_1 _14724_ (.A(net475),
    .B(net942),
    .X(_01950_));
 sky130_fd_sc_hd__o211a_1 _14725_ (.A1(net946),
    .A2(_01949_),
    .B1(_01950_),
    .C1(_01919_),
    .X(_01951_));
 sky130_fd_sc_hd__o21ba_1 _14726_ (.A1(_01917_),
    .A2(_01918_),
    .B1_N(_07044_),
    .X(_01952_));
 sky130_fd_sc_hd__o21ai_2 _14727_ (.A1(net672),
    .A2(_01951_),
    .B1(net1277),
    .Y(_01953_));
 sky130_fd_sc_hd__mux2_8 _14728_ (.A0(net76),
    .A1(net71),
    .S(net1741),
    .X(_01954_));
 sky130_fd_sc_hd__o21bai_4 _14729_ (.A1(_01925_),
    .A2(_01954_),
    .B1_N(net1909),
    .Y(_01955_));
 sky130_fd_sc_hd__a21oi_4 _14730_ (.A1(_01953_),
    .A2(_01955_),
    .B1(net489),
    .Y(_01956_));
 sky130_fd_sc_hd__a211o_1 _14731_ (.A1(net435),
    .A2(net491),
    .B1(_01956_),
    .C1(net1880),
    .X(_00716_));
 sky130_fd_sc_hd__or2_1 _14732_ (.A(\core.csr.currentInstruction[4] ),
    .B(net938),
    .X(_01957_));
 sky130_fd_sc_hd__a221o_1 _14733_ (.A1(net1021),
    .A2(_07676_),
    .B1(net934),
    .B2(\core.registers[0][4] ),
    .C1(net940),
    .X(_01958_));
 sky130_fd_sc_hd__a21o_1 _14734_ (.A1(_01957_),
    .A2(_01958_),
    .B1(net948),
    .X(_01959_));
 sky130_fd_sc_hd__o211a_1 _14735_ (.A1(net1748),
    .A2(net942),
    .B1(_01919_),
    .C1(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__o21ai_2 _14736_ (.A1(net672),
    .A2(_01960_),
    .B1(net1276),
    .Y(_01961_));
 sky130_fd_sc_hd__mux2_8 _14737_ (.A0(net87),
    .A1(net72),
    .S(net1741),
    .X(_01962_));
 sky130_fd_sc_hd__o21bai_4 _14738_ (.A1(_01925_),
    .A2(_01962_),
    .B1_N(net1909),
    .Y(_01963_));
 sky130_fd_sc_hd__a21oi_4 _14739_ (.A1(_01961_),
    .A2(_01963_),
    .B1(net488),
    .Y(_01964_));
 sky130_fd_sc_hd__a211o_1 _14740_ (.A1(net436),
    .A2(net492),
    .B1(_01964_),
    .C1(net1881),
    .X(_00717_));
 sky130_fd_sc_hd__nand2_1 _14741_ (.A(_03847_),
    .B(net940),
    .Y(_01965_));
 sky130_fd_sc_hd__a221o_1 _14742_ (.A1(net1021),
    .A2(_07721_),
    .B1(net934),
    .B2(\core.registers[0][5] ),
    .C1(net940),
    .X(_01966_));
 sky130_fd_sc_hd__a21o_1 _14743_ (.A1(_01965_),
    .A2(_01966_),
    .B1(net947),
    .X(_01967_));
 sky130_fd_sc_hd__o211a_1 _14744_ (.A1(net477),
    .A2(net942),
    .B1(_01919_),
    .C1(_01967_),
    .X(_01968_));
 sky130_fd_sc_hd__o21ai_2 _14745_ (.A1(net672),
    .A2(_01968_),
    .B1(net1276),
    .Y(_01969_));
 sky130_fd_sc_hd__mux2_8 _14746_ (.A0(net98),
    .A1(net73),
    .S(net1741),
    .X(_01970_));
 sky130_fd_sc_hd__o21bai_4 _14747_ (.A1(_01925_),
    .A2(_01970_),
    .B1_N(net1909),
    .Y(_01971_));
 sky130_fd_sc_hd__a21oi_4 _14748_ (.A1(_01969_),
    .A2(_01971_),
    .B1(net488),
    .Y(_01972_));
 sky130_fd_sc_hd__a211o_1 _14749_ (.A1(net437),
    .A2(net491),
    .B1(_01972_),
    .C1(net1882),
    .X(_00718_));
 sky130_fd_sc_hd__or2_1 _14750_ (.A(\core.csr.currentInstruction[6] ),
    .B(net938),
    .X(_01973_));
 sky130_fd_sc_hd__a221o_1 _14751_ (.A1(net1020),
    .A2(_07772_),
    .B1(net934),
    .B2(\core.registers[0][6] ),
    .C1(net940),
    .X(_01974_));
 sky130_fd_sc_hd__a21o_1 _14752_ (.A1(_01973_),
    .A2(_01974_),
    .B1(net947),
    .X(_01975_));
 sky130_fd_sc_hd__o211a_1 _14753_ (.A1(net478),
    .A2(net942),
    .B1(_01919_),
    .C1(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__o21ai_2 _14754_ (.A1(net672),
    .A2(_01976_),
    .B1(net1276),
    .Y(_01977_));
 sky130_fd_sc_hd__mux2_8 _14755_ (.A0(net103),
    .A1(net74),
    .S(net1741),
    .X(_01978_));
 sky130_fd_sc_hd__o21bai_4 _14756_ (.A1(_01925_),
    .A2(_01978_),
    .B1_N(net1909),
    .Y(_01979_));
 sky130_fd_sc_hd__a21oi_4 _14757_ (.A1(_01977_),
    .A2(_01979_),
    .B1(net488),
    .Y(_01980_));
 sky130_fd_sc_hd__a211o_1 _14758_ (.A1(net438),
    .A2(net491),
    .B1(_01980_),
    .C1(net1883),
    .X(_00719_));
 sky130_fd_sc_hd__or2_1 _14759_ (.A(\core.csr.currentInstruction[7] ),
    .B(net937),
    .X(_01981_));
 sky130_fd_sc_hd__a221o_2 _14760_ (.A1(net1021),
    .A2(_07813_),
    .B1(net934),
    .B2(\core.registers[0][7] ),
    .C1(net940),
    .X(_01982_));
 sky130_fd_sc_hd__a21o_1 _14761_ (.A1(_01981_),
    .A2(_01982_),
    .B1(net946),
    .X(_01983_));
 sky130_fd_sc_hd__o211a_1 _14762_ (.A1(net479),
    .A2(net942),
    .B1(_01919_),
    .C1(_01983_),
    .X(_01984_));
 sky130_fd_sc_hd__o21ai_2 _14763_ (.A1(net672),
    .A2(_01984_),
    .B1(net1276),
    .Y(_01985_));
 sky130_fd_sc_hd__mux2_8 _14764_ (.A0(net104),
    .A1(net75),
    .S(net1741),
    .X(_01986_));
 sky130_fd_sc_hd__o21bai_4 _14765_ (.A1(_01925_),
    .A2(_01986_),
    .B1_N(net1909),
    .Y(_01987_));
 sky130_fd_sc_hd__a21oi_4 _14766_ (.A1(_01985_),
    .A2(_01987_),
    .B1(net488),
    .Y(_01988_));
 sky130_fd_sc_hd__a211o_1 _14767_ (.A1(net439),
    .A2(net491),
    .B1(_01988_),
    .C1(net1883),
    .X(_00720_));
 sky130_fd_sc_hd__or2_1 _14768_ (.A(\core.csr.currentInstruction[8] ),
    .B(net937),
    .X(_01989_));
 sky130_fd_sc_hd__a221o_2 _14769_ (.A1(net1022),
    .A2(_07874_),
    .B1(net934),
    .B2(\core.registers[0][8] ),
    .C1(net940),
    .X(_01990_));
 sky130_fd_sc_hd__a21o_1 _14770_ (.A1(_01989_),
    .A2(_01990_),
    .B1(net946),
    .X(_01991_));
 sky130_fd_sc_hd__and4_4 _14771_ (.A(\wbSRAMInterface.currentByteSelect[1] ),
    .B(net1614),
    .C(net1230),
    .D(_07042_),
    .X(_01992_));
 sky130_fd_sc_hd__o211a_1 _14772_ (.A1(net480),
    .A2(net942),
    .B1(_01991_),
    .C1(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__o21ai_2 _14773_ (.A1(net672),
    .A2(_01993_),
    .B1(net1276),
    .Y(_01994_));
 sky130_fd_sc_hd__mux2_1 _14774_ (.A0(net105),
    .A1(net77),
    .S(net1741),
    .X(_01995_));
 sky130_fd_sc_hd__inv_2 _14775_ (.A(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__a31o_1 _14776_ (.A1(net1738),
    .A2(\localMemoryInterface.lastWBByteSelect[1] ),
    .A3(_01996_),
    .B1(net1909),
    .X(_01997_));
 sky130_fd_sc_hd__a21oi_4 _14777_ (.A1(_01994_),
    .A2(_01997_),
    .B1(net488),
    .Y(_01998_));
 sky130_fd_sc_hd__a211o_1 _14778_ (.A1(net440),
    .A2(net492),
    .B1(_01998_),
    .C1(net1883),
    .X(_00721_));
 sky130_fd_sc_hd__or2_1 _14779_ (.A(net1801),
    .B(net938),
    .X(_01999_));
 sky130_fd_sc_hd__a221o_1 _14780_ (.A1(net1021),
    .A2(_07910_),
    .B1(net934),
    .B2(\core.registers[0][9] ),
    .C1(net940),
    .X(_02000_));
 sky130_fd_sc_hd__a21o_1 _14781_ (.A1(_01999_),
    .A2(_02000_),
    .B1(net947),
    .X(_02001_));
 sky130_fd_sc_hd__o211a_1 _14782_ (.A1(net481),
    .A2(net944),
    .B1(_01992_),
    .C1(_02001_),
    .X(_02002_));
 sky130_fd_sc_hd__o21ai_2 _14783_ (.A1(net673),
    .A2(_02002_),
    .B1(net1276),
    .Y(_02003_));
 sky130_fd_sc_hd__mux2_1 _14784_ (.A0(net106),
    .A1(net78),
    .S(net1741),
    .X(_02004_));
 sky130_fd_sc_hd__inv_2 _14785_ (.A(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__a31o_1 _14786_ (.A1(net1738),
    .A2(\localMemoryInterface.lastWBByteSelect[1] ),
    .A3(_02005_),
    .B1(net1909),
    .X(_02006_));
 sky130_fd_sc_hd__a21oi_4 _14787_ (.A1(_02003_),
    .A2(_02006_),
    .B1(net488),
    .Y(_02007_));
 sky130_fd_sc_hd__a211o_1 _14788_ (.A1(net441),
    .A2(net492),
    .B1(_02007_),
    .C1(net1883),
    .X(_00722_));
 sky130_fd_sc_hd__or2_1 _14789_ (.A(\core.csr.currentInstruction[10] ),
    .B(net938),
    .X(_02008_));
 sky130_fd_sc_hd__a221o_1 _14790_ (.A1(net1021),
    .A2(_07943_),
    .B1(net934),
    .B2(\core.registers[0][10] ),
    .C1(net940),
    .X(_02009_));
 sky130_fd_sc_hd__a21o_1 _14791_ (.A1(_02008_),
    .A2(_02009_),
    .B1(net947),
    .X(_02010_));
 sky130_fd_sc_hd__o211a_1 _14792_ (.A1(net451),
    .A2(net944),
    .B1(_01992_),
    .C1(_02010_),
    .X(_02011_));
 sky130_fd_sc_hd__o21ai_2 _14793_ (.A1(net672),
    .A2(_02011_),
    .B1(net1276),
    .Y(_02012_));
 sky130_fd_sc_hd__mux2_1 _14794_ (.A0(net44),
    .A1(net79),
    .S(net1742),
    .X(_02013_));
 sky130_fd_sc_hd__inv_2 _14795_ (.A(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__a31o_1 _14796_ (.A1(net1738),
    .A2(\localMemoryInterface.lastWBByteSelect[1] ),
    .A3(_02014_),
    .B1(net1909),
    .X(_02015_));
 sky130_fd_sc_hd__a21oi_4 _14797_ (.A1(_02012_),
    .A2(_02015_),
    .B1(net489),
    .Y(_02016_));
 sky130_fd_sc_hd__a211o_1 _14798_ (.A1(net411),
    .A2(net492),
    .B1(_02016_),
    .C1(net1884),
    .X(_00723_));
 sky130_fd_sc_hd__a2bb2o_1 _14799_ (.A1_N(_07161_),
    .A2_N(_07977_),
    .B1(_01912_),
    .B2(\core.registers[0][11] ),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _14800_ (.A0(\core.csr.currentInstruction[11] ),
    .A1(_02017_),
    .S(_01909_),
    .X(_02018_));
 sky130_fd_sc_hd__or2_1 _14801_ (.A(net452),
    .B(net942),
    .X(_02019_));
 sky130_fd_sc_hd__o211a_1 _14802_ (.A1(net947),
    .A2(_02018_),
    .B1(_02019_),
    .C1(_01992_),
    .X(_02020_));
 sky130_fd_sc_hd__o21ai_2 _14803_ (.A1(net673),
    .A2(_02020_),
    .B1(net1277),
    .Y(_02021_));
 sky130_fd_sc_hd__mux2_1 _14804_ (.A0(net45),
    .A1(net80),
    .S(net1742),
    .X(_02022_));
 sky130_fd_sc_hd__inv_2 _14805_ (.A(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__a31o_1 _14806_ (.A1(net1738),
    .A2(\localMemoryInterface.lastWBByteSelect[1] ),
    .A3(_02023_),
    .B1(net1909),
    .X(_02024_));
 sky130_fd_sc_hd__a21oi_4 _14807_ (.A1(_02021_),
    .A2(_02024_),
    .B1(net489),
    .Y(_02025_));
 sky130_fd_sc_hd__a211o_1 _14808_ (.A1(net412),
    .A2(net494),
    .B1(_02025_),
    .C1(net1884),
    .X(_00724_));
 sky130_fd_sc_hd__a2bb2o_1 _14809_ (.A1_N(_07161_),
    .A2_N(_07997_),
    .B1(_01912_),
    .B2(\core.registers[0][12] ),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _14810_ (.A0(\core.csr.currentInstruction[12] ),
    .A1(_02026_),
    .S(_01909_),
    .X(_02027_));
 sky130_fd_sc_hd__or2_1 _14811_ (.A(net453),
    .B(net944),
    .X(_02028_));
 sky130_fd_sc_hd__o211a_1 _14812_ (.A1(net947),
    .A2(_02027_),
    .B1(_02028_),
    .C1(_01992_),
    .X(_02029_));
 sky130_fd_sc_hd__o21ai_2 _14813_ (.A1(net674),
    .A2(_02029_),
    .B1(net1277),
    .Y(_02030_));
 sky130_fd_sc_hd__mux2_2 _14814_ (.A0(net46),
    .A1(net81),
    .S(net1742),
    .X(_02031_));
 sky130_fd_sc_hd__clkinv_4 _14815_ (.A(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__a31o_2 _14816_ (.A1(net1738),
    .A2(\localMemoryInterface.lastWBByteSelect[1] ),
    .A3(_02032_),
    .B1(net1907),
    .X(_02033_));
 sky130_fd_sc_hd__a21oi_4 _14817_ (.A1(_02030_),
    .A2(_02033_),
    .B1(net489),
    .Y(_02034_));
 sky130_fd_sc_hd__a211o_1 _14818_ (.A1(net413),
    .A2(net494),
    .B1(_02034_),
    .C1(net1884),
    .X(_00725_));
 sky130_fd_sc_hd__a2bb2o_1 _14819_ (.A1_N(_07161_),
    .A2_N(_08034_),
    .B1(_01912_),
    .B2(\core.registers[0][13] ),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _14820_ (.A0(net1800),
    .A1(_02035_),
    .S(_01909_),
    .X(_02036_));
 sky130_fd_sc_hd__or2_1 _14821_ (.A(net454),
    .B(net944),
    .X(_02037_));
 sky130_fd_sc_hd__o211a_1 _14822_ (.A1(net948),
    .A2(_02036_),
    .B1(_02037_),
    .C1(_01992_),
    .X(_02038_));
 sky130_fd_sc_hd__o21ai_2 _14823_ (.A1(net674),
    .A2(_02038_),
    .B1(net1277),
    .Y(_02039_));
 sky130_fd_sc_hd__mux2_1 _14824_ (.A0(net47),
    .A1(net82),
    .S(net1742),
    .X(_02040_));
 sky130_fd_sc_hd__inv_2 _14825_ (.A(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__a31o_2 _14826_ (.A1(net1740),
    .A2(\localMemoryInterface.lastWBByteSelect[1] ),
    .A3(_02041_),
    .B1(net1907),
    .X(_02042_));
 sky130_fd_sc_hd__a21oi_4 _14827_ (.A1(_02039_),
    .A2(_02042_),
    .B1(net489),
    .Y(_02043_));
 sky130_fd_sc_hd__a211o_1 _14828_ (.A1(net414),
    .A2(net494),
    .B1(_02043_),
    .C1(net1884),
    .X(_00726_));
 sky130_fd_sc_hd__a2bb2o_1 _14829_ (.A1_N(_07161_),
    .A2_N(_08069_),
    .B1(_01912_),
    .B2(\core.registers[0][14] ),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _14830_ (.A0(net1799),
    .A1(_02044_),
    .S(_01909_),
    .X(_02045_));
 sky130_fd_sc_hd__or2_1 _14831_ (.A(net455),
    .B(net944),
    .X(_02046_));
 sky130_fd_sc_hd__o211a_1 _14832_ (.A1(net947),
    .A2(_02045_),
    .B1(_02046_),
    .C1(_01992_),
    .X(_02047_));
 sky130_fd_sc_hd__o21ai_2 _14833_ (.A1(net674),
    .A2(_02047_),
    .B1(net1277),
    .Y(_02048_));
 sky130_fd_sc_hd__mux2_1 _14834_ (.A0(net48),
    .A1(net83),
    .S(net1742),
    .X(_02049_));
 sky130_fd_sc_hd__inv_2 _14835_ (.A(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__a31o_2 _14836_ (.A1(net1740),
    .A2(\localMemoryInterface.lastWBByteSelect[1] ),
    .A3(_02050_),
    .B1(net1907),
    .X(_02051_));
 sky130_fd_sc_hd__a21oi_4 _14837_ (.A1(_02048_),
    .A2(_02051_),
    .B1(net489),
    .Y(_02052_));
 sky130_fd_sc_hd__a211o_1 _14838_ (.A1(net415),
    .A2(net494),
    .B1(_02052_),
    .C1(net1894),
    .X(_00727_));
 sky130_fd_sc_hd__or2_1 _14839_ (.A(\core.csr.currentInstruction[15] ),
    .B(net936),
    .X(_02053_));
 sky130_fd_sc_hd__a221o_1 _14840_ (.A1(net1019),
    .A2(_08123_),
    .B1(net933),
    .B2(\core.registers[0][15] ),
    .C1(net939),
    .X(_02054_));
 sky130_fd_sc_hd__a21o_1 _14841_ (.A1(_02053_),
    .A2(_02054_),
    .B1(net945),
    .X(_02055_));
 sky130_fd_sc_hd__o211a_1 _14842_ (.A1(net456),
    .A2(net944),
    .B1(_01992_),
    .C1(_02055_),
    .X(_02056_));
 sky130_fd_sc_hd__o21ai_2 _14843_ (.A1(net672),
    .A2(_02056_),
    .B1(net1276),
    .Y(_02057_));
 sky130_fd_sc_hd__mux2_2 _14844_ (.A0(net49),
    .A1(net84),
    .S(net1742),
    .X(_02058_));
 sky130_fd_sc_hd__clkinv_4 _14845_ (.A(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__a31o_1 _14846_ (.A1(net1738),
    .A2(\localMemoryInterface.lastWBByteSelect[1] ),
    .A3(_02059_),
    .B1(net1909),
    .X(_02060_));
 sky130_fd_sc_hd__a21oi_4 _14847_ (.A1(_02057_),
    .A2(_02060_),
    .B1(net488),
    .Y(_02061_));
 sky130_fd_sc_hd__a211o_1 _14848_ (.A1(net416),
    .A2(net494),
    .B1(_02061_),
    .C1(net1894),
    .X(_00728_));
 sky130_fd_sc_hd__or2_1 _14849_ (.A(\core.csr.currentInstruction[16] ),
    .B(net936),
    .X(_02062_));
 sky130_fd_sc_hd__a221o_1 _14850_ (.A1(net1020),
    .A2(_08145_),
    .B1(net933),
    .B2(\core.registers[0][16] ),
    .C1(net939),
    .X(_02063_));
 sky130_fd_sc_hd__a21o_1 _14851_ (.A1(_02062_),
    .A2(_02063_),
    .B1(net945),
    .X(_02064_));
 sky130_fd_sc_hd__and4_4 _14852_ (.A(\wbSRAMInterface.currentByteSelect[2] ),
    .B(net1614),
    .C(net1230),
    .D(_07042_),
    .X(_02065_));
 sky130_fd_sc_hd__o211a_1 _14853_ (.A1(net1747),
    .A2(net943),
    .B1(_02064_),
    .C1(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__and4_1 _14854_ (.A(\wbSRAMInterface.currentByteSelect[2] ),
    .B(net1614),
    .C(net1230),
    .D(_07044_),
    .X(_02067_));
 sky130_fd_sc_hd__o21ai_4 _14855_ (.A1(net672),
    .A2(_02066_),
    .B1(net1276),
    .Y(_02068_));
 sky130_fd_sc_hd__mux2_2 _14856_ (.A0(net50),
    .A1(net85),
    .S(net1743),
    .X(_02069_));
 sky130_fd_sc_hd__clkinv_4 _14857_ (.A(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__a31o_1 _14858_ (.A1(net1738),
    .A2(\localMemoryInterface.lastWBByteSelect[2] ),
    .A3(_02070_),
    .B1(net1907),
    .X(_02071_));
 sky130_fd_sc_hd__a21oi_4 _14859_ (.A1(_02068_),
    .A2(_02071_),
    .B1(net488),
    .Y(_02072_));
 sky130_fd_sc_hd__a211o_1 _14860_ (.A1(net417),
    .A2(net494),
    .B1(_02072_),
    .C1(net1894),
    .X(_00729_));
 sky130_fd_sc_hd__or2_1 _14861_ (.A(\core.csr.currentInstruction[17] ),
    .B(net936),
    .X(_02073_));
 sky130_fd_sc_hd__a221o_1 _14862_ (.A1(net1019),
    .A2(_08190_),
    .B1(net933),
    .B2(\core.registers[0][17] ),
    .C1(net939),
    .X(_02074_));
 sky130_fd_sc_hd__a21o_1 _14863_ (.A1(_02073_),
    .A2(_02074_),
    .B1(net945),
    .X(_02075_));
 sky130_fd_sc_hd__o211a_2 _14864_ (.A1(net458),
    .A2(net943),
    .B1(_02065_),
    .C1(_02075_),
    .X(_02076_));
 sky130_fd_sc_hd__o21ai_4 _14865_ (.A1(net672),
    .A2(_02076_),
    .B1(net1276),
    .Y(_02077_));
 sky130_fd_sc_hd__mux2_2 _14866_ (.A0(net51),
    .A1(net86),
    .S(net1743),
    .X(_02078_));
 sky130_fd_sc_hd__clkinv_4 _14867_ (.A(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__a31o_1 _14868_ (.A1(net1740),
    .A2(\localMemoryInterface.lastWBByteSelect[2] ),
    .A3(_02079_),
    .B1(net1907),
    .X(_02080_));
 sky130_fd_sc_hd__a21oi_4 _14869_ (.A1(_02077_),
    .A2(_02080_),
    .B1(net488),
    .Y(_02081_));
 sky130_fd_sc_hd__a211o_1 _14870_ (.A1(net418),
    .A2(net494),
    .B1(_02081_),
    .C1(net1896),
    .X(_00730_));
 sky130_fd_sc_hd__or2_1 _14871_ (.A(\core.csr.currentInstruction[18] ),
    .B(net937),
    .X(_02082_));
 sky130_fd_sc_hd__a221o_1 _14872_ (.A1(net1019),
    .A2(_08211_),
    .B1(net935),
    .B2(\core.registers[0][18] ),
    .C1(net941),
    .X(_02083_));
 sky130_fd_sc_hd__a21o_1 _14873_ (.A1(_02082_),
    .A2(_02083_),
    .B1(net946),
    .X(_02084_));
 sky130_fd_sc_hd__o211a_1 _14874_ (.A1(net459),
    .A2(net942),
    .B1(_02065_),
    .C1(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__o21ai_2 _14875_ (.A1(net673),
    .A2(_02085_),
    .B1(net1277),
    .Y(_02086_));
 sky130_fd_sc_hd__mux2_2 _14876_ (.A0(net52),
    .A1(net88),
    .S(net1743),
    .X(_02087_));
 sky130_fd_sc_hd__clkinv_4 _14877_ (.A(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__a31o_1 _14878_ (.A1(net1738),
    .A2(\localMemoryInterface.lastWBByteSelect[2] ),
    .A3(_02088_),
    .B1(net1907),
    .X(_02089_));
 sky130_fd_sc_hd__a21oi_4 _14879_ (.A1(_02086_),
    .A2(_02089_),
    .B1(net488),
    .Y(_02090_));
 sky130_fd_sc_hd__a211o_1 _14880_ (.A1(net419),
    .A2(net494),
    .B1(_02090_),
    .C1(net1895),
    .X(_00731_));
 sky130_fd_sc_hd__a221o_1 _14881_ (.A1(net1019),
    .A2(_08244_),
    .B1(net933),
    .B2(\core.registers[0][19] ),
    .C1(net939),
    .X(_02091_));
 sky130_fd_sc_hd__o21a_1 _14882_ (.A1(\core.csr.currentInstruction[19] ),
    .A2(net936),
    .B1(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__mux2_2 _14883_ (.A0(net460),
    .A1(_02092_),
    .S(net943),
    .X(_02093_));
 sky130_fd_sc_hd__a21oi_1 _14884_ (.A1(_02067_),
    .A2(_02093_),
    .B1(_01952_),
    .Y(_02094_));
 sky130_fd_sc_hd__a21bo_1 _14885_ (.A1(_07005_),
    .A2(_02094_),
    .B1_N(net1278),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_2 _14886_ (.A0(net53),
    .A1(net89),
    .S(net1743),
    .X(_02096_));
 sky130_fd_sc_hd__clkinv_4 _14887_ (.A(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__a31o_2 _14888_ (.A1(net1739),
    .A2(\localMemoryInterface.lastWBByteSelect[2] ),
    .A3(_02097_),
    .B1(net1907),
    .X(_02098_));
 sky130_fd_sc_hd__a21oi_4 _14889_ (.A1(_02095_),
    .A2(_02098_),
    .B1(net492),
    .Y(_02099_));
 sky130_fd_sc_hd__a211o_1 _14890_ (.A1(net420),
    .A2(net493),
    .B1(_02099_),
    .C1(net1895),
    .X(_00732_));
 sky130_fd_sc_hd__a221o_1 _14891_ (.A1(net1019),
    .A2(_08276_),
    .B1(net933),
    .B2(\core.registers[0][20] ),
    .C1(net939),
    .X(_02100_));
 sky130_fd_sc_hd__o21a_1 _14892_ (.A1(\core.csr.currentInstruction[20] ),
    .A2(net936),
    .B1(_02100_),
    .X(_02101_));
 sky130_fd_sc_hd__mux2_4 _14893_ (.A0(net462),
    .A1(_02101_),
    .S(net943),
    .X(_02102_));
 sky130_fd_sc_hd__a21oi_2 _14894_ (.A1(_02067_),
    .A2(_02102_),
    .B1(_01952_),
    .Y(_02103_));
 sky130_fd_sc_hd__a21bo_1 _14895_ (.A1(_07005_),
    .A2(_02103_),
    .B1_N(net1279),
    .X(_02104_));
 sky130_fd_sc_hd__mux2_2 _14896_ (.A0(net55),
    .A1(net90),
    .S(net1743),
    .X(_02105_));
 sky130_fd_sc_hd__clkinv_4 _14897_ (.A(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__a31o_2 _14898_ (.A1(net1739),
    .A2(\localMemoryInterface.lastWBByteSelect[2] ),
    .A3(_02106_),
    .B1(net1907),
    .X(_02107_));
 sky130_fd_sc_hd__a21oi_4 _14899_ (.A1(_02104_),
    .A2(_02107_),
    .B1(net490),
    .Y(_02108_));
 sky130_fd_sc_hd__a211o_1 _14900_ (.A1(net422),
    .A2(net493),
    .B1(_02108_),
    .C1(net1895),
    .X(_00733_));
 sky130_fd_sc_hd__or2_1 _14901_ (.A(\core.csr.currentInstruction[21] ),
    .B(net936),
    .X(_02109_));
 sky130_fd_sc_hd__a221o_1 _14902_ (.A1(net1019),
    .A2(_08317_),
    .B1(net933),
    .B2(\core.registers[0][21] ),
    .C1(net939),
    .X(_02110_));
 sky130_fd_sc_hd__a21o_1 _14903_ (.A1(_02109_),
    .A2(_02110_),
    .B1(net945),
    .X(_02111_));
 sky130_fd_sc_hd__o211a_2 _14904_ (.A1(net463),
    .A2(net943),
    .B1(_02065_),
    .C1(_02111_),
    .X(_02112_));
 sky130_fd_sc_hd__o21ai_2 _14905_ (.A1(net674),
    .A2(_02112_),
    .B1(net1278),
    .Y(_02113_));
 sky130_fd_sc_hd__mux2_2 _14906_ (.A0(net56),
    .A1(net91),
    .S(net1743),
    .X(_02114_));
 sky130_fd_sc_hd__clkinv_4 _14907_ (.A(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__a31o_1 _14908_ (.A1(net1739),
    .A2(\localMemoryInterface.lastWBByteSelect[2] ),
    .A3(_02115_),
    .B1(net1907),
    .X(_02116_));
 sky130_fd_sc_hd__a21oi_4 _14909_ (.A1(_02113_),
    .A2(_02116_),
    .B1(net490),
    .Y(_02117_));
 sky130_fd_sc_hd__a211o_1 _14910_ (.A1(net423),
    .A2(net493),
    .B1(_02117_),
    .C1(net1896),
    .X(_00734_));
 sky130_fd_sc_hd__or2_1 _14911_ (.A(\core.csr.currentInstruction[22] ),
    .B(net937),
    .X(_02118_));
 sky130_fd_sc_hd__a221o_1 _14912_ (.A1(net1020),
    .A2(_08339_),
    .B1(net935),
    .B2(\core.registers[0][22] ),
    .C1(net941),
    .X(_02119_));
 sky130_fd_sc_hd__a21o_1 _14913_ (.A1(_02118_),
    .A2(_02119_),
    .B1(net946),
    .X(_02120_));
 sky130_fd_sc_hd__o211a_1 _14914_ (.A1(net464),
    .A2(net942),
    .B1(_02065_),
    .C1(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__o21ai_2 _14915_ (.A1(net674),
    .A2(_02121_),
    .B1(net1278),
    .Y(_02122_));
 sky130_fd_sc_hd__mux2_2 _14916_ (.A0(net57),
    .A1(net92),
    .S(net1743),
    .X(_02123_));
 sky130_fd_sc_hd__clkinv_4 _14917_ (.A(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__a31o_1 _14918_ (.A1(net1739),
    .A2(\localMemoryInterface.lastWBByteSelect[2] ),
    .A3(_02124_),
    .B1(net1907),
    .X(_02125_));
 sky130_fd_sc_hd__a21oi_4 _14919_ (.A1(_02122_),
    .A2(_02125_),
    .B1(net489),
    .Y(_02126_));
 sky130_fd_sc_hd__a211o_1 _14920_ (.A1(net424),
    .A2(net493),
    .B1(_02126_),
    .C1(net1902),
    .X(_00735_));
 sky130_fd_sc_hd__or2_1 _14921_ (.A(\core.csr.currentInstruction[23] ),
    .B(net936),
    .X(_02127_));
 sky130_fd_sc_hd__a221o_1 _14922_ (.A1(net1019),
    .A2(_08370_),
    .B1(net933),
    .B2(\core.registers[0][23] ),
    .C1(net939),
    .X(_02128_));
 sky130_fd_sc_hd__a21o_1 _14923_ (.A1(_02127_),
    .A2(_02128_),
    .B1(net945),
    .X(_02129_));
 sky130_fd_sc_hd__o211a_2 _14924_ (.A1(net465),
    .A2(net943),
    .B1(_02065_),
    .C1(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__o21ai_2 _14925_ (.A1(net674),
    .A2(_02130_),
    .B1(net1278),
    .Y(_02131_));
 sky130_fd_sc_hd__mux2_2 _14926_ (.A0(net58),
    .A1(net93),
    .S(net1743),
    .X(_02132_));
 sky130_fd_sc_hd__clkinv_4 _14927_ (.A(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__a31o_1 _14928_ (.A1(net1739),
    .A2(\localMemoryInterface.lastWBByteSelect[2] ),
    .A3(_02133_),
    .B1(net1908),
    .X(_02134_));
 sky130_fd_sc_hd__a21oi_4 _14929_ (.A1(_02131_),
    .A2(_02134_),
    .B1(net489),
    .Y(_02135_));
 sky130_fd_sc_hd__a211o_1 _14930_ (.A1(net425),
    .A2(net493),
    .B1(_02135_),
    .C1(net1902),
    .X(_00736_));
 sky130_fd_sc_hd__or2_1 _14931_ (.A(\core.csr.currentInstruction[24] ),
    .B(net936),
    .X(_02136_));
 sky130_fd_sc_hd__a221o_1 _14932_ (.A1(net1019),
    .A2(_08401_),
    .B1(net933),
    .B2(\core.registers[0][24] ),
    .C1(net939),
    .X(_02137_));
 sky130_fd_sc_hd__a21o_1 _14933_ (.A1(_02136_),
    .A2(_02137_),
    .B1(net945),
    .X(_02138_));
 sky130_fd_sc_hd__and4_4 _14934_ (.A(\wbSRAMInterface.currentByteSelect[3] ),
    .B(net1614),
    .C(net1230),
    .D(_07042_),
    .X(_02139_));
 sky130_fd_sc_hd__o211a_2 _14935_ (.A1(net466),
    .A2(net943),
    .B1(_02138_),
    .C1(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__o21ai_2 _14936_ (.A1(net674),
    .A2(_02140_),
    .B1(net1278),
    .Y(_02141_));
 sky130_fd_sc_hd__mux2_2 _14937_ (.A0(net59),
    .A1(net94),
    .S(net1743),
    .X(_02142_));
 sky130_fd_sc_hd__clkinv_4 _14938_ (.A(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__a31o_1 _14939_ (.A1(net1739),
    .A2(\localMemoryInterface.lastWBByteSelect[3] ),
    .A3(_02143_),
    .B1(net1910),
    .X(_02144_));
 sky130_fd_sc_hd__a21oi_4 _14940_ (.A1(_02141_),
    .A2(_02144_),
    .B1(net490),
    .Y(_02145_));
 sky130_fd_sc_hd__a211o_1 _14941_ (.A1(net426),
    .A2(_01896_),
    .B1(_02145_),
    .C1(net1902),
    .X(_00737_));
 sky130_fd_sc_hd__or2_1 _14942_ (.A(\core.csr.currentInstruction[25] ),
    .B(net936),
    .X(_02146_));
 sky130_fd_sc_hd__a221o_1 _14943_ (.A1(net1019),
    .A2(_08433_),
    .B1(net933),
    .B2(\core.registers[0][25] ),
    .C1(net939),
    .X(_02147_));
 sky130_fd_sc_hd__a21o_1 _14944_ (.A1(_02146_),
    .A2(_02147_),
    .B1(net945),
    .X(_02148_));
 sky130_fd_sc_hd__o211a_2 _14945_ (.A1(net467),
    .A2(net943),
    .B1(_02139_),
    .C1(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__o21ai_2 _14946_ (.A1(net674),
    .A2(_02149_),
    .B1(net1278),
    .Y(_02150_));
 sky130_fd_sc_hd__mux2_2 _14947_ (.A0(net60),
    .A1(net95),
    .S(net1743),
    .X(_02151_));
 sky130_fd_sc_hd__clkinv_4 _14948_ (.A(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__a31o_1 _14949_ (.A1(net1739),
    .A2(\localMemoryInterface.lastWBByteSelect[3] ),
    .A3(_02152_),
    .B1(net1910),
    .X(_02153_));
 sky130_fd_sc_hd__a21oi_4 _14950_ (.A1(_02150_),
    .A2(_02153_),
    .B1(net489),
    .Y(_02154_));
 sky130_fd_sc_hd__a211o_1 _14951_ (.A1(net427),
    .A2(net493),
    .B1(_02154_),
    .C1(net1902),
    .X(_00738_));
 sky130_fd_sc_hd__or2_1 _14952_ (.A(\core.csr.currentInstruction[26] ),
    .B(net938),
    .X(_02155_));
 sky130_fd_sc_hd__a221o_1 _14953_ (.A1(net1022),
    .A2(_08464_),
    .B1(net934),
    .B2(\core.registers[0][26] ),
    .C1(net940),
    .X(_02156_));
 sky130_fd_sc_hd__a21o_1 _14954_ (.A1(_02155_),
    .A2(_02156_),
    .B1(net948),
    .X(_02157_));
 sky130_fd_sc_hd__o211a_1 _14955_ (.A1(net468),
    .A2(net944),
    .B1(_02139_),
    .C1(_02157_),
    .X(_02158_));
 sky130_fd_sc_hd__o21ai_2 _14956_ (.A1(net674),
    .A2(_02158_),
    .B1(net1279),
    .Y(_02159_));
 sky130_fd_sc_hd__mux2_2 _14957_ (.A0(net61),
    .A1(net96),
    .S(net1744),
    .X(_02160_));
 sky130_fd_sc_hd__clkinv_4 _14958_ (.A(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__a31o_1 _14959_ (.A1(net1739),
    .A2(\localMemoryInterface.lastWBByteSelect[3] ),
    .A3(_02161_),
    .B1(net1910),
    .X(_02162_));
 sky130_fd_sc_hd__a21oi_4 _14960_ (.A1(_02159_),
    .A2(_02162_),
    .B1(net490),
    .Y(_02163_));
 sky130_fd_sc_hd__a211o_1 _14961_ (.A1(net428),
    .A2(net493),
    .B1(_02163_),
    .C1(net1902),
    .X(_00739_));
 sky130_fd_sc_hd__or2_1 _14962_ (.A(\core.csr.currentInstruction[27] ),
    .B(net938),
    .X(_02164_));
 sky130_fd_sc_hd__a221o_1 _14963_ (.A1(net1021),
    .A2(_08506_),
    .B1(net934),
    .B2(\core.registers[0][27] ),
    .C1(net941),
    .X(_02165_));
 sky130_fd_sc_hd__a21o_1 _14964_ (.A1(_02164_),
    .A2(_02165_),
    .B1(net947),
    .X(_02166_));
 sky130_fd_sc_hd__o211a_1 _14965_ (.A1(net469),
    .A2(_01900_),
    .B1(_02139_),
    .C1(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__o21ai_2 _14966_ (.A1(net675),
    .A2(_02167_),
    .B1(net1278),
    .Y(_02168_));
 sky130_fd_sc_hd__mux2_2 _14967_ (.A0(net62),
    .A1(net97),
    .S(net1744),
    .X(_02169_));
 sky130_fd_sc_hd__clkinv_4 _14968_ (.A(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__a31o_1 _14969_ (.A1(net1739),
    .A2(\localMemoryInterface.lastWBByteSelect[3] ),
    .A3(_02170_),
    .B1(net1910),
    .X(_02171_));
 sky130_fd_sc_hd__a21oi_4 _14970_ (.A1(_02168_),
    .A2(_02171_),
    .B1(net490),
    .Y(_02172_));
 sky130_fd_sc_hd__a211o_1 _14971_ (.A1(net429),
    .A2(net493),
    .B1(_02172_),
    .C1(net1903),
    .X(_00740_));
 sky130_fd_sc_hd__or2_1 _14972_ (.A(\core.csr.currentInstruction[28] ),
    .B(net938),
    .X(_02173_));
 sky130_fd_sc_hd__a221o_1 _14973_ (.A1(net1022),
    .A2(_08530_),
    .B1(net934),
    .B2(\core.registers[0][28] ),
    .C1(net941),
    .X(_02174_));
 sky130_fd_sc_hd__a21o_1 _14974_ (.A1(_02173_),
    .A2(_02174_),
    .B1(net948),
    .X(_02175_));
 sky130_fd_sc_hd__o211a_1 _14975_ (.A1(net470),
    .A2(_01900_),
    .B1(_02139_),
    .C1(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__o21ai_2 _14976_ (.A1(net675),
    .A2(_02176_),
    .B1(net1278),
    .Y(_02177_));
 sky130_fd_sc_hd__mux2_2 _14977_ (.A0(net63),
    .A1(net99),
    .S(net1744),
    .X(_02178_));
 sky130_fd_sc_hd__clkinv_4 _14978_ (.A(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__a31o_2 _14979_ (.A1(net1739),
    .A2(\localMemoryInterface.lastWBByteSelect[3] ),
    .A3(_02179_),
    .B1(net1910),
    .X(_02180_));
 sky130_fd_sc_hd__a21oi_4 _14980_ (.A1(_02177_),
    .A2(_02180_),
    .B1(net490),
    .Y(_02181_));
 sky130_fd_sc_hd__a211o_1 _14981_ (.A1(net430),
    .A2(net493),
    .B1(_02181_),
    .C1(net1903),
    .X(_00741_));
 sky130_fd_sc_hd__or2_1 _14982_ (.A(\core.csr.currentInstruction[29] ),
    .B(net938),
    .X(_02182_));
 sky130_fd_sc_hd__a221o_1 _14983_ (.A1(net1021),
    .A2(_08559_),
    .B1(net935),
    .B2(\core.registers[0][29] ),
    .C1(net940),
    .X(_02183_));
 sky130_fd_sc_hd__a21o_1 _14984_ (.A1(_02182_),
    .A2(_02183_),
    .B1(net948),
    .X(_02184_));
 sky130_fd_sc_hd__o211a_1 _14985_ (.A1(net471),
    .A2(_01900_),
    .B1(_02139_),
    .C1(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__o21ai_2 _14986_ (.A1(net675),
    .A2(_02185_),
    .B1(net1278),
    .Y(_02186_));
 sky130_fd_sc_hd__mux2_2 _14987_ (.A0(net64),
    .A1(net100),
    .S(net1744),
    .X(_02187_));
 sky130_fd_sc_hd__clkinv_4 _14988_ (.A(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__a31o_1 _14989_ (.A1(net1740),
    .A2(\localMemoryInterface.lastWBByteSelect[3] ),
    .A3(_02188_),
    .B1(net1910),
    .X(_02189_));
 sky130_fd_sc_hd__a21oi_4 _14990_ (.A1(_02186_),
    .A2(_02189_),
    .B1(net490),
    .Y(_02190_));
 sky130_fd_sc_hd__a211o_1 _14991_ (.A1(net431),
    .A2(net494),
    .B1(_02190_),
    .C1(net1903),
    .X(_00742_));
 sky130_fd_sc_hd__a22o_1 _14992_ (.A1(net1021),
    .A2(_08600_),
    .B1(_01912_),
    .B2(\core.registers[0][30] ),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _14993_ (.A0(\core.csr.currentInstruction[30] ),
    .A1(_02191_),
    .S(_01909_),
    .X(_02192_));
 sky130_fd_sc_hd__or2_1 _14994_ (.A(net473),
    .B(net944),
    .X(_02193_));
 sky130_fd_sc_hd__o211a_1 _14995_ (.A1(net948),
    .A2(_02192_),
    .B1(_02193_),
    .C1(_02139_),
    .X(_02194_));
 sky130_fd_sc_hd__o21ai_2 _14996_ (.A1(net675),
    .A2(_02194_),
    .B1(net1279),
    .Y(_02195_));
 sky130_fd_sc_hd__mux2_2 _14997_ (.A0(net66),
    .A1(net101),
    .S(net1744),
    .X(_02196_));
 sky130_fd_sc_hd__clkinv_4 _14998_ (.A(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__a31o_1 _14999_ (.A1(net1740),
    .A2(\localMemoryInterface.lastWBByteSelect[3] ),
    .A3(_02197_),
    .B1(net1910),
    .X(_02198_));
 sky130_fd_sc_hd__a21oi_4 _15000_ (.A1(_02195_),
    .A2(_02198_),
    .B1(net490),
    .Y(_02199_));
 sky130_fd_sc_hd__a211o_1 _15001_ (.A1(net433),
    .A2(net494),
    .B1(_02199_),
    .C1(net1902),
    .X(_00743_));
 sky130_fd_sc_hd__or2_1 _15002_ (.A(\core.csr.currentInstruction[31] ),
    .B(net936),
    .X(_02200_));
 sky130_fd_sc_hd__a221o_1 _15003_ (.A1(net1019),
    .A2(_08625_),
    .B1(net933),
    .B2(\core.registers[0][31] ),
    .C1(net939),
    .X(_02201_));
 sky130_fd_sc_hd__a21o_1 _15004_ (.A1(_02200_),
    .A2(_02201_),
    .B1(net945),
    .X(_02202_));
 sky130_fd_sc_hd__o211a_2 _15005_ (.A1(net474),
    .A2(net943),
    .B1(_02139_),
    .C1(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__o21ai_2 _15006_ (.A1(net674),
    .A2(_02203_),
    .B1(net1278),
    .Y(_02204_));
 sky130_fd_sc_hd__mux2_2 _15007_ (.A0(net67),
    .A1(net102),
    .S(net1744),
    .X(_02205_));
 sky130_fd_sc_hd__clkinv_4 _15008_ (.A(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__a31o_2 _15009_ (.A1(net1740),
    .A2(\localMemoryInterface.lastWBByteSelect[3] ),
    .A3(_02206_),
    .B1(net205),
    .X(_02207_));
 sky130_fd_sc_hd__a21oi_4 _15010_ (.A1(_02204_),
    .A2(_02207_),
    .B1(net490),
    .Y(_02208_));
 sky130_fd_sc_hd__a211o_1 _15011_ (.A1(net434),
    .A2(net493),
    .B1(_02208_),
    .C1(net1896),
    .X(_00744_));
 sky130_fd_sc_hd__a211oi_1 _15012_ (.A1(_03822_),
    .A2(_01895_),
    .B1(_06697_),
    .C1(net1880),
    .Y(_00745_));
 sky130_fd_sc_hd__nand2_1 _15013_ (.A(net251),
    .B(net214),
    .Y(_02209_));
 sky130_fd_sc_hd__nor3_1 _15014_ (.A(net1880),
    .B(net1614),
    .C(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__mux2_1 _15015_ (.A0(\wbSRAMInterface.currentAddress[0] ),
    .A1(net190),
    .S(net1287),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _15016_ (.A0(\wbSRAMInterface.currentAddress[1] ),
    .A1(net201),
    .S(net1287),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _15017_ (.A0(\wbSRAMInterface.currentAddress[2] ),
    .A1(net206),
    .S(net1287),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _15018_ (.A0(\wbSRAMInterface.currentAddress[3] ),
    .A1(net207),
    .S(net1287),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _15019_ (.A0(\wbSRAMInterface.currentAddress[4] ),
    .A1(net208),
    .S(net1287),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _15020_ (.A0(\wbSRAMInterface.currentAddress[5] ),
    .A1(net209),
    .S(net1288),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _15021_ (.A0(\wbSRAMInterface.currentAddress[6] ),
    .A1(net210),
    .S(net1288),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _15022_ (.A0(\wbSRAMInterface.currentAddress[7] ),
    .A1(net211),
    .S(net1288),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _15023_ (.A0(\wbSRAMInterface.currentAddress[8] ),
    .A1(net212),
    .S(net1288),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _15024_ (.A0(\wbSRAMInterface.currentAddress[9] ),
    .A1(net213),
    .S(net1288),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _15025_ (.A0(\wbSRAMInterface.currentAddress[10] ),
    .A1(net191),
    .S(net1289),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _15026_ (.A0(\wbSRAMInterface.currentAddress[11] ),
    .A1(net192),
    .S(net1289),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _15027_ (.A0(\wbSRAMInterface.currentAddress[12] ),
    .A1(net193),
    .S(net1289),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _15028_ (.A0(\wbSRAMInterface.currentAddress[13] ),
    .A1(net194),
    .S(net1289),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _15029_ (.A0(\wbSRAMInterface.currentAddress[14] ),
    .A1(net195),
    .S(net1289),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _15030_ (.A0(\wbSRAMInterface.currentAddress[15] ),
    .A1(net196),
    .S(net1290),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _15031_ (.A0(\wbSRAMInterface.currentAddress[16] ),
    .A1(net197),
    .S(net1289),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _15032_ (.A0(\wbSRAMInterface.currentAddress[17] ),
    .A1(net198),
    .S(net1289),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _15033_ (.A0(\wbSRAMInterface.currentAddress[18] ),
    .A1(net199),
    .S(net1289),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _15034_ (.A0(\wbSRAMInterface.currentAddress[19] ),
    .A1(net200),
    .S(net1289),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _15035_ (.A0(\wbSRAMInterface.currentAddress[20] ),
    .A1(net202),
    .S(net1290),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _15036_ (.A0(\wbSRAMInterface.currentAddress[21] ),
    .A1(net203),
    .S(net1290),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _15037_ (.A0(\wbSRAMInterface.currentAddress[22] ),
    .A1(net204),
    .S(net1290),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _15038_ (.A0(\wbSRAMInterface.currentAddress[23] ),
    .A1(net205),
    .S(net1289),
    .X(_00769_));
 sky130_fd_sc_hd__and2_4 _15039_ (.A(net1805),
    .B(_06709_),
    .X(_00770_));
 sky130_fd_sc_hd__a41o_1 _15040_ (.A1(net442),
    .A2(net1849),
    .A3(net1615),
    .A4(_06696_),
    .B1(net1287),
    .X(_00771_));
 sky130_fd_sc_hd__a31o_1 _15041_ (.A1(net251),
    .A2(net214),
    .A3(net252),
    .B1(net1615),
    .X(_02211_));
 sky130_fd_sc_hd__o21ai_1 _15042_ (.A1(\wbSRAMInterface.state[0] ),
    .A2(_01895_),
    .B1(\wbSRAMInterface.state[1] ),
    .Y(_02212_));
 sky130_fd_sc_hd__and3_1 _15043_ (.A(net1849),
    .B(_02211_),
    .C(_02212_),
    .X(_00772_));
 sky130_fd_sc_hd__o21ba_1 _15044_ (.A1(net252),
    .A2(_02209_),
    .B1_N(net1614),
    .X(_02213_));
 sky130_fd_sc_hd__a211o_1 _15045_ (.A1(\wbSRAMInterface.state[1] ),
    .A2(\wbSRAMInterface.state[0] ),
    .B1(net1880),
    .C1(_02213_),
    .X(_02214_));
 sky130_fd_sc_hd__a21oi_1 _15046_ (.A1(\wbSRAMInterface.state[0] ),
    .A2(_01895_),
    .B1(_02214_),
    .Y(_00773_));
 sky130_fd_sc_hd__nor2_8 _15047_ (.A(_06849_),
    .B(_07061_),
    .Y(_02215_));
 sky130_fd_sc_hd__mux2_1 _15048_ (.A0(\core.registers[16][0] ),
    .A1(net1078),
    .S(net1012),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _15049_ (.A0(\core.registers[16][1] ),
    .A1(net1083),
    .S(net1014),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _15050_ (.A0(\core.registers[16][2] ),
    .A1(net1085),
    .S(net1012),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _15051_ (.A0(\core.registers[16][3] ),
    .A1(net1091),
    .S(net1011),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _15052_ (.A0(\core.registers[16][4] ),
    .A1(net1027),
    .S(net1014),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _15053_ (.A0(\core.registers[16][5] ),
    .A1(net1033),
    .S(net1014),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _15054_ (.A0(\core.registers[16][6] ),
    .A1(net1035),
    .S(net1014),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _15055_ (.A0(\core.registers[16][7] ),
    .A1(net1139),
    .S(net1014),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _15056_ (.A0(\core.registers[16][8] ),
    .A1(net898),
    .S(net1013),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _15057_ (.A0(\core.registers[16][9] ),
    .A1(net902),
    .S(net1013),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _15058_ (.A0(\core.registers[16][10] ),
    .A1(net759),
    .S(net1013),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _15059_ (.A0(\core.registers[16][11] ),
    .A1(net762),
    .S(net1013),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _15060_ (.A0(\core.registers[16][12] ),
    .A1(net729),
    .S(net1014),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _15061_ (.A0(\core.registers[16][13] ),
    .A1(net733),
    .S(net1013),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _15062_ (.A0(\core.registers[16][14] ),
    .A1(net738),
    .S(net1011),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _15063_ (.A0(\core.registers[16][15] ),
    .A1(net740),
    .S(net1012),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _15064_ (.A0(\core.registers[16][16] ),
    .A1(net830),
    .S(net1012),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _15065_ (.A0(\core.registers[16][17] ),
    .A1(net835),
    .S(net1011),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _15066_ (.A0(\core.registers[16][18] ),
    .A1(net838),
    .S(net1013),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _15067_ (.A0(\core.registers[16][19] ),
    .A1(net844),
    .S(net1011),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _15068_ (.A0(\core.registers[16][20] ),
    .A1(net847),
    .S(net1011),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _15069_ (.A0(\core.registers[16][21] ),
    .A1(net852),
    .S(net1011),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _15070_ (.A0(\core.registers[16][22] ),
    .A1(net857),
    .S(net1012),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _15071_ (.A0(\core.registers[16][23] ),
    .A1(net862),
    .S(net1011),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _15072_ (.A0(\core.registers[16][24] ),
    .A1(net994),
    .S(net1011),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _15073_ (.A0(\core.registers[16][25] ),
    .A1(net998),
    .S(net1011),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _15074_ (.A0(\core.registers[16][26] ),
    .A1(net1003),
    .S(net1013),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _15075_ (.A0(\core.registers[16][27] ),
    .A1(net867),
    .S(net1013),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _15076_ (.A0(\core.registers[16][28] ),
    .A1(net871),
    .S(net1014),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _15077_ (.A0(\core.registers[16][29] ),
    .A1(net874),
    .S(net1013),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _15078_ (.A0(\core.registers[16][30] ),
    .A1(net879),
    .S(net1013),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _15079_ (.A0(\core.registers[16][31] ),
    .A1(net1023),
    .S(net1011),
    .X(_00805_));
 sky130_fd_sc_hd__nor2_1 _15080_ (.A(_04070_),
    .B(_06648_),
    .Y(_02216_));
 sky130_fd_sc_hd__or2_2 _15081_ (.A(_04070_),
    .B(_06648_),
    .X(_02217_));
 sky130_fd_sc_hd__or4b_2 _15082_ (.A(net1634),
    .B(_04071_),
    .C(_07003_),
    .D_N(_03861_),
    .X(_02218_));
 sky130_fd_sc_hd__nor2_2 _15083_ (.A(_07150_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__and3_1 _15084_ (.A(\core.csr.traps.mie.currentValue[20] ),
    .B(net1732),
    .C(net181),
    .X(_02220_));
 sky130_fd_sc_hd__and3_1 _15085_ (.A(\core.csr.traps.mie.currentValue[23] ),
    .B(net1732),
    .C(net184),
    .X(_02221_));
 sky130_fd_sc_hd__and3_1 _15086_ (.A(\core.csr.traps.mie.currentValue[21] ),
    .B(net1731),
    .C(net182),
    .X(_02222_));
 sky130_fd_sc_hd__and3_1 _15087_ (.A(\core.csr.traps.mie.currentValue[30] ),
    .B(net1733),
    .C(net176),
    .X(_02223_));
 sky130_fd_sc_hd__and3_1 _15088_ (.A(\core.csr.traps.mie.currentValue[27] ),
    .B(net1733),
    .C(net173),
    .X(_02224_));
 sky130_fd_sc_hd__and3_1 _15089_ (.A(\core.csr.traps.mie.currentValue[28] ),
    .B(net1732),
    .C(net174),
    .X(_02225_));
 sky130_fd_sc_hd__and3_1 _15090_ (.A(\core.csr.traps.mie.currentValue[25] ),
    .B(net1732),
    .C(net186),
    .X(_02226_));
 sky130_fd_sc_hd__and3_2 _15091_ (.A(\core.csr.traps.mie.currentValue[26] ),
    .B(net1732),
    .C(net172),
    .X(_02227_));
 sky130_fd_sc_hd__and3_1 _15092_ (.A(\core.csr.traps.mie.currentValue[19] ),
    .B(net1732),
    .C(net180),
    .X(_02228_));
 sky130_fd_sc_hd__or4_4 _15093_ (.A(_02220_),
    .B(_02225_),
    .C(_02226_),
    .D(_02227_),
    .X(_02229_));
 sky130_fd_sc_hd__a31o_1 _15094_ (.A1(\core.csr.traps.mie.currentValue[16] ),
    .A2(net1731),
    .A3(net171),
    .B1(_02222_),
    .X(_02230_));
 sky130_fd_sc_hd__a31o_1 _15095_ (.A1(\core.csr.traps.mie.currentValue[22] ),
    .A2(net1731),
    .A3(net183),
    .B1(_02230_),
    .X(_02231_));
 sky130_fd_sc_hd__a31o_1 _15096_ (.A1(\core.csr.traps.mie.currentValue[24] ),
    .A2(net1731),
    .A3(net185),
    .B1(_02224_),
    .X(_02232_));
 sky130_fd_sc_hd__a31o_1 _15097_ (.A1(\core.csr.traps.mie.currentValue[18] ),
    .A2(net1731),
    .A3(net179),
    .B1(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__a31o_1 _15098_ (.A1(\core.csr.traps.mie.currentValue[17] ),
    .A2(net1731),
    .A3(net178),
    .B1(_02233_),
    .X(_02234_));
 sky130_fd_sc_hd__a31o_1 _15099_ (.A1(\core.csr.traps.mie.currentValue[29] ),
    .A2(net1732),
    .A3(net175),
    .B1(_02228_),
    .X(_02235_));
 sky130_fd_sc_hd__a311o_1 _15100_ (.A1(\core.csr.traps.mie.currentValue[31] ),
    .A2(net1732),
    .A3(net177),
    .B1(_02221_),
    .C1(_02235_),
    .X(_02236_));
 sky130_fd_sc_hd__or4_4 _15101_ (.A(_02223_),
    .B(_02231_),
    .C(_02234_),
    .D(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__nor2_4 _15102_ (.A(_02229_),
    .B(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__nor2_4 _15103_ (.A(\core.fetchProgramCounter[1] ),
    .B(\core.fetchProgramCounter[0] ),
    .Y(_02239_));
 sky130_fd_sc_hd__or2_2 _15104_ (.A(\core.fetchProgramCounter[1] ),
    .B(\core.fetchProgramCounter[0] ),
    .X(_02240_));
 sky130_fd_sc_hd__o31ai_4 _15105_ (.A1(_08695_),
    .A2(_08696_),
    .A3(_08699_),
    .B1(_06998_),
    .Y(_02241_));
 sky130_fd_sc_hd__o22a_2 _15106_ (.A1(net1700),
    .A2(_07053_),
    .B1(net571),
    .B2(_03845_),
    .X(_02242_));
 sky130_fd_sc_hd__mux2_4 _15107_ (.A0(_04968_),
    .A1(_07490_),
    .S(net1181),
    .X(_02243_));
 sky130_fd_sc_hd__xor2_2 _15108_ (.A(_02242_),
    .B(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__o211a_2 _15109_ (.A1(_05049_),
    .A2(net1229),
    .B1(net1185),
    .C1(net1776),
    .X(_02245_));
 sky130_fd_sc_hd__and2_2 _15110_ (.A(net1179),
    .B(net570),
    .X(_02246_));
 sky130_fd_sc_hd__nand2_4 _15111_ (.A(net1179),
    .B(net570),
    .Y(_02247_));
 sky130_fd_sc_hd__nor2_4 _15112_ (.A(net1227),
    .B(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__nand2_4 _15113_ (.A(net1136),
    .B(_02241_),
    .Y(_02249_));
 sky130_fd_sc_hd__a21oi_1 _15114_ (.A1(_02244_),
    .A2(net568),
    .B1(_02245_),
    .Y(_02250_));
 sky130_fd_sc_hd__a21oi_2 _15115_ (.A1(_02244_),
    .A2(_02245_),
    .B1(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__or3b_4 _15116_ (.A(_02251_),
    .B(net1605),
    .C_N(net1102),
    .X(_02252_));
 sky130_fd_sc_hd__nor2_2 _15117_ (.A(net931),
    .B(_02252_),
    .Y(_02253_));
 sky130_fd_sc_hd__nand2_1 _15118_ (.A(net604),
    .B(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__o21ai_2 _15119_ (.A1(_03871_),
    .A2(net1606),
    .B1(net1102),
    .Y(_02255_));
 sky130_fd_sc_hd__nor2_2 _15120_ (.A(net1154),
    .B(_06648_),
    .Y(_02256_));
 sky130_fd_sc_hd__o311a_4 _15121_ (.A1(_03871_),
    .A2(net931),
    .A3(_02256_),
    .B1(net1609),
    .C1(net1103),
    .X(_02257_));
 sky130_fd_sc_hd__a211oi_4 _15122_ (.A1(net604),
    .A2(_02253_),
    .B1(_02257_),
    .C1(_02252_),
    .Y(_02258_));
 sky130_fd_sc_hd__or3b_1 _15123_ (.A(_02257_),
    .B(_02252_),
    .C_N(_02254_),
    .X(_02259_));
 sky130_fd_sc_hd__and3_4 _15124_ (.A(net1136),
    .B(net1129),
    .C(_02241_),
    .X(_02260_));
 sky130_fd_sc_hd__a21o_2 _15125_ (.A1(net554),
    .A2(net567),
    .B1(net596),
    .X(_02261_));
 sky130_fd_sc_hd__a31o_1 _15126_ (.A1(_07047_),
    .A2(net554),
    .A3(net567),
    .B1(net596),
    .X(_02262_));
 sky130_fd_sc_hd__o21ai_4 _15127_ (.A1(net596),
    .A2(_07047_),
    .B1(_02261_),
    .Y(_02263_));
 sky130_fd_sc_hd__a2bb2o_1 _15128_ (.A1_N(_02242_),
    .A2_N(_02243_),
    .B1(_02244_),
    .B2(_02245_),
    .X(_02264_));
 sky130_fd_sc_hd__a32o_4 _15129_ (.A1(\core.pipe0_currentInstruction[9] ),
    .A2(_06998_),
    .A3(_08700_),
    .B1(net1133),
    .B2(net1767),
    .X(_02265_));
 sky130_fd_sc_hd__and2_1 _15130_ (.A(_04882_),
    .B(net1185),
    .X(_02266_));
 sky130_fd_sc_hd__a31o_1 _15131_ (.A1(net1181),
    .A2(_07569_),
    .A3(net571),
    .B1(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__and2_4 _15132_ (.A(net1221),
    .B(net570),
    .X(_02268_));
 sky130_fd_sc_hd__nand2_8 _15133_ (.A(net1221),
    .B(net570),
    .Y(_02269_));
 sky130_fd_sc_hd__o2bb2a_2 _15134_ (.A1_N(net1226),
    .A2_N(_02267_),
    .B1(net566),
    .B2(net472),
    .X(_02270_));
 sky130_fd_sc_hd__xor2_2 _15135_ (.A(_02265_),
    .B(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__nor2_1 _15136_ (.A(_02264_),
    .B(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__and2_1 _15137_ (.A(_02264_),
    .B(_02271_),
    .X(_02273_));
 sky130_fd_sc_hd__or3_1 _15138_ (.A(net562),
    .B(_02272_),
    .C(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__o211a_1 _15139_ (.A1(\core.fetchProgramCounter[2] ),
    .A2(net568),
    .B1(_02274_),
    .C1(net1128),
    .X(_02275_));
 sky130_fd_sc_hd__nor2_1 _15140_ (.A(\core.csr.trapReturnVector[2] ),
    .B(net1128),
    .Y(_02276_));
 sky130_fd_sc_hd__nor3b_4 _15141_ (.A(\core.csr.traps.mtvec.csrReadData[1] ),
    .B(net1103),
    .C_N(\core.csr.traps.mtvec.csrReadData[0] ),
    .Y(_02277_));
 sky130_fd_sc_hd__a21oi_1 _15142_ (.A1(\core.csr.traps.mcause.csrReadData[0] ),
    .A2(net1057),
    .B1(\core.csr.traps.mtvec.csrReadData[2] ),
    .Y(_02278_));
 sky130_fd_sc_hd__nand2_1 _15143_ (.A(\core.csr.traps.mtvec.csrReadData[2] ),
    .B(\core.csr.traps.mcause.csrReadData[0] ),
    .Y(_02279_));
 sky130_fd_sc_hd__and3_1 _15144_ (.A(\core.csr.traps.mtvec.csrReadData[2] ),
    .B(\core.csr.traps.mcause.csrReadData[0] ),
    .C(net1057),
    .X(_02280_));
 sky130_fd_sc_hd__or3_1 _15145_ (.A(net555),
    .B(_02278_),
    .C(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__o311a_1 _15146_ (.A1(net546),
    .A2(_02275_),
    .A3(_02276_),
    .B1(_02281_),
    .C1(net523),
    .X(_02282_));
 sky130_fd_sc_hd__nor2_1 _15147_ (.A(net1877),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__o21a_1 _15148_ (.A1(\core.fetchProgramCounter[2] ),
    .A2(net523),
    .B1(_02283_),
    .X(_00806_));
 sky130_fd_sc_hd__a21oi_1 _15149_ (.A1(_02265_),
    .A2(_02270_),
    .B1(_02273_),
    .Y(_02284_));
 sky130_fd_sc_hd__a2bb2o_1 _15150_ (.A1_N(_03844_),
    .A2_N(net572),
    .B1(net1133),
    .B2(net1762),
    .X(_02285_));
 sky130_fd_sc_hd__nor2_1 _15151_ (.A(_04801_),
    .B(net1181),
    .Y(_02286_));
 sky130_fd_sc_hd__a31o_1 _15152_ (.A1(net1181),
    .A2(_07626_),
    .A3(net571),
    .B1(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__a22o_1 _15153_ (.A1(net475),
    .A2(_02269_),
    .B1(_02287_),
    .B2(net1226),
    .X(_02288_));
 sky130_fd_sc_hd__or2_2 _15154_ (.A(_02285_),
    .B(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__nand2_1 _15155_ (.A(_02285_),
    .B(_02288_),
    .Y(_02290_));
 sky130_fd_sc_hd__and2_1 _15156_ (.A(_02289_),
    .B(_02290_),
    .X(_02291_));
 sky130_fd_sc_hd__a22o_1 _15157_ (.A1(_02265_),
    .A2(_02270_),
    .B1(_02285_),
    .B2(_02288_),
    .X(_02292_));
 sky130_fd_sc_hd__a21o_1 _15158_ (.A1(_02264_),
    .A2(_02271_),
    .B1(_02292_),
    .X(_02293_));
 sky130_fd_sc_hd__a21oi_1 _15159_ (.A1(_02284_),
    .A2(_02291_),
    .B1(net562),
    .Y(_02294_));
 sky130_fd_sc_hd__o21a_1 _15160_ (.A1(_02284_),
    .A2(_02291_),
    .B1(_02294_),
    .X(_02295_));
 sky130_fd_sc_hd__xnor2_1 _15161_ (.A(\core.fetchProgramCounter[3] ),
    .B(\core.fetchProgramCounter[2] ),
    .Y(_02296_));
 sky130_fd_sc_hd__a221o_1 _15162_ (.A1(_03812_),
    .A2(net1131),
    .B1(net567),
    .B2(_02296_),
    .C1(net544),
    .X(_02297_));
 sky130_fd_sc_hd__nor2_1 _15163_ (.A(_02295_),
    .B(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__and2_1 _15164_ (.A(\core.csr.traps.mtvec.csrReadData[3] ),
    .B(\core.csr.traps.mcause.csrReadData[1] ),
    .X(_02299_));
 sky130_fd_sc_hd__nor2_1 _15165_ (.A(\core.csr.traps.mtvec.csrReadData[3] ),
    .B(\core.csr.traps.mcause.csrReadData[1] ),
    .Y(_02300_));
 sky130_fd_sc_hd__nor2_1 _15166_ (.A(_02299_),
    .B(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__xnor2_1 _15167_ (.A(_02279_),
    .B(_02301_),
    .Y(_02302_));
 sky130_fd_sc_hd__mux2_1 _15168_ (.A0(\core.csr.traps.mtvec.csrReadData[3] ),
    .A1(_02302_),
    .S(net1057),
    .X(_02303_));
 sky130_fd_sc_hd__a211o_1 _15169_ (.A1(net544),
    .A2(_02303_),
    .B1(_02298_),
    .C1(net538),
    .X(_02304_));
 sky130_fd_sc_hd__o211a_1 _15170_ (.A1(\core.fetchProgramCounter[3] ),
    .A2(net523),
    .B1(_02304_),
    .C1(net1825),
    .X(_00807_));
 sky130_fd_sc_hd__nand2_1 _15171_ (.A(_02289_),
    .B(_02293_),
    .Y(_02305_));
 sky130_fd_sc_hd__a32o_2 _15172_ (.A1(\core.pipe0_currentInstruction[11] ),
    .A2(_06998_),
    .A3(_08700_),
    .B1(net1133),
    .B2(\core.pipe0_currentInstruction[24] ),
    .X(_02306_));
 sky130_fd_sc_hd__nor2_1 _15173_ (.A(_04719_),
    .B(net1181),
    .Y(_02307_));
 sky130_fd_sc_hd__a31oi_4 _15174_ (.A1(net1181),
    .A2(_07679_),
    .A3(net571),
    .B1(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__o22a_1 _15175_ (.A1(net1748),
    .A2(_02268_),
    .B1(_02308_),
    .B2(net1229),
    .X(_02309_));
 sky130_fd_sc_hd__o221a_1 _15176_ (.A1(net1748),
    .A2(_02268_),
    .B1(_02308_),
    .B2(net1229),
    .C1(_02306_),
    .X(_02310_));
 sky130_fd_sc_hd__xnor2_2 _15177_ (.A(_02306_),
    .B(_02309_),
    .Y(_02311_));
 sky130_fd_sc_hd__nor2_2 _15178_ (.A(_02305_),
    .B(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__and2_1 _15179_ (.A(_02305_),
    .B(_02311_),
    .X(_02313_));
 sky130_fd_sc_hd__o21a_1 _15180_ (.A1(_02312_),
    .A2(_02313_),
    .B1(_02249_),
    .X(_02314_));
 sky130_fd_sc_hd__and3_2 _15181_ (.A(\core.fetchProgramCounter[4] ),
    .B(\core.fetchProgramCounter[3] ),
    .C(\core.fetchProgramCounter[2] ),
    .X(_02315_));
 sky130_fd_sc_hd__a21oi_1 _15182_ (.A1(\core.fetchProgramCounter[3] ),
    .A2(\core.fetchProgramCounter[2] ),
    .B1(\core.fetchProgramCounter[4] ),
    .Y(_02316_));
 sky130_fd_sc_hd__or2_1 _15183_ (.A(_02315_),
    .B(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__a2bb2o_1 _15184_ (.A1_N(\core.csr.trapReturnVector[4] ),
    .A2_N(net1128),
    .B1(net567),
    .B2(_02317_),
    .X(_02318_));
 sky130_fd_sc_hd__o21ba_1 _15185_ (.A1(_02279_),
    .A2(_02300_),
    .B1_N(_02299_),
    .X(_02319_));
 sky130_fd_sc_hd__nor2_1 _15186_ (.A(\core.csr.traps.mtvec.csrReadData[4] ),
    .B(\core.csr.traps.mcause.csrReadData[2] ),
    .Y(_02320_));
 sky130_fd_sc_hd__nand2_1 _15187_ (.A(\core.csr.traps.mtvec.csrReadData[4] ),
    .B(\core.csr.traps.mcause.csrReadData[2] ),
    .Y(_02321_));
 sky130_fd_sc_hd__and2b_1 _15188_ (.A_N(_02320_),
    .B(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__xnor2_1 _15189_ (.A(_02319_),
    .B(_02322_),
    .Y(_02323_));
 sky130_fd_sc_hd__mux2_1 _15190_ (.A0(\core.csr.traps.mtvec.csrReadData[4] ),
    .A1(_02323_),
    .S(net1057),
    .X(_02324_));
 sky130_fd_sc_hd__a21o_1 _15191_ (.A1(net546),
    .A2(_02324_),
    .B1(net538),
    .X(_02325_));
 sky130_fd_sc_hd__nor3_1 _15192_ (.A(net544),
    .B(_02314_),
    .C(_02318_),
    .Y(_02326_));
 sky130_fd_sc_hd__o221a_1 _15193_ (.A1(\core.fetchProgramCounter[4] ),
    .A2(net523),
    .B1(_02325_),
    .B2(_02326_),
    .C1(net1830),
    .X(_00808_));
 sky130_fd_sc_hd__nor2_1 _15194_ (.A(_04597_),
    .B(net1181),
    .Y(_02327_));
 sky130_fd_sc_hd__a31o_1 _15195_ (.A1(net1181),
    .A2(_07727_),
    .A3(net571),
    .B1(_02327_),
    .X(_02328_));
 sky130_fd_sc_hd__a22o_1 _15196_ (.A1(net477),
    .A2(_02269_),
    .B1(_02328_),
    .B2(net1226),
    .X(_02329_));
 sky130_fd_sc_hd__and2_1 _15197_ (.A(\core.pipe0_currentInstruction[25] ),
    .B(net568),
    .X(_02330_));
 sky130_fd_sc_hd__or2_1 _15198_ (.A(_02329_),
    .B(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__xnor2_1 _15199_ (.A(_02329_),
    .B(_02330_),
    .Y(_02332_));
 sky130_fd_sc_hd__nor2_1 _15200_ (.A(_02310_),
    .B(_02312_),
    .Y(_02333_));
 sky130_fd_sc_hd__a21o_1 _15201_ (.A1(_02329_),
    .A2(_02330_),
    .B1(_02310_),
    .X(_02334_));
 sky130_fd_sc_hd__xnor2_1 _15202_ (.A(\core.csr.traps.mtvec.csrReadData[5] ),
    .B(\core.csr.traps.mcause.csrReadData[3] ),
    .Y(_02335_));
 sky130_fd_sc_hd__o21ai_2 _15203_ (.A1(_02319_),
    .A2(_02320_),
    .B1(_02321_),
    .Y(_02336_));
 sky130_fd_sc_hd__xnor2_1 _15204_ (.A(_02335_),
    .B(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__mux2_1 _15205_ (.A0(\core.csr.traps.mtvec.csrReadData[5] ),
    .A1(_02337_),
    .S(net1057),
    .X(_02338_));
 sky130_fd_sc_hd__xor2_1 _15206_ (.A(\core.fetchProgramCounter[5] ),
    .B(_02315_),
    .X(_02339_));
 sky130_fd_sc_hd__xnor2_1 _15207_ (.A(_02332_),
    .B(_02333_),
    .Y(_02340_));
 sky130_fd_sc_hd__a21oi_1 _15208_ (.A1(net1300),
    .A2(_02340_),
    .B1(net562),
    .Y(_02341_));
 sky130_fd_sc_hd__a211o_1 _15209_ (.A1(net563),
    .A2(_02339_),
    .B1(_02341_),
    .C1(net1131),
    .X(_02342_));
 sky130_fd_sc_hd__o211a_1 _15210_ (.A1(\core.csr.trapReturnVector[5] ),
    .A2(net1127),
    .B1(net556),
    .C1(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__a211o_1 _15211_ (.A1(net546),
    .A2(_02338_),
    .B1(_02343_),
    .C1(net538),
    .X(_02344_));
 sky130_fd_sc_hd__o211a_1 _15212_ (.A1(\core.fetchProgramCounter[5] ),
    .A2(net523),
    .B1(_02344_),
    .C1(net1830),
    .X(_00809_));
 sky130_fd_sc_hd__nand2_2 _15213_ (.A(\core.pipe0_currentInstruction[26] ),
    .B(net568),
    .Y(_02345_));
 sky130_fd_sc_hd__and2_1 _15214_ (.A(_04512_),
    .B(_07051_),
    .X(_02346_));
 sky130_fd_sc_hd__a31oi_4 _15215_ (.A1(net1182),
    .A2(_07752_),
    .A3(net571),
    .B1(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__a21o_1 _15216_ (.A1(net1226),
    .A2(net571),
    .B1(net478),
    .X(_02348_));
 sky130_fd_sc_hd__o21a_2 _15217_ (.A1(net1229),
    .A2(_02347_),
    .B1(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__o2111ai_4 _15218_ (.A1(net1229),
    .A2(_02347_),
    .B1(_02348_),
    .C1(net568),
    .D1(\core.pipe0_currentInstruction[26] ),
    .Y(_02350_));
 sky130_fd_sc_hd__xnor2_4 _15219_ (.A(_02345_),
    .B(_02349_),
    .Y(_02351_));
 sky130_fd_sc_hd__inv_2 _15220_ (.A(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__o21ai_2 _15221_ (.A1(_02312_),
    .A2(_02334_),
    .B1(_02331_),
    .Y(_02353_));
 sky130_fd_sc_hd__xnor2_1 _15222_ (.A(_02351_),
    .B(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__nor2_1 _15223_ (.A(net563),
    .B(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__and3_1 _15224_ (.A(\core.fetchProgramCounter[6] ),
    .B(\core.fetchProgramCounter[5] ),
    .C(_02315_),
    .X(_02356_));
 sky130_fd_sc_hd__a21oi_1 _15225_ (.A1(\core.fetchProgramCounter[5] ),
    .A2(_02315_),
    .B1(\core.fetchProgramCounter[6] ),
    .Y(_02357_));
 sky130_fd_sc_hd__or2_1 _15226_ (.A(_02356_),
    .B(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__a2bb2o_1 _15227_ (.A1_N(\core.csr.trapReturnVector[6] ),
    .A2_N(net1127),
    .B1(net567),
    .B2(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__nor2_2 _15228_ (.A(\core.csr.traps.mtvec.csrReadData[6] ),
    .B(\core.csr.traps.mcause.csrReadData[4] ),
    .Y(_02360_));
 sky130_fd_sc_hd__nand2_2 _15229_ (.A(\core.csr.traps.mtvec.csrReadData[6] ),
    .B(\core.csr.traps.mcause.csrReadData[4] ),
    .Y(_02361_));
 sky130_fd_sc_hd__and2b_1 _15230_ (.A_N(_02360_),
    .B(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__a21o_1 _15231_ (.A1(\core.csr.traps.mtvec.csrReadData[5] ),
    .A2(\core.csr.traps.mcause.csrReadData[3] ),
    .B1(_02336_),
    .X(_02363_));
 sky130_fd_sc_hd__o21ai_4 _15232_ (.A1(\core.csr.traps.mtvec.csrReadData[5] ),
    .A2(\core.csr.traps.mcause.csrReadData[3] ),
    .B1(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__xnor2_1 _15233_ (.A(_02362_),
    .B(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__mux2_1 _15234_ (.A0(\core.csr.traps.mtvec.csrReadData[6] ),
    .A1(_02365_),
    .S(net1057),
    .X(_02366_));
 sky130_fd_sc_hd__a21o_1 _15235_ (.A1(net547),
    .A2(_02366_),
    .B1(net538),
    .X(_02367_));
 sky130_fd_sc_hd__nor3_1 _15236_ (.A(net546),
    .B(_02355_),
    .C(_02359_),
    .Y(_02368_));
 sky130_fd_sc_hd__o221a_1 _15237_ (.A1(\core.fetchProgramCounter[6] ),
    .A2(net524),
    .B1(_02367_),
    .B2(_02368_),
    .C1(net1830),
    .X(_00810_));
 sky130_fd_sc_hd__and2_1 _15238_ (.A(_04423_),
    .B(_07051_),
    .X(_02369_));
 sky130_fd_sc_hd__a31oi_4 _15239_ (.A1(net1182),
    .A2(_07817_),
    .A3(net571),
    .B1(_02369_),
    .Y(_02370_));
 sky130_fd_sc_hd__o22a_4 _15240_ (.A1(_03826_),
    .A2(net566),
    .B1(_02370_),
    .B2(net1229),
    .X(_02371_));
 sky130_fd_sc_hd__a21o_2 _15241_ (.A1(_07053_),
    .A2(net572),
    .B1(_03832_),
    .X(_02372_));
 sky130_fd_sc_hd__o221a_1 _15242_ (.A1(_03826_),
    .A2(net566),
    .B1(_02370_),
    .B2(net1229),
    .C1(_02372_),
    .X(_02373_));
 sky130_fd_sc_hd__xor2_4 _15243_ (.A(_02371_),
    .B(_02372_),
    .X(_02374_));
 sky130_fd_sc_hd__o21ai_1 _15244_ (.A1(_02352_),
    .A2(_02353_),
    .B1(_02350_),
    .Y(_02375_));
 sky130_fd_sc_hd__and2_1 _15245_ (.A(\core.fetchProgramCounter[7] ),
    .B(_02356_),
    .X(_02376_));
 sky130_fd_sc_hd__o21ai_1 _15246_ (.A1(\core.fetchProgramCounter[7] ),
    .A2(_02356_),
    .B1(net563),
    .Y(_02377_));
 sky130_fd_sc_hd__nor2_1 _15247_ (.A(_02376_),
    .B(_02377_),
    .Y(_02378_));
 sky130_fd_sc_hd__xnor2_1 _15248_ (.A(_02374_),
    .B(_02375_),
    .Y(_02379_));
 sky130_fd_sc_hd__a21oi_2 _15249_ (.A1(net1300),
    .A2(_02379_),
    .B1(net562),
    .Y(_02380_));
 sky130_fd_sc_hd__or3_1 _15250_ (.A(net1131),
    .B(_02378_),
    .C(_02380_),
    .X(_02381_));
 sky130_fd_sc_hd__o211a_1 _15251_ (.A1(\core.csr.trapReturnVector[7] ),
    .A2(net1127),
    .B1(net556),
    .C1(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__xnor2_1 _15252_ (.A(\core.csr.traps.mtvec.csrReadData[7] ),
    .B(\core.csr.traps.mcause.csrReadData[5] ),
    .Y(_02383_));
 sky130_fd_sc_hd__o21ai_4 _15253_ (.A1(_02360_),
    .A2(_02364_),
    .B1(_02361_),
    .Y(_02384_));
 sky130_fd_sc_hd__xnor2_1 _15254_ (.A(_02383_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__mux2_1 _15255_ (.A0(\core.csr.traps.mtvec.csrReadData[7] ),
    .A1(_02385_),
    .S(net1057),
    .X(_02386_));
 sky130_fd_sc_hd__a21o_1 _15256_ (.A1(net547),
    .A2(_02386_),
    .B1(net538),
    .X(_02387_));
 sky130_fd_sc_hd__o221a_1 _15257_ (.A1(\core.fetchProgramCounter[7] ),
    .A2(net523),
    .B1(_02382_),
    .B2(_02387_),
    .C1(net1831),
    .X(_00811_));
 sky130_fd_sc_hd__nand2_2 _15258_ (.A(\core.pipe0_currentInstruction[28] ),
    .B(net568),
    .Y(_02388_));
 sky130_fd_sc_hd__nor2_1 _15259_ (.A(_04387_),
    .B(net1181),
    .Y(_02389_));
 sky130_fd_sc_hd__a31o_1 _15260_ (.A1(net1182),
    .A2(_07855_),
    .A3(net571),
    .B1(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__a2bb2o_2 _15261_ (.A1_N(net480),
    .A2_N(_02268_),
    .B1(_02390_),
    .B2(net1225),
    .X(_02391_));
 sky130_fd_sc_hd__xor2_2 _15262_ (.A(_02388_),
    .B(_02391_),
    .X(_02392_));
 sky130_fd_sc_hd__and4bb_1 _15263_ (.A_N(_02311_),
    .B_N(_02332_),
    .C(_02351_),
    .D(_02374_),
    .X(_02393_));
 sky130_fd_sc_hd__o32ai_4 _15264_ (.A1(_03832_),
    .A2(net562),
    .A3(_02371_),
    .B1(_02373_),
    .B2(_02350_),
    .Y(_02394_));
 sky130_fd_sc_hd__a41o_1 _15265_ (.A1(_02331_),
    .A2(_02334_),
    .A3(_02351_),
    .A4(_02374_),
    .B1(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__a31o_4 _15266_ (.A1(_02289_),
    .A2(_02293_),
    .A3(_02393_),
    .B1(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__or2_1 _15267_ (.A(_02392_),
    .B(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__nand2_1 _15268_ (.A(_02392_),
    .B(_02396_),
    .Y(_02398_));
 sky130_fd_sc_hd__a21o_1 _15269_ (.A1(_02397_),
    .A2(_02398_),
    .B1(net562),
    .X(_02399_));
 sky130_fd_sc_hd__and3_2 _15270_ (.A(\core.fetchProgramCounter[8] ),
    .B(\core.fetchProgramCounter[7] ),
    .C(_02356_),
    .X(_02400_));
 sky130_fd_sc_hd__nor2_1 _15271_ (.A(\core.fetchProgramCounter[8] ),
    .B(_02376_),
    .Y(_02401_));
 sky130_fd_sc_hd__or2_1 _15272_ (.A(_02400_),
    .B(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__o2bb2a_1 _15273_ (.A1_N(net567),
    .A2_N(_02402_),
    .B1(\core.csr.trapReturnVector[8] ),
    .B2(net1127),
    .X(_02403_));
 sky130_fd_sc_hd__and3_1 _15274_ (.A(net553),
    .B(_02399_),
    .C(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__nor2_2 _15275_ (.A(\core.csr.traps.mtvec.csrReadData[8] ),
    .B(\core.csr.traps.mcause.csrReadData[6] ),
    .Y(_02405_));
 sky130_fd_sc_hd__nand2_2 _15276_ (.A(\core.csr.traps.mtvec.csrReadData[8] ),
    .B(\core.csr.traps.mcause.csrReadData[6] ),
    .Y(_02406_));
 sky130_fd_sc_hd__nand2b_1 _15277_ (.A_N(_02405_),
    .B(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__a21o_1 _15278_ (.A1(\core.csr.traps.mtvec.csrReadData[7] ),
    .A2(\core.csr.traps.mcause.csrReadData[5] ),
    .B1(_02384_),
    .X(_02408_));
 sky130_fd_sc_hd__o21ai_4 _15279_ (.A1(\core.csr.traps.mtvec.csrReadData[7] ),
    .A2(\core.csr.traps.mcause.csrReadData[5] ),
    .B1(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__xor2_1 _15280_ (.A(_02407_),
    .B(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__mux2_1 _15281_ (.A0(\core.csr.traps.mtvec.csrReadData[8] ),
    .A1(_02410_),
    .S(net1057),
    .X(_02411_));
 sky130_fd_sc_hd__a211o_1 _15282_ (.A1(net547),
    .A2(_02411_),
    .B1(_02404_),
    .C1(net538),
    .X(_02412_));
 sky130_fd_sc_hd__o211a_1 _15283_ (.A1(\core.fetchProgramCounter[8] ),
    .A2(net523),
    .B1(_02412_),
    .C1(net1831),
    .X(_00812_));
 sky130_fd_sc_hd__and2_1 _15284_ (.A(_04301_),
    .B(_07051_),
    .X(_02413_));
 sky130_fd_sc_hd__a31o_1 _15285_ (.A1(net1182),
    .A2(_07896_),
    .A3(net571),
    .B1(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__o2bb2a_2 _15286_ (.A1_N(net1225),
    .A2_N(_02414_),
    .B1(net566),
    .B2(_03825_),
    .X(_02415_));
 sky130_fd_sc_hd__nand2_1 _15287_ (.A(\core.pipe0_currentInstruction[29] ),
    .B(net568),
    .Y(_02416_));
 sky130_fd_sc_hd__nand2_1 _15288_ (.A(_02415_),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__or2_1 _15289_ (.A(_02415_),
    .B(_02416_),
    .X(_02418_));
 sky130_fd_sc_hd__and2_1 _15290_ (.A(_02417_),
    .B(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__o21a_1 _15291_ (.A1(_02388_),
    .A2(_02391_),
    .B1(_02398_),
    .X(_02420_));
 sky130_fd_sc_hd__xor2_1 _15292_ (.A(\core.fetchProgramCounter[9] ),
    .B(_02400_),
    .X(_02421_));
 sky130_fd_sc_hd__xor2_1 _15293_ (.A(_02419_),
    .B(_02420_),
    .X(_02422_));
 sky130_fd_sc_hd__a21oi_2 _15294_ (.A1(net1300),
    .A2(_02422_),
    .B1(net562),
    .Y(_02423_));
 sky130_fd_sc_hd__a211o_1 _15295_ (.A1(net562),
    .A2(_02421_),
    .B1(_02423_),
    .C1(net1131),
    .X(_02424_));
 sky130_fd_sc_hd__o211a_1 _15296_ (.A1(\core.csr.trapReturnVector[9] ),
    .A2(net1127),
    .B1(net553),
    .C1(_02424_),
    .X(_02425_));
 sky130_fd_sc_hd__xnor2_1 _15297_ (.A(\core.csr.traps.mtvec.csrReadData[9] ),
    .B(\core.csr.traps.mcause.csrReadData[7] ),
    .Y(_02426_));
 sky130_fd_sc_hd__o21ai_4 _15298_ (.A1(_02405_),
    .A2(_02409_),
    .B1(_02406_),
    .Y(_02427_));
 sky130_fd_sc_hd__xnor2_1 _15299_ (.A(_02426_),
    .B(_02427_),
    .Y(_02428_));
 sky130_fd_sc_hd__mux2_1 _15300_ (.A0(\core.csr.traps.mtvec.csrReadData[9] ),
    .A1(_02428_),
    .S(net1058),
    .X(_02429_));
 sky130_fd_sc_hd__a21o_1 _15301_ (.A1(net545),
    .A2(_02429_),
    .B1(net538),
    .X(_02430_));
 sky130_fd_sc_hd__o221a_1 _15302_ (.A1(\core.fetchProgramCounter[9] ),
    .A2(net523),
    .B1(_02425_),
    .B2(_02430_),
    .C1(net1827),
    .X(_00813_));
 sky130_fd_sc_hd__and2_1 _15303_ (.A(_04213_),
    .B(_07051_),
    .X(_02431_));
 sky130_fd_sc_hd__a31o_1 _15304_ (.A1(net1182),
    .A2(_07928_),
    .A3(net572),
    .B1(_02431_),
    .X(_02432_));
 sky130_fd_sc_hd__a22o_1 _15305_ (.A1(net451),
    .A2(_02269_),
    .B1(_02432_),
    .B2(net1225),
    .X(_02433_));
 sky130_fd_sc_hd__a21oi_1 _15306_ (.A1(net1752),
    .A2(_02249_),
    .B1(_02433_),
    .Y(_02434_));
 sky130_fd_sc_hd__or3b_4 _15307_ (.A(_03831_),
    .B(net562),
    .C_N(_02433_),
    .X(_02435_));
 sky130_fd_sc_hd__and2b_1 _15308_ (.A_N(_02434_),
    .B(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__a21o_1 _15309_ (.A1(_02415_),
    .A2(_02416_),
    .B1(_02420_),
    .X(_02437_));
 sky130_fd_sc_hd__nand2_1 _15310_ (.A(_02418_),
    .B(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__or2_1 _15311_ (.A(_02436_),
    .B(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__nand2_1 _15312_ (.A(_02436_),
    .B(_02438_),
    .Y(_02440_));
 sky130_fd_sc_hd__nand2_1 _15313_ (.A(_02439_),
    .B(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__and3_1 _15314_ (.A(\core.fetchProgramCounter[10] ),
    .B(\core.fetchProgramCounter[9] ),
    .C(_02400_),
    .X(_02442_));
 sky130_fd_sc_hd__a21oi_1 _15315_ (.A1(\core.fetchProgramCounter[9] ),
    .A2(_02400_),
    .B1(\core.fetchProgramCounter[10] ),
    .Y(_02443_));
 sky130_fd_sc_hd__o21ai_1 _15316_ (.A1(_02442_),
    .A2(_02443_),
    .B1(net567),
    .Y(_02444_));
 sky130_fd_sc_hd__o211ai_1 _15317_ (.A1(\core.csr.trapReturnVector[10] ),
    .A2(net1127),
    .B1(net554),
    .C1(_02444_),
    .Y(_02445_));
 sky130_fd_sc_hd__a21oi_1 _15318_ (.A1(net568),
    .A2(_02441_),
    .B1(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__nor2_1 _15319_ (.A(\core.csr.traps.mtvec.csrReadData[10] ),
    .B(\core.csr.traps.mcause.csrReadData[8] ),
    .Y(_02447_));
 sky130_fd_sc_hd__nand2_1 _15320_ (.A(\core.csr.traps.mtvec.csrReadData[10] ),
    .B(\core.csr.traps.mcause.csrReadData[8] ),
    .Y(_02448_));
 sky130_fd_sc_hd__nand2b_1 _15321_ (.A_N(_02447_),
    .B(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__a21o_1 _15322_ (.A1(\core.csr.traps.mtvec.csrReadData[9] ),
    .A2(\core.csr.traps.mcause.csrReadData[7] ),
    .B1(_02427_),
    .X(_02450_));
 sky130_fd_sc_hd__o21ai_2 _15323_ (.A1(\core.csr.traps.mtvec.csrReadData[9] ),
    .A2(\core.csr.traps.mcause.csrReadData[7] ),
    .B1(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__xor2_1 _15324_ (.A(_02449_),
    .B(_02451_),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _15325_ (.A0(\core.csr.traps.mtvec.csrReadData[10] ),
    .A1(_02452_),
    .S(net1057),
    .X(_02453_));
 sky130_fd_sc_hd__a21o_1 _15326_ (.A1(net545),
    .A2(_02453_),
    .B1(net538),
    .X(_02454_));
 sky130_fd_sc_hd__o221a_1 _15327_ (.A1(\core.fetchProgramCounter[10] ),
    .A2(net523),
    .B1(_02446_),
    .B2(_02454_),
    .C1(net1827),
    .X(_00814_));
 sky130_fd_sc_hd__and3_1 _15328_ (.A(\core.pipe0_currentInstruction[7] ),
    .B(_06998_),
    .C(_08700_),
    .X(_02455_));
 sky130_fd_sc_hd__nor2_2 _15329_ (.A(net1751),
    .B(_07048_),
    .Y(_02456_));
 sky130_fd_sc_hd__nor2_1 _15330_ (.A(net1136),
    .B(_02456_),
    .Y(_02457_));
 sky130_fd_sc_hd__o22a_1 _15331_ (.A1(net1776),
    .A2(net1225),
    .B1(_02455_),
    .B2(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__and2_1 _15332_ (.A(_04044_),
    .B(net1185),
    .X(_02459_));
 sky130_fd_sc_hd__a31o_1 _15333_ (.A1(net1183),
    .A2(_07964_),
    .A3(net572),
    .B1(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__a22oi_2 _15334_ (.A1(net452),
    .A2(_02269_),
    .B1(_02460_),
    .B2(net1225),
    .Y(_02461_));
 sky130_fd_sc_hd__and2b_1 _15335_ (.A_N(_02458_),
    .B(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__nand2b_2 _15336_ (.A_N(_02461_),
    .B(_02458_),
    .Y(_02463_));
 sky130_fd_sc_hd__and2b_1 _15337_ (.A_N(_02462_),
    .B(_02463_),
    .X(_02464_));
 sky130_fd_sc_hd__a21oi_1 _15338_ (.A1(_02435_),
    .A2(_02440_),
    .B1(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__a31o_1 _15339_ (.A1(_02435_),
    .A2(_02440_),
    .A3(_02464_),
    .B1(net562),
    .X(_02466_));
 sky130_fd_sc_hd__nor2_2 _15340_ (.A(_02465_),
    .B(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__and2_2 _15341_ (.A(\core.fetchProgramCounter[11] ),
    .B(_02442_),
    .X(_02468_));
 sky130_fd_sc_hd__nor2_1 _15342_ (.A(\core.fetchProgramCounter[11] ),
    .B(_02442_),
    .Y(_02469_));
 sky130_fd_sc_hd__o21ai_1 _15343_ (.A1(_02468_),
    .A2(_02469_),
    .B1(_02260_),
    .Y(_02470_));
 sky130_fd_sc_hd__o211ai_1 _15344_ (.A1(\core.csr.trapReturnVector[11] ),
    .A2(net1127),
    .B1(net554),
    .C1(_02470_),
    .Y(_02471_));
 sky130_fd_sc_hd__xnor2_1 _15345_ (.A(\core.csr.traps.mtvec.csrReadData[11] ),
    .B(\core.csr.traps.mcause.csrReadData[9] ),
    .Y(_02472_));
 sky130_fd_sc_hd__o21ai_2 _15346_ (.A1(_02447_),
    .A2(_02451_),
    .B1(_02448_),
    .Y(_02473_));
 sky130_fd_sc_hd__xnor2_1 _15347_ (.A(_02472_),
    .B(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__mux2_1 _15348_ (.A0(\core.csr.traps.mtvec.csrReadData[11] ),
    .A1(_02474_),
    .S(net1058),
    .X(_02475_));
 sky130_fd_sc_hd__a21oi_1 _15349_ (.A1(net545),
    .A2(_02475_),
    .B1(net538),
    .Y(_02476_));
 sky130_fd_sc_hd__o21ai_1 _15350_ (.A1(_02467_),
    .A2(_02471_),
    .B1(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__o211a_1 _15351_ (.A1(\core.fetchProgramCounter[11] ),
    .A2(net523),
    .B1(_02477_),
    .C1(net1827),
    .X(_00815_));
 sky130_fd_sc_hd__nand2_1 _15352_ (.A(\core.fetchProgramCounter[12] ),
    .B(_02468_),
    .Y(_02478_));
 sky130_fd_sc_hd__or2_1 _15353_ (.A(\core.fetchProgramCounter[12] ),
    .B(_02468_),
    .X(_02479_));
 sky130_fd_sc_hd__a31o_1 _15354_ (.A1(net563),
    .A2(_02478_),
    .A3(_02479_),
    .B1(net1131),
    .X(_02480_));
 sky130_fd_sc_hd__a21oi_4 _15355_ (.A1(net1136),
    .A2(net572),
    .B1(_02456_),
    .Y(_02481_));
 sky130_fd_sc_hd__o21a_1 _15356_ (.A1(\core.pipe0_currentInstruction[12] ),
    .A2(net1224),
    .B1(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__nor2_1 _15357_ (.A(_06506_),
    .B(net1183),
    .Y(_02483_));
 sky130_fd_sc_hd__a31o_1 _15358_ (.A1(net1183),
    .A2(_08017_),
    .A3(net572),
    .B1(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__a2bb2o_2 _15359_ (.A1_N(net453),
    .A2_N(_02268_),
    .B1(_02484_),
    .B2(net1224),
    .X(_02485_));
 sky130_fd_sc_hd__a2111o_1 _15360_ (.A1(_03843_),
    .A2(net1229),
    .B1(net564),
    .C1(_02456_),
    .D1(_02485_),
    .X(_02486_));
 sky130_fd_sc_hd__xor2_2 _15361_ (.A(_02482_),
    .B(_02485_),
    .X(_02487_));
 sky130_fd_sc_hd__a211o_1 _15362_ (.A1(_02415_),
    .A2(_02416_),
    .B1(_02388_),
    .C1(_02391_),
    .X(_02488_));
 sky130_fd_sc_hd__a311o_2 _15363_ (.A1(_02418_),
    .A2(_02435_),
    .A3(_02488_),
    .B1(_02462_),
    .C1(_02434_),
    .X(_02489_));
 sky130_fd_sc_hd__nand2_1 _15364_ (.A(_02463_),
    .B(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__and4_2 _15365_ (.A(_02392_),
    .B(_02419_),
    .C(_02436_),
    .D(_02464_),
    .X(_02491_));
 sky130_fd_sc_hd__a21oi_1 _15366_ (.A1(_02396_),
    .A2(_02491_),
    .B1(_02490_),
    .Y(_02492_));
 sky130_fd_sc_hd__or2_1 _15367_ (.A(_02487_),
    .B(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__nand2_1 _15368_ (.A(_02487_),
    .B(_02492_),
    .Y(_02494_));
 sky130_fd_sc_hd__and3_1 _15369_ (.A(net568),
    .B(_02493_),
    .C(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__o221a_1 _15370_ (.A1(\core.csr.trapReturnVector[12] ),
    .A2(net1129),
    .B1(_02480_),
    .B2(_02495_),
    .C1(net553),
    .X(_02496_));
 sky130_fd_sc_hd__nand2_2 _15371_ (.A(\core.csr.traps.mtvec.csrReadData[12] ),
    .B(\core.csr.traps.mcause.csrReadData[10] ),
    .Y(_02497_));
 sky130_fd_sc_hd__or2_1 _15372_ (.A(\core.csr.traps.mtvec.csrReadData[12] ),
    .B(\core.csr.traps.mcause.csrReadData[10] ),
    .X(_02498_));
 sky130_fd_sc_hd__nand2_2 _15373_ (.A(_02497_),
    .B(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__a21o_1 _15374_ (.A1(\core.csr.traps.mtvec.csrReadData[11] ),
    .A2(\core.csr.traps.mcause.csrReadData[9] ),
    .B1(_02473_),
    .X(_02500_));
 sky130_fd_sc_hd__o21ai_4 _15375_ (.A1(\core.csr.traps.mtvec.csrReadData[11] ),
    .A2(\core.csr.traps.mcause.csrReadData[9] ),
    .B1(_02500_),
    .Y(_02501_));
 sky130_fd_sc_hd__xor2_1 _15376_ (.A(_02499_),
    .B(_02501_),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _15377_ (.A0(\core.csr.traps.mtvec.csrReadData[12] ),
    .A1(_02502_),
    .S(net1058),
    .X(_02503_));
 sky130_fd_sc_hd__a21o_1 _15378_ (.A1(net547),
    .A2(_02503_),
    .B1(net539),
    .X(_02504_));
 sky130_fd_sc_hd__o221a_1 _15379_ (.A1(\core.fetchProgramCounter[12] ),
    .A2(net524),
    .B1(_02496_),
    .B2(_02504_),
    .C1(net1827),
    .X(_00816_));
 sky130_fd_sc_hd__and2_1 _15380_ (.A(_06428_),
    .B(net1185),
    .X(_02505_));
 sky130_fd_sc_hd__a31o_1 _15381_ (.A1(net1183),
    .A2(_08052_),
    .A3(net572),
    .B1(_02505_),
    .X(_02506_));
 sky130_fd_sc_hd__a22o_1 _15382_ (.A1(net454),
    .A2(_02269_),
    .B1(_02506_),
    .B2(net1225),
    .X(_02507_));
 sky130_fd_sc_hd__o21a_1 _15383_ (.A1(\core.pipe0_currentInstruction[13] ),
    .A2(net1224),
    .B1(_02481_),
    .X(_02508_));
 sky130_fd_sc_hd__nor2_1 _15384_ (.A(_02507_),
    .B(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__and2_1 _15385_ (.A(_02486_),
    .B(_02493_),
    .X(_02510_));
 sky130_fd_sc_hd__nand2_1 _15386_ (.A(_02507_),
    .B(_02508_),
    .Y(_02511_));
 sky130_fd_sc_hd__xnor2_1 _15387_ (.A(_02507_),
    .B(_02508_),
    .Y(_02512_));
 sky130_fd_sc_hd__and3_1 _15388_ (.A(\core.fetchProgramCounter[13] ),
    .B(\core.fetchProgramCounter[12] ),
    .C(_02468_),
    .X(_02513_));
 sky130_fd_sc_hd__a21oi_1 _15389_ (.A1(\core.fetchProgramCounter[12] ),
    .A2(_02468_),
    .B1(\core.fetchProgramCounter[13] ),
    .Y(_02514_));
 sky130_fd_sc_hd__nor2_1 _15390_ (.A(_02513_),
    .B(_02514_),
    .Y(_02515_));
 sky130_fd_sc_hd__xnor2_1 _15391_ (.A(_02510_),
    .B(_02512_),
    .Y(_02516_));
 sky130_fd_sc_hd__a21oi_2 _15392_ (.A1(net1300),
    .A2(_02516_),
    .B1(net564),
    .Y(_02517_));
 sky130_fd_sc_hd__a211o_1 _15393_ (.A1(net563),
    .A2(_02515_),
    .B1(_02517_),
    .C1(net1131),
    .X(_02518_));
 sky130_fd_sc_hd__o211a_1 _15394_ (.A1(\core.csr.trapReturnVector[13] ),
    .A2(net1127),
    .B1(net553),
    .C1(_02518_),
    .X(_02519_));
 sky130_fd_sc_hd__o21ai_4 _15395_ (.A1(_02499_),
    .A2(_02501_),
    .B1(_02497_),
    .Y(_02520_));
 sky130_fd_sc_hd__nand2_1 _15396_ (.A(\core.csr.traps.mtvec.csrReadData[13] ),
    .B(\core.csr.traps.mcause.csrReadData[11] ),
    .Y(_02521_));
 sky130_fd_sc_hd__or2_1 _15397_ (.A(\core.csr.traps.mtvec.csrReadData[13] ),
    .B(\core.csr.traps.mcause.csrReadData[11] ),
    .X(_02522_));
 sky130_fd_sc_hd__nand2_1 _15398_ (.A(_02521_),
    .B(_02522_),
    .Y(_02523_));
 sky130_fd_sc_hd__xnor2_1 _15399_ (.A(_02520_),
    .B(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__mux2_2 _15400_ (.A0(\core.csr.traps.mtvec.csrReadData[13] ),
    .A1(_02524_),
    .S(net1057),
    .X(_02525_));
 sky130_fd_sc_hd__a21o_1 _15401_ (.A1(net545),
    .A2(_02525_),
    .B1(net539),
    .X(_02526_));
 sky130_fd_sc_hd__o221a_1 _15402_ (.A1(\core.fetchProgramCounter[13] ),
    .A2(net524),
    .B1(_02519_),
    .B2(_02526_),
    .C1(net1827),
    .X(_00817_));
 sky130_fd_sc_hd__o21ai_4 _15403_ (.A1(net1795),
    .A2(net1224),
    .B1(_02481_),
    .Y(_02527_));
 sky130_fd_sc_hd__nor2_1 _15404_ (.A(_06353_),
    .B(net1183),
    .Y(_02528_));
 sky130_fd_sc_hd__a31o_1 _15405_ (.A1(net1183),
    .A2(_08087_),
    .A3(net570),
    .B1(_02528_),
    .X(_02529_));
 sky130_fd_sc_hd__a2bb2o_2 _15406_ (.A1_N(net455),
    .A2_N(net566),
    .B1(_02529_),
    .B2(net1224),
    .X(_02530_));
 sky130_fd_sc_hd__or2_2 _15407_ (.A(_02527_),
    .B(_02530_),
    .X(_02531_));
 sky130_fd_sc_hd__xnor2_4 _15408_ (.A(_02527_),
    .B(_02530_),
    .Y(_02532_));
 sky130_fd_sc_hd__a31o_1 _15409_ (.A1(_02486_),
    .A2(_02493_),
    .A3(_02511_),
    .B1(_02509_),
    .X(_02533_));
 sky130_fd_sc_hd__xnor2_1 _15410_ (.A(_02532_),
    .B(_02533_),
    .Y(_02534_));
 sky130_fd_sc_hd__or2_1 _15411_ (.A(\core.csr.trapReturnVector[14] ),
    .B(net1127),
    .X(_02535_));
 sky130_fd_sc_hd__and2_2 _15412_ (.A(\core.fetchProgramCounter[14] ),
    .B(_02513_),
    .X(_02536_));
 sky130_fd_sc_hd__o21ai_1 _15413_ (.A1(\core.fetchProgramCounter[14] ),
    .A2(_02513_),
    .B1(net564),
    .Y(_02537_));
 sky130_fd_sc_hd__nor2_1 _15414_ (.A(_02536_),
    .B(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__a21oi_2 _15415_ (.A1(net1299),
    .A2(_02534_),
    .B1(net564),
    .Y(_02539_));
 sky130_fd_sc_hd__or3_1 _15416_ (.A(net1131),
    .B(_02538_),
    .C(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__nand2_1 _15417_ (.A(\core.csr.traps.mtvec.csrReadData[14] ),
    .B(\core.csr.traps.mcause.csrReadData[12] ),
    .Y(_02541_));
 sky130_fd_sc_hd__or2_1 _15418_ (.A(\core.csr.traps.mtvec.csrReadData[14] ),
    .B(\core.csr.traps.mcause.csrReadData[12] ),
    .X(_02542_));
 sky130_fd_sc_hd__nand2_1 _15419_ (.A(_02541_),
    .B(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__a21boi_2 _15420_ (.A1(_02520_),
    .A2(_02522_),
    .B1_N(_02521_),
    .Y(_02544_));
 sky130_fd_sc_hd__xnor2_1 _15421_ (.A(_02543_),
    .B(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__nand2_1 _15422_ (.A(net1058),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__o211a_1 _15423_ (.A1(\core.csr.traps.mtvec.csrReadData[14] ),
    .A2(net1058),
    .B1(_02546_),
    .C1(net548),
    .X(_02547_));
 sky130_fd_sc_hd__a311o_1 _15424_ (.A1(net554),
    .A2(_02535_),
    .A3(_02540_),
    .B1(_02547_),
    .C1(net538),
    .X(_02548_));
 sky130_fd_sc_hd__o211a_1 _15425_ (.A1(\core.fetchProgramCounter[14] ),
    .A2(net524),
    .B1(_02548_),
    .C1(net1827),
    .X(_00818_));
 sky130_fd_sc_hd__and2_1 _15426_ (.A(_06277_),
    .B(net1185),
    .X(_02549_));
 sky130_fd_sc_hd__a31o_1 _15427_ (.A1(net1183),
    .A2(_08095_),
    .A3(net570),
    .B1(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__a22o_2 _15428_ (.A1(net456),
    .A2(_02269_),
    .B1(_02550_),
    .B2(net1224),
    .X(_02551_));
 sky130_fd_sc_hd__o21a_2 _15429_ (.A1(net1793),
    .A2(net1224),
    .B1(_02481_),
    .X(_02552_));
 sky130_fd_sc_hd__nor2_1 _15430_ (.A(_02551_),
    .B(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__nand2_1 _15431_ (.A(_02551_),
    .B(_02552_),
    .Y(_02554_));
 sky130_fd_sc_hd__xnor2_2 _15432_ (.A(_02551_),
    .B(_02552_),
    .Y(_02555_));
 sky130_fd_sc_hd__o21ai_1 _15433_ (.A1(_02532_),
    .A2(_02533_),
    .B1(_02531_),
    .Y(_02556_));
 sky130_fd_sc_hd__o21ai_1 _15434_ (.A1(\core.fetchProgramCounter[15] ),
    .A2(_02536_),
    .B1(net564),
    .Y(_02557_));
 sky130_fd_sc_hd__a21o_1 _15435_ (.A1(\core.fetchProgramCounter[15] ),
    .A2(_02536_),
    .B1(_02557_),
    .X(_02558_));
 sky130_fd_sc_hd__xor2_1 _15436_ (.A(_02555_),
    .B(_02556_),
    .X(_02559_));
 sky130_fd_sc_hd__a21o_1 _15437_ (.A1(net1300),
    .A2(_02559_),
    .B1(net564),
    .X(_02560_));
 sky130_fd_sc_hd__o21ai_1 _15438_ (.A1(\core.csr.trapReturnVector[15] ),
    .A2(net1129),
    .B1(net553),
    .Y(_02561_));
 sky130_fd_sc_hd__a31o_1 _15439_ (.A1(net1129),
    .A2(_02558_),
    .A3(_02560_),
    .B1(_02561_),
    .X(_02562_));
 sky130_fd_sc_hd__nor2_1 _15440_ (.A(\core.csr.traps.mtvec.csrReadData[15] ),
    .B(net1058),
    .Y(_02563_));
 sky130_fd_sc_hd__o21a_2 _15441_ (.A1(_02543_),
    .A2(_02544_),
    .B1(_02541_),
    .X(_02564_));
 sky130_fd_sc_hd__nand2_1 _15442_ (.A(\core.csr.traps.mtvec.csrReadData[15] ),
    .B(\core.csr.traps.mcause.csrReadData[13] ),
    .Y(_02565_));
 sky130_fd_sc_hd__or2_1 _15443_ (.A(\core.csr.traps.mtvec.csrReadData[15] ),
    .B(\core.csr.traps.mcause.csrReadData[13] ),
    .X(_02566_));
 sky130_fd_sc_hd__nand2_1 _15444_ (.A(_02565_),
    .B(_02566_),
    .Y(_02567_));
 sky130_fd_sc_hd__xnor2_1 _15445_ (.A(_02564_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__a211o_1 _15446_ (.A1(net1058),
    .A2(_02568_),
    .B1(_02563_),
    .C1(net553),
    .X(_02569_));
 sky130_fd_sc_hd__nor2_1 _15447_ (.A(\core.fetchProgramCounter[15] ),
    .B(net524),
    .Y(_02570_));
 sky130_fd_sc_hd__a311oi_1 _15448_ (.A1(net524),
    .A2(_02562_),
    .A3(_02569_),
    .B1(_02570_),
    .C1(net1876),
    .Y(_00819_));
 sky130_fd_sc_hd__o21a_1 _15449_ (.A1(net1789),
    .A2(net1222),
    .B1(_02481_),
    .X(_02571_));
 sky130_fd_sc_hd__nor2_1 _15450_ (.A(_06198_),
    .B(net1180),
    .Y(_02572_));
 sky130_fd_sc_hd__a31o_1 _15451_ (.A1(net1180),
    .A2(_08159_),
    .A3(net570),
    .B1(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__nand2_1 _15452_ (.A(net1222),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__o21a_1 _15453_ (.A1(net1747),
    .A2(net566),
    .B1(_02574_),
    .X(_02575_));
 sky130_fd_sc_hd__o211a_1 _15454_ (.A1(net1747),
    .A2(net566),
    .B1(_02571_),
    .C1(_02574_),
    .X(_02576_));
 sky130_fd_sc_hd__xnor2_2 _15455_ (.A(_02571_),
    .B(_02575_),
    .Y(_02577_));
 sky130_fd_sc_hd__or4_2 _15456_ (.A(_02487_),
    .B(_02512_),
    .C(_02532_),
    .D(_02555_),
    .X(_02578_));
 sky130_fd_sc_hd__inv_2 _15457_ (.A(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__a21oi_2 _15458_ (.A1(_02463_),
    .A2(_02489_),
    .B1(_02578_),
    .Y(_02580_));
 sky130_fd_sc_hd__a2111o_2 _15459_ (.A1(_02486_),
    .A2(_02511_),
    .B1(_02532_),
    .C1(_02555_),
    .D1(_02509_),
    .X(_02581_));
 sky130_fd_sc_hd__o211ai_4 _15460_ (.A1(_02531_),
    .A2(_02553_),
    .B1(_02554_),
    .C1(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__a311oi_4 _15461_ (.A1(_02396_),
    .A2(_02491_),
    .A3(_02579_),
    .B1(_02580_),
    .C1(_02582_),
    .Y(_02583_));
 sky130_fd_sc_hd__and2_1 _15462_ (.A(_02577_),
    .B(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__nor2_1 _15463_ (.A(_02577_),
    .B(_02583_),
    .Y(_02585_));
 sky130_fd_sc_hd__or2_1 _15464_ (.A(_02584_),
    .B(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__and3_2 _15465_ (.A(\core.fetchProgramCounter[16] ),
    .B(\core.fetchProgramCounter[15] ),
    .C(_02536_),
    .X(_02587_));
 sky130_fd_sc_hd__a21oi_1 _15466_ (.A1(\core.fetchProgramCounter[15] ),
    .A2(_02536_),
    .B1(\core.fetchProgramCounter[16] ),
    .Y(_02588_));
 sky130_fd_sc_hd__or2_1 _15467_ (.A(_02587_),
    .B(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__a2bb2o_1 _15468_ (.A1_N(\core.csr.trapReturnVector[16] ),
    .A2_N(net1129),
    .B1(net567),
    .B2(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__a211oi_1 _15469_ (.A1(net568),
    .A2(_02586_),
    .B1(_02590_),
    .C1(net543),
    .Y(_02591_));
 sky130_fd_sc_hd__nand2_1 _15470_ (.A(\core.csr.traps.mtvec.csrReadData[16] ),
    .B(\core.csr.traps.mcause.csrReadData[14] ),
    .Y(_02592_));
 sky130_fd_sc_hd__or2_1 _15471_ (.A(\core.csr.traps.mtvec.csrReadData[16] ),
    .B(\core.csr.traps.mcause.csrReadData[14] ),
    .X(_02593_));
 sky130_fd_sc_hd__nand2_1 _15472_ (.A(_02592_),
    .B(_02593_),
    .Y(_02594_));
 sky130_fd_sc_hd__o21ai_2 _15473_ (.A1(_02564_),
    .A2(_02567_),
    .B1(_02565_),
    .Y(_02595_));
 sky130_fd_sc_hd__xnor2_1 _15474_ (.A(_02594_),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__mux2_1 _15475_ (.A0(\core.csr.traps.mtvec.csrReadData[16] ),
    .A1(_02596_),
    .S(net1058),
    .X(_02597_));
 sky130_fd_sc_hd__a21o_1 _15476_ (.A1(net548),
    .A2(_02597_),
    .B1(net539),
    .X(_02598_));
 sky130_fd_sc_hd__o221a_1 _15477_ (.A1(\core.fetchProgramCounter[16] ),
    .A2(net524),
    .B1(_02591_),
    .B2(_02598_),
    .C1(net1826),
    .X(_00820_));
 sky130_fd_sc_hd__nor2_1 _15478_ (.A(_06121_),
    .B(net1180),
    .Y(_02599_));
 sky130_fd_sc_hd__a31o_1 _15479_ (.A1(net1180),
    .A2(_08167_),
    .A3(net570),
    .B1(_02599_),
    .X(_02600_));
 sky130_fd_sc_hd__a22o_2 _15480_ (.A1(net458),
    .A2(_02269_),
    .B1(_02600_),
    .B2(net1222),
    .X(_02601_));
 sky130_fd_sc_hd__nand2_2 _15481_ (.A(net1669),
    .B(net1228),
    .Y(_02602_));
 sky130_fd_sc_hd__a21oi_2 _15482_ (.A1(_02481_),
    .A2(_02602_),
    .B1(_02601_),
    .Y(_02603_));
 sky130_fd_sc_hd__a21o_1 _15483_ (.A1(_02481_),
    .A2(_02602_),
    .B1(_02601_),
    .X(_02604_));
 sky130_fd_sc_hd__nand3_2 _15484_ (.A(_02481_),
    .B(_02601_),
    .C(_02602_),
    .Y(_02605_));
 sky130_fd_sc_hd__inv_2 _15485_ (.A(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__nand2_1 _15486_ (.A(_02604_),
    .B(_02605_),
    .Y(_02607_));
 sky130_fd_sc_hd__nor2_1 _15487_ (.A(_02576_),
    .B(_02585_),
    .Y(_02608_));
 sky130_fd_sc_hd__xor2_1 _15488_ (.A(\core.fetchProgramCounter[17] ),
    .B(_02587_),
    .X(_02609_));
 sky130_fd_sc_hd__xnor2_1 _15489_ (.A(_02607_),
    .B(_02608_),
    .Y(_02610_));
 sky130_fd_sc_hd__a21oi_1 _15490_ (.A1(net1299),
    .A2(_02610_),
    .B1(net561),
    .Y(_02611_));
 sky130_fd_sc_hd__a211o_1 _15491_ (.A1(net561),
    .A2(_02609_),
    .B1(_02611_),
    .C1(net1130),
    .X(_02612_));
 sky130_fd_sc_hd__o211a_1 _15492_ (.A1(\core.csr.trapReturnVector[17] ),
    .A2(net1129),
    .B1(net554),
    .C1(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__a21bo_2 _15493_ (.A1(_02593_),
    .A2(_02595_),
    .B1_N(_02592_),
    .X(_02614_));
 sky130_fd_sc_hd__nand2_1 _15494_ (.A(\core.csr.traps.mtvec.csrReadData[17] ),
    .B(\core.csr.traps.mcause.csrReadData[15] ),
    .Y(_02615_));
 sky130_fd_sc_hd__or2_2 _15495_ (.A(\core.csr.traps.mtvec.csrReadData[17] ),
    .B(\core.csr.traps.mcause.csrReadData[15] ),
    .X(_02616_));
 sky130_fd_sc_hd__nand2_1 _15496_ (.A(_02615_),
    .B(_02616_),
    .Y(_02617_));
 sky130_fd_sc_hd__xnor2_1 _15497_ (.A(_02614_),
    .B(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__mux2_1 _15498_ (.A0(\core.csr.traps.mtvec.csrReadData[17] ),
    .A1(_02618_),
    .S(net1058),
    .X(_02619_));
 sky130_fd_sc_hd__a21o_1 _15499_ (.A1(net544),
    .A2(_02619_),
    .B1(net539),
    .X(_02620_));
 sky130_fd_sc_hd__o221a_1 _15500_ (.A1(\core.fetchProgramCounter[17] ),
    .A2(net524),
    .B1(_02613_),
    .B2(_02620_),
    .C1(net1826),
    .X(_00821_));
 sky130_fd_sc_hd__o21ai_2 _15501_ (.A1(\core.pipe0_currentInstruction[18] ),
    .A2(net1222),
    .B1(_02481_),
    .Y(_02621_));
 sky130_fd_sc_hd__nor2_1 _15502_ (.A(_06044_),
    .B(net1180),
    .Y(_02622_));
 sky130_fd_sc_hd__a31o_1 _15503_ (.A1(net1184),
    .A2(_08226_),
    .A3(net570),
    .B1(_02622_),
    .X(_02623_));
 sky130_fd_sc_hd__a2bb2o_1 _15504_ (.A1_N(net459),
    .A2_N(net566),
    .B1(_02623_),
    .B2(net1222),
    .X(_02624_));
 sky130_fd_sc_hd__nor2_1 _15505_ (.A(_02621_),
    .B(_02624_),
    .Y(_02625_));
 sky130_fd_sc_hd__xnor2_1 _15506_ (.A(_02621_),
    .B(_02624_),
    .Y(_02626_));
 sky130_fd_sc_hd__inv_2 _15507_ (.A(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__and2b_1 _15508_ (.A_N(_02576_),
    .B(_02605_),
    .X(_02628_));
 sky130_fd_sc_hd__a21oi_1 _15509_ (.A1(_02605_),
    .A2(_02608_),
    .B1(_02603_),
    .Y(_02629_));
 sky130_fd_sc_hd__o311a_1 _15510_ (.A1(_02576_),
    .A2(_02585_),
    .A3(_02606_),
    .B1(_02627_),
    .C1(_02604_),
    .X(_02630_));
 sky130_fd_sc_hd__xnor2_1 _15511_ (.A(_02627_),
    .B(_02629_),
    .Y(_02631_));
 sky130_fd_sc_hd__and3_2 _15512_ (.A(\core.fetchProgramCounter[18] ),
    .B(\core.fetchProgramCounter[17] ),
    .C(_02587_),
    .X(_02632_));
 sky130_fd_sc_hd__a21oi_1 _15513_ (.A1(\core.fetchProgramCounter[17] ),
    .A2(_02587_),
    .B1(\core.fetchProgramCounter[18] ),
    .Y(_02633_));
 sky130_fd_sc_hd__nor2_1 _15514_ (.A(_02632_),
    .B(_02633_),
    .Y(_02634_));
 sky130_fd_sc_hd__a21oi_1 _15515_ (.A1(net1299),
    .A2(_02631_),
    .B1(net561),
    .Y(_02635_));
 sky130_fd_sc_hd__a211o_1 _15516_ (.A1(net561),
    .A2(_02634_),
    .B1(_02635_),
    .C1(net1130),
    .X(_02636_));
 sky130_fd_sc_hd__o21a_1 _15517_ (.A1(\core.csr.trapReturnVector[18] ),
    .A2(net1126),
    .B1(net551),
    .X(_02637_));
 sky130_fd_sc_hd__a21boi_4 _15518_ (.A1(_02614_),
    .A2(_02616_),
    .B1_N(_02615_),
    .Y(_02638_));
 sky130_fd_sc_hd__nor2_1 _15519_ (.A(\core.csr.traps.mtvec.csrReadData[18] ),
    .B(\core.csr.traps.mcause.csrReadData[16] ),
    .Y(_02639_));
 sky130_fd_sc_hd__nand2_1 _15520_ (.A(\core.csr.traps.mtvec.csrReadData[18] ),
    .B(\core.csr.traps.mcause.csrReadData[16] ),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2b_1 _15521_ (.A_N(_02639_),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__xor2_1 _15522_ (.A(_02638_),
    .B(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__mux2_1 _15523_ (.A0(\core.csr.traps.mtvec.csrReadData[18] ),
    .A1(_02642_),
    .S(_02277_),
    .X(_02643_));
 sky130_fd_sc_hd__a221o_1 _15524_ (.A1(_02636_),
    .A2(_02637_),
    .B1(_02643_),
    .B2(net543),
    .C1(net540),
    .X(_02644_));
 sky130_fd_sc_hd__o211a_1 _15525_ (.A1(\core.fetchProgramCounter[18] ),
    .A2(net522),
    .B1(_02644_),
    .C1(net1815),
    .X(_00822_));
 sky130_fd_sc_hd__nor2_1 _15526_ (.A(_05967_),
    .B(net1184),
    .Y(_02645_));
 sky130_fd_sc_hd__a31o_1 _15527_ (.A1(net1184),
    .A2(_08259_),
    .A3(net570),
    .B1(_02645_),
    .X(_02646_));
 sky130_fd_sc_hd__a22o_1 _15528_ (.A1(net460),
    .A2(_02269_),
    .B1(_02646_),
    .B2(net1222),
    .X(_02647_));
 sky130_fd_sc_hd__o21a_1 _15529_ (.A1(net1780),
    .A2(net1222),
    .B1(_02481_),
    .X(_02648_));
 sky130_fd_sc_hd__nand2_1 _15530_ (.A(_02647_),
    .B(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__xnor2_1 _15531_ (.A(_02647_),
    .B(_02648_),
    .Y(_02650_));
 sky130_fd_sc_hd__nor2_1 _15532_ (.A(_02625_),
    .B(_02630_),
    .Y(_02651_));
 sky130_fd_sc_hd__and2_1 _15533_ (.A(\core.fetchProgramCounter[19] ),
    .B(_02632_),
    .X(_02652_));
 sky130_fd_sc_hd__o21ai_1 _15534_ (.A1(\core.fetchProgramCounter[19] ),
    .A2(_02632_),
    .B1(net561),
    .Y(_02653_));
 sky130_fd_sc_hd__nor2_1 _15535_ (.A(_02652_),
    .B(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__xnor2_1 _15536_ (.A(_02650_),
    .B(_02651_),
    .Y(_02655_));
 sky130_fd_sc_hd__a21oi_1 _15537_ (.A1(net1299),
    .A2(_02655_),
    .B1(net561),
    .Y(_02656_));
 sky130_fd_sc_hd__or3_1 _15538_ (.A(net1130),
    .B(_02654_),
    .C(_02656_),
    .X(_02657_));
 sky130_fd_sc_hd__o21a_1 _15539_ (.A1(\core.csr.trapReturnVector[19] ),
    .A2(net1126),
    .B1(net550),
    .X(_02658_));
 sky130_fd_sc_hd__nor2_1 _15540_ (.A(\core.csr.traps.mtvec.csrReadData[19] ),
    .B(\core.csr.traps.mcause.csrReadData[17] ),
    .Y(_02659_));
 sky130_fd_sc_hd__nand2_1 _15541_ (.A(\core.csr.traps.mtvec.csrReadData[19] ),
    .B(\core.csr.traps.mcause.csrReadData[17] ),
    .Y(_02660_));
 sky130_fd_sc_hd__nand2b_1 _15542_ (.A_N(_02659_),
    .B(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__o21a_1 _15543_ (.A1(_02638_),
    .A2(_02639_),
    .B1(_02640_),
    .X(_02662_));
 sky130_fd_sc_hd__xor2_1 _15544_ (.A(_02661_),
    .B(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__mux2_1 _15545_ (.A0(\core.csr.traps.mtvec.csrReadData[19] ),
    .A1(_02663_),
    .S(net1055),
    .X(_02664_));
 sky130_fd_sc_hd__a221o_1 _15546_ (.A1(_02657_),
    .A2(_02658_),
    .B1(_02664_),
    .B2(net541),
    .C1(net540),
    .X(_02665_));
 sky130_fd_sc_hd__o211a_1 _15547_ (.A1(\core.fetchProgramCounter[19] ),
    .A2(net522),
    .B1(_02665_),
    .C1(net1814),
    .X(_00823_));
 sky130_fd_sc_hd__and2_1 _15548_ (.A(net1751),
    .B(net569),
    .X(_02666_));
 sky130_fd_sc_hd__nand2_8 _15549_ (.A(net1751),
    .B(net569),
    .Y(_02667_));
 sky130_fd_sc_hd__a22o_1 _15550_ (.A1(_05891_),
    .A2(net1185),
    .B1(_08290_),
    .B2(_02246_),
    .X(_02668_));
 sky130_fd_sc_hd__a2bb2o_4 _15551_ (.A1_N(net462),
    .A2_N(net565),
    .B1(_02668_),
    .B2(net1223),
    .X(_02669_));
 sky130_fd_sc_hd__nor2_2 _15552_ (.A(_02667_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__xnor2_4 _15553_ (.A(_02667_),
    .B(_02669_),
    .Y(_02671_));
 sky130_fd_sc_hd__or2_1 _15554_ (.A(_02626_),
    .B(_02650_),
    .X(_02672_));
 sky130_fd_sc_hd__o21ai_1 _15555_ (.A1(_02647_),
    .A2(_02648_),
    .B1(_02625_),
    .Y(_02673_));
 sky130_fd_sc_hd__o311a_4 _15556_ (.A1(_02603_),
    .A2(_02628_),
    .A3(_02672_),
    .B1(_02673_),
    .C1(_02649_),
    .X(_02674_));
 sky130_fd_sc_hd__or3_2 _15557_ (.A(_02577_),
    .B(_02607_),
    .C(_02672_),
    .X(_02675_));
 sky130_fd_sc_hd__or2_2 _15558_ (.A(_02583_),
    .B(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__a21oi_4 _15559_ (.A1(_02674_),
    .A2(_02676_),
    .B1(_02671_),
    .Y(_02677_));
 sky130_fd_sc_hd__a311o_1 _15560_ (.A1(_02671_),
    .A2(_02674_),
    .A3(_02676_),
    .B1(_02677_),
    .C1(net559),
    .X(_02678_));
 sky130_fd_sc_hd__and3_1 _15561_ (.A(\core.fetchProgramCounter[20] ),
    .B(\core.fetchProgramCounter[19] ),
    .C(_02632_),
    .X(_02679_));
 sky130_fd_sc_hd__nor2_1 _15562_ (.A(\core.fetchProgramCounter[20] ),
    .B(_02652_),
    .Y(_02680_));
 sky130_fd_sc_hd__o31a_1 _15563_ (.A1(net569),
    .A2(_02679_),
    .A3(_02680_),
    .B1(net1125),
    .X(_02681_));
 sky130_fd_sc_hd__o21ai_1 _15564_ (.A1(\core.csr.trapReturnVector[20] ),
    .A2(net1125),
    .B1(net549),
    .Y(_02682_));
 sky130_fd_sc_hd__a21oi_1 _15565_ (.A1(_02678_),
    .A2(_02681_),
    .B1(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand2_1 _15566_ (.A(\core.csr.traps.mtvec.csrReadData[20] ),
    .B(\core.csr.traps.mcause.csrReadData[18] ),
    .Y(_02684_));
 sky130_fd_sc_hd__or2_1 _15567_ (.A(\core.csr.traps.mtvec.csrReadData[20] ),
    .B(\core.csr.traps.mcause.csrReadData[18] ),
    .X(_02685_));
 sky130_fd_sc_hd__nand2_1 _15568_ (.A(_02684_),
    .B(_02685_),
    .Y(_02686_));
 sky130_fd_sc_hd__o21a_1 _15569_ (.A1(_02659_),
    .A2(_02662_),
    .B1(_02660_),
    .X(_02687_));
 sky130_fd_sc_hd__xor2_1 _15570_ (.A(_02686_),
    .B(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__mux2_1 _15571_ (.A0(\core.csr.traps.mtvec.csrReadData[20] ),
    .A1(_02688_),
    .S(net1055),
    .X(_02689_));
 sky130_fd_sc_hd__a21o_1 _15572_ (.A1(net541),
    .A2(_02689_),
    .B1(net537),
    .X(_02690_));
 sky130_fd_sc_hd__o221a_1 _15573_ (.A1(\core.fetchProgramCounter[20] ),
    .A2(net521),
    .B1(_02683_),
    .B2(_02690_),
    .C1(net1810),
    .X(_00824_));
 sky130_fd_sc_hd__o2bb2a_1 _15574_ (.A1_N(_08324_),
    .A2_N(_02246_),
    .B1(_05816_),
    .B2(net1179),
    .X(_02691_));
 sky130_fd_sc_hd__o22a_2 _15575_ (.A1(net463),
    .A2(net565),
    .B1(_02691_),
    .B2(net1228),
    .X(_02692_));
 sky130_fd_sc_hd__or2_1 _15576_ (.A(net558),
    .B(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__and2_1 _15577_ (.A(net558),
    .B(_02692_),
    .X(_02694_));
 sky130_fd_sc_hd__xnor2_1 _15578_ (.A(net558),
    .B(_02692_),
    .Y(_02695_));
 sky130_fd_sc_hd__o21ai_1 _15579_ (.A1(_02670_),
    .A2(_02677_),
    .B1(_02695_),
    .Y(_02696_));
 sky130_fd_sc_hd__or3_1 _15580_ (.A(_02670_),
    .B(_02677_),
    .C(_02695_),
    .X(_02697_));
 sky130_fd_sc_hd__and3_2 _15581_ (.A(\core.fetchProgramCounter[21] ),
    .B(\core.fetchProgramCounter[20] ),
    .C(_02652_),
    .X(_02698_));
 sky130_fd_sc_hd__a21oi_1 _15582_ (.A1(\core.fetchProgramCounter[20] ),
    .A2(_02652_),
    .B1(\core.fetchProgramCounter[21] ),
    .Y(_02699_));
 sky130_fd_sc_hd__nor2_1 _15583_ (.A(_02698_),
    .B(_02699_),
    .Y(_02700_));
 sky130_fd_sc_hd__a31oi_1 _15584_ (.A1(net1299),
    .A2(_02696_),
    .A3(_02697_),
    .B1(net559),
    .Y(_02701_));
 sky130_fd_sc_hd__a211o_1 _15585_ (.A1(net559),
    .A2(_02700_),
    .B1(_02701_),
    .C1(_07057_),
    .X(_02702_));
 sky130_fd_sc_hd__o211a_1 _15586_ (.A1(\core.csr.trapReturnVector[21] ),
    .A2(net1125),
    .B1(net550),
    .C1(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__o21a_1 _15587_ (.A1(_02686_),
    .A2(_02687_),
    .B1(_02684_),
    .X(_02704_));
 sky130_fd_sc_hd__and2_1 _15588_ (.A(\core.csr.traps.mtvec.csrReadData[21] ),
    .B(\core.csr.traps.mcause.csrReadData[19] ),
    .X(_02705_));
 sky130_fd_sc_hd__nor2_1 _15589_ (.A(\core.csr.traps.mtvec.csrReadData[21] ),
    .B(\core.csr.traps.mcause.csrReadData[19] ),
    .Y(_02706_));
 sky130_fd_sc_hd__nor2_1 _15590_ (.A(_02705_),
    .B(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__xnor2_1 _15591_ (.A(_02704_),
    .B(_02707_),
    .Y(_02708_));
 sky130_fd_sc_hd__mux2_1 _15592_ (.A0(\core.csr.traps.mtvec.csrReadData[21] ),
    .A1(_02708_),
    .S(net1055),
    .X(_02709_));
 sky130_fd_sc_hd__a21o_1 _15593_ (.A1(net541),
    .A2(_02709_),
    .B1(net537),
    .X(_02710_));
 sky130_fd_sc_hd__o221a_1 _15594_ (.A1(\core.fetchProgramCounter[21] ),
    .A2(net521),
    .B1(_02703_),
    .B2(_02710_),
    .C1(net1810),
    .X(_00825_));
 sky130_fd_sc_hd__o2bb2a_1 _15595_ (.A1_N(_08353_),
    .A2_N(_02246_),
    .B1(_05738_),
    .B2(net1179),
    .X(_02711_));
 sky130_fd_sc_hd__o22a_4 _15596_ (.A1(net464),
    .A2(net565),
    .B1(_02711_),
    .B2(net1227),
    .X(_02712_));
 sky130_fd_sc_hd__and2_1 _15597_ (.A(net558),
    .B(_02712_),
    .X(_02713_));
 sky130_fd_sc_hd__xnor2_4 _15598_ (.A(net558),
    .B(_02712_),
    .Y(_02714_));
 sky130_fd_sc_hd__inv_2 _15599_ (.A(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__o31a_1 _15600_ (.A1(_02670_),
    .A2(_02677_),
    .A3(_02694_),
    .B1(_02693_),
    .X(_02716_));
 sky130_fd_sc_hd__o311a_1 _15601_ (.A1(_02670_),
    .A2(_02677_),
    .A3(_02694_),
    .B1(_02715_),
    .C1(_02693_),
    .X(_02717_));
 sky130_fd_sc_hd__xnor2_2 _15602_ (.A(_02714_),
    .B(_02716_),
    .Y(_02718_));
 sky130_fd_sc_hd__nand2_1 _15603_ (.A(\core.fetchProgramCounter[22] ),
    .B(_02698_),
    .Y(_02719_));
 sky130_fd_sc_hd__or2_1 _15604_ (.A(\core.fetchProgramCounter[22] ),
    .B(_02698_),
    .X(_02720_));
 sky130_fd_sc_hd__a31o_1 _15605_ (.A1(net560),
    .A2(_02719_),
    .A3(_02720_),
    .B1(net1130),
    .X(_02721_));
 sky130_fd_sc_hd__a21o_1 _15606_ (.A1(net569),
    .A2(_02718_),
    .B1(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__o211a_1 _15607_ (.A1(\core.csr.trapReturnVector[22] ),
    .A2(net1125),
    .B1(net552),
    .C1(_02722_),
    .X(_02723_));
 sky130_fd_sc_hd__and2_1 _15608_ (.A(\core.csr.traps.mtvec.csrReadData[22] ),
    .B(\core.csr.traps.mcause.csrReadData[20] ),
    .X(_02724_));
 sky130_fd_sc_hd__nor2_1 _15609_ (.A(\core.csr.traps.mtvec.csrReadData[22] ),
    .B(\core.csr.traps.mcause.csrReadData[20] ),
    .Y(_02725_));
 sky130_fd_sc_hd__nor2_1 _15610_ (.A(_02724_),
    .B(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__o21ba_2 _15611_ (.A1(_02704_),
    .A2(_02706_),
    .B1_N(_02705_),
    .X(_02727_));
 sky130_fd_sc_hd__xnor2_1 _15612_ (.A(_02726_),
    .B(_02727_),
    .Y(_02728_));
 sky130_fd_sc_hd__mux2_1 _15613_ (.A0(\core.csr.traps.mtvec.csrReadData[22] ),
    .A1(_02728_),
    .S(net1056),
    .X(_02729_));
 sky130_fd_sc_hd__a21o_1 _15614_ (.A1(net543),
    .A2(_02729_),
    .B1(net537),
    .X(_02730_));
 sky130_fd_sc_hd__o221a_1 _15615_ (.A1(\core.fetchProgramCounter[22] ),
    .A2(net521),
    .B1(_02723_),
    .B2(_02730_),
    .C1(net1816),
    .X(_00826_));
 sky130_fd_sc_hd__o22a_1 _15616_ (.A1(_05661_),
    .A2(net1179),
    .B1(_08385_),
    .B2(_02247_),
    .X(_02731_));
 sky130_fd_sc_hd__o22a_1 _15617_ (.A1(_03824_),
    .A2(net565),
    .B1(_02731_),
    .B2(net1227),
    .X(_02732_));
 sky130_fd_sc_hd__xnor2_1 _15618_ (.A(_02667_),
    .B(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__o21ai_1 _15619_ (.A1(_02713_),
    .A2(_02717_),
    .B1(_02733_),
    .Y(_02734_));
 sky130_fd_sc_hd__or3_1 _15620_ (.A(_02713_),
    .B(_02717_),
    .C(_02733_),
    .X(_02735_));
 sky130_fd_sc_hd__and3_2 _15621_ (.A(\core.fetchProgramCounter[23] ),
    .B(\core.fetchProgramCounter[22] ),
    .C(_02698_),
    .X(_02736_));
 sky130_fd_sc_hd__a21oi_1 _15622_ (.A1(\core.fetchProgramCounter[22] ),
    .A2(_02698_),
    .B1(\core.fetchProgramCounter[23] ),
    .Y(_02737_));
 sky130_fd_sc_hd__or3_1 _15623_ (.A(net569),
    .B(_02736_),
    .C(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__a31o_1 _15624_ (.A1(net1299),
    .A2(_02734_),
    .A3(_02735_),
    .B1(net559),
    .X(_02739_));
 sky130_fd_sc_hd__nand3_1 _15625_ (.A(net1126),
    .B(_02738_),
    .C(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__o21a_1 _15626_ (.A1(\core.csr.trapReturnVector[23] ),
    .A2(net1126),
    .B1(net550),
    .X(_02741_));
 sky130_fd_sc_hd__o21bai_2 _15627_ (.A1(_02725_),
    .A2(_02727_),
    .B1_N(_02724_),
    .Y(_02742_));
 sky130_fd_sc_hd__and2_1 _15628_ (.A(\core.csr.traps.mtvec.csrReadData[23] ),
    .B(\core.csr.traps.mcause.csrReadData[21] ),
    .X(_02743_));
 sky130_fd_sc_hd__or2_1 _15629_ (.A(\core.csr.traps.mtvec.csrReadData[23] ),
    .B(\core.csr.traps.mcause.csrReadData[21] ),
    .X(_02744_));
 sky130_fd_sc_hd__nand2b_1 _15630_ (.A_N(_02743_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__xnor2_1 _15631_ (.A(_02742_),
    .B(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__mux2_1 _15632_ (.A0(\core.csr.traps.mtvec.csrReadData[23] ),
    .A1(_02746_),
    .S(net1055),
    .X(_02747_));
 sky130_fd_sc_hd__a221o_1 _15633_ (.A1(_02740_),
    .A2(_02741_),
    .B1(_02747_),
    .B2(net542),
    .C1(net540),
    .X(_02748_));
 sky130_fd_sc_hd__o211a_1 _15634_ (.A1(\core.fetchProgramCounter[23] ),
    .A2(net522),
    .B1(_02748_),
    .C1(net1813),
    .X(_00827_));
 sky130_fd_sc_hd__o2bb2a_1 _15635_ (.A1_N(_08415_),
    .A2_N(_02246_),
    .B1(_05587_),
    .B2(net1179),
    .X(_02749_));
 sky130_fd_sc_hd__o22a_2 _15636_ (.A1(net466),
    .A2(net565),
    .B1(_02749_),
    .B2(net1227),
    .X(_02750_));
 sky130_fd_sc_hd__xnor2_1 _15637_ (.A(net557),
    .B(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__or4_1 _15638_ (.A(_02671_),
    .B(_02695_),
    .C(_02714_),
    .D(_02733_),
    .X(_02752_));
 sky130_fd_sc_hd__or3b_1 _15639_ (.A(_02692_),
    .B(_02712_),
    .C_N(_02732_),
    .X(_02753_));
 sky130_fd_sc_hd__nand2_1 _15640_ (.A(net558),
    .B(_02753_),
    .Y(_02754_));
 sky130_fd_sc_hd__o221a_1 _15641_ (.A1(_02667_),
    .A2(_02669_),
    .B1(_02674_),
    .B2(_02752_),
    .C1(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__o31a_2 _15642_ (.A1(_02583_),
    .A2(_02675_),
    .A3(_02752_),
    .B1(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__and2_1 _15643_ (.A(_02751_),
    .B(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__nor2_1 _15644_ (.A(_02751_),
    .B(_02756_),
    .Y(_02758_));
 sky130_fd_sc_hd__or2_2 _15645_ (.A(_02757_),
    .B(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__xnor2_1 _15646_ (.A(\core.fetchProgramCounter[24] ),
    .B(_02736_),
    .Y(_02760_));
 sky130_fd_sc_hd__a221o_1 _15647_ (.A1(_03811_),
    .A2(net1130),
    .B1(net567),
    .B2(_02760_),
    .C1(net542),
    .X(_02761_));
 sky130_fd_sc_hd__a21oi_1 _15648_ (.A1(net569),
    .A2(_02759_),
    .B1(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__nand2_1 _15649_ (.A(\core.csr.traps.mtvec.csrReadData[24] ),
    .B(\core.csr.traps.mcause.csrReadData[22] ),
    .Y(_02763_));
 sky130_fd_sc_hd__or2_1 _15650_ (.A(\core.csr.traps.mtvec.csrReadData[24] ),
    .B(\core.csr.traps.mcause.csrReadData[22] ),
    .X(_02764_));
 sky130_fd_sc_hd__nand2_1 _15651_ (.A(_02763_),
    .B(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__a21o_1 _15652_ (.A1(_02742_),
    .A2(_02744_),
    .B1(_02743_),
    .X(_02766_));
 sky130_fd_sc_hd__xnor2_1 _15653_ (.A(_02765_),
    .B(_02766_),
    .Y(_02767_));
 sky130_fd_sc_hd__mux2_1 _15654_ (.A0(\core.csr.traps.mtvec.csrReadData[24] ),
    .A1(_02767_),
    .S(net1056),
    .X(_02768_));
 sky130_fd_sc_hd__a21o_1 _15655_ (.A1(net542),
    .A2(_02768_),
    .B1(net537),
    .X(_02769_));
 sky130_fd_sc_hd__o221a_1 _15656_ (.A1(\core.fetchProgramCounter[24] ),
    .A2(net522),
    .B1(_02762_),
    .B2(_02769_),
    .C1(net1812),
    .X(_00828_));
 sky130_fd_sc_hd__o2bb2a_1 _15657_ (.A1_N(_08447_),
    .A2_N(_02246_),
    .B1(_05512_),
    .B2(net1179),
    .X(_02770_));
 sky130_fd_sc_hd__o22a_1 _15658_ (.A1(net467),
    .A2(net565),
    .B1(_02770_),
    .B2(net1227),
    .X(_02771_));
 sky130_fd_sc_hd__xnor2_1 _15659_ (.A(net557),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__a21o_1 _15660_ (.A1(net557),
    .A2(_02750_),
    .B1(_02758_),
    .X(_02773_));
 sky130_fd_sc_hd__or2_1 _15661_ (.A(\core.csr.trapReturnVector[25] ),
    .B(net1126),
    .X(_02774_));
 sky130_fd_sc_hd__and3_2 _15662_ (.A(\core.fetchProgramCounter[25] ),
    .B(\core.fetchProgramCounter[24] ),
    .C(_02736_),
    .X(_02775_));
 sky130_fd_sc_hd__a21oi_1 _15663_ (.A1(\core.fetchProgramCounter[24] ),
    .A2(_02736_),
    .B1(\core.fetchProgramCounter[25] ),
    .Y(_02776_));
 sky130_fd_sc_hd__nor2_1 _15664_ (.A(_02775_),
    .B(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__xor2_1 _15665_ (.A(_02772_),
    .B(_02773_),
    .X(_02778_));
 sky130_fd_sc_hd__a21oi_2 _15666_ (.A1(net1299),
    .A2(_02778_),
    .B1(net559),
    .Y(_02779_));
 sky130_fd_sc_hd__a211o_1 _15667_ (.A1(net560),
    .A2(_02777_),
    .B1(_02779_),
    .C1(net1130),
    .X(_02780_));
 sky130_fd_sc_hd__a21bo_1 _15668_ (.A1(_02764_),
    .A2(_02766_),
    .B1_N(_02763_),
    .X(_02781_));
 sky130_fd_sc_hd__and2_1 _15669_ (.A(\core.csr.traps.mtvec.csrReadData[25] ),
    .B(\core.csr.traps.mcause.csrReadData[23] ),
    .X(_02782_));
 sky130_fd_sc_hd__nor2_1 _15670_ (.A(\core.csr.traps.mtvec.csrReadData[25] ),
    .B(\core.csr.traps.mcause.csrReadData[23] ),
    .Y(_02783_));
 sky130_fd_sc_hd__nor2_1 _15671_ (.A(_02782_),
    .B(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__xnor2_1 _15672_ (.A(_02781_),
    .B(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__nand2_1 _15673_ (.A(net1056),
    .B(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__o211a_1 _15674_ (.A1(\core.csr.traps.mtvec.csrReadData[25] ),
    .A2(net1055),
    .B1(_02786_),
    .C1(net542),
    .X(_02787_));
 sky130_fd_sc_hd__a311o_1 _15675_ (.A1(net550),
    .A2(_02774_),
    .A3(_02780_),
    .B1(_02787_),
    .C1(net537),
    .X(_02788_));
 sky130_fd_sc_hd__o211a_1 _15676_ (.A1(\core.fetchProgramCounter[25] ),
    .A2(net521),
    .B1(_02788_),
    .C1(net1812),
    .X(_00829_));
 sky130_fd_sc_hd__nand2_1 _15677_ (.A(\core.fetchProgramCounter[26] ),
    .B(_02775_),
    .Y(_02789_));
 sky130_fd_sc_hd__or2_1 _15678_ (.A(\core.fetchProgramCounter[26] ),
    .B(_02775_),
    .X(_02790_));
 sky130_fd_sc_hd__a31o_1 _15679_ (.A1(net560),
    .A2(_02789_),
    .A3(_02790_),
    .B1(net1130),
    .X(_02791_));
 sky130_fd_sc_hd__o2bb2a_1 _15680_ (.A1_N(_08480_),
    .A2_N(_02246_),
    .B1(_05438_),
    .B2(net1179),
    .X(_02792_));
 sky130_fd_sc_hd__o22a_1 _15681_ (.A1(net468),
    .A2(net565),
    .B1(_02792_),
    .B2(net1227),
    .X(_02793_));
 sky130_fd_sc_hd__nor2_1 _15682_ (.A(net557),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__and2_1 _15683_ (.A(net557),
    .B(_02793_),
    .X(_02795_));
 sky130_fd_sc_hd__or2_1 _15684_ (.A(_02794_),
    .B(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__inv_2 _15685_ (.A(_02796_),
    .Y(_02797_));
 sky130_fd_sc_hd__or2_1 _15686_ (.A(_02751_),
    .B(_02772_),
    .X(_02798_));
 sky130_fd_sc_hd__or2_1 _15687_ (.A(_02750_),
    .B(_02771_),
    .X(_02799_));
 sky130_fd_sc_hd__a2bb2o_2 _15688_ (.A1_N(_02756_),
    .A2_N(_02798_),
    .B1(_02799_),
    .B2(net557),
    .X(_02800_));
 sky130_fd_sc_hd__xnor2_2 _15689_ (.A(_02797_),
    .B(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__nor2_1 _15690_ (.A(net560),
    .B(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__o221a_1 _15691_ (.A1(\core.csr.trapReturnVector[26] ),
    .A2(net1125),
    .B1(_02791_),
    .B2(_02802_),
    .C1(net550),
    .X(_02803_));
 sky130_fd_sc_hd__a21oi_2 _15692_ (.A1(_02781_),
    .A2(_02784_),
    .B1(_02782_),
    .Y(_02804_));
 sky130_fd_sc_hd__nor2_1 _15693_ (.A(\core.csr.traps.mtvec.csrReadData[26] ),
    .B(\core.csr.traps.mcause.csrReadData[24] ),
    .Y(_02805_));
 sky130_fd_sc_hd__nand2_1 _15694_ (.A(\core.csr.traps.mtvec.csrReadData[26] ),
    .B(\core.csr.traps.mcause.csrReadData[24] ),
    .Y(_02806_));
 sky130_fd_sc_hd__and2b_1 _15695_ (.A_N(_02805_),
    .B(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__xnor2_1 _15696_ (.A(_02804_),
    .B(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__mux2_1 _15697_ (.A0(\core.csr.traps.mtvec.csrReadData[26] ),
    .A1(_02808_),
    .S(net1056),
    .X(_02809_));
 sky130_fd_sc_hd__a21o_1 _15698_ (.A1(net542),
    .A2(_02809_),
    .B1(net537),
    .X(_02810_));
 sky130_fd_sc_hd__o221a_1 _15699_ (.A1(\core.fetchProgramCounter[26] ),
    .A2(net521),
    .B1(_02803_),
    .B2(_02810_),
    .C1(net1812),
    .X(_00830_));
 sky130_fd_sc_hd__o22a_1 _15700_ (.A1(_05364_),
    .A2(net1179),
    .B1(_08513_),
    .B2(_02247_),
    .X(_02811_));
 sky130_fd_sc_hd__o2bb2a_2 _15701_ (.A1_N(net469),
    .A2_N(_02269_),
    .B1(_02811_),
    .B2(net1227),
    .X(_02812_));
 sky130_fd_sc_hd__xnor2_2 _15702_ (.A(_02667_),
    .B(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__a21oi_1 _15703_ (.A1(_02797_),
    .A2(_02800_),
    .B1(_02795_),
    .Y(_02814_));
 sky130_fd_sc_hd__and3_2 _15704_ (.A(\core.fetchProgramCounter[27] ),
    .B(\core.fetchProgramCounter[26] ),
    .C(_02775_),
    .X(_02815_));
 sky130_fd_sc_hd__a21oi_1 _15705_ (.A1(\core.fetchProgramCounter[26] ),
    .A2(_02775_),
    .B1(\core.fetchProgramCounter[27] ),
    .Y(_02816_));
 sky130_fd_sc_hd__nor2_1 _15706_ (.A(_02815_),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__xnor2_1 _15707_ (.A(_02813_),
    .B(_02814_),
    .Y(_02818_));
 sky130_fd_sc_hd__a21oi_2 _15708_ (.A1(net1299),
    .A2(_02818_),
    .B1(net559),
    .Y(_02819_));
 sky130_fd_sc_hd__a211o_1 _15709_ (.A1(net560),
    .A2(_02817_),
    .B1(_02819_),
    .C1(net1130),
    .X(_02820_));
 sky130_fd_sc_hd__o21a_1 _15710_ (.A1(\core.csr.trapReturnVector[27] ),
    .A2(net1126),
    .B1(net552),
    .X(_02821_));
 sky130_fd_sc_hd__or2_1 _15711_ (.A(\core.csr.traps.mtvec.csrReadData[27] ),
    .B(\core.csr.traps.mcause.csrReadData[25] ),
    .X(_02822_));
 sky130_fd_sc_hd__nand2_1 _15712_ (.A(\core.csr.traps.mtvec.csrReadData[27] ),
    .B(\core.csr.traps.mcause.csrReadData[25] ),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_1 _15713_ (.A(_02822_),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__o21ai_2 _15714_ (.A1(_02804_),
    .A2(_02805_),
    .B1(_02806_),
    .Y(_02825_));
 sky130_fd_sc_hd__xnor2_1 _15715_ (.A(_02824_),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__mux2_1 _15716_ (.A0(\core.csr.traps.mtvec.csrReadData[27] ),
    .A1(_02826_),
    .S(net1056),
    .X(_02827_));
 sky130_fd_sc_hd__a221o_1 _15717_ (.A1(_02820_),
    .A2(_02821_),
    .B1(_02827_),
    .B2(net542),
    .C1(net537),
    .X(_02828_));
 sky130_fd_sc_hd__o211a_1 _15718_ (.A1(\core.fetchProgramCounter[27] ),
    .A2(net522),
    .B1(_02828_),
    .C1(net1812),
    .X(_00831_));
 sky130_fd_sc_hd__o2bb2a_1 _15719_ (.A1_N(_08542_),
    .A2_N(_02246_),
    .B1(_05292_),
    .B2(net1180),
    .X(_02829_));
 sky130_fd_sc_hd__o22a_1 _15720_ (.A1(net470),
    .A2(net565),
    .B1(_02829_),
    .B2(net1227),
    .X(_02830_));
 sky130_fd_sc_hd__nor2_1 _15721_ (.A(net557),
    .B(_02830_),
    .Y(_02831_));
 sky130_fd_sc_hd__and2_1 _15722_ (.A(net557),
    .B(_02830_),
    .X(_02832_));
 sky130_fd_sc_hd__nor2_1 _15723_ (.A(_02831_),
    .B(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__inv_2 _15724_ (.A(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__or3b_1 _15725_ (.A(_02793_),
    .B(_02799_),
    .C_N(_02812_),
    .X(_02835_));
 sky130_fd_sc_hd__nand2_1 _15726_ (.A(net557),
    .B(_02835_),
    .Y(_02836_));
 sky130_fd_sc_hd__o41a_2 _15727_ (.A1(_02756_),
    .A2(_02796_),
    .A3(_02798_),
    .A4(_02813_),
    .B1(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__xnor2_1 _15728_ (.A(_02834_),
    .B(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__and2_1 _15729_ (.A(\core.fetchProgramCounter[28] ),
    .B(_02815_),
    .X(_02839_));
 sky130_fd_sc_hd__nor2_1 _15730_ (.A(\core.fetchProgramCounter[28] ),
    .B(_02815_),
    .Y(_02840_));
 sky130_fd_sc_hd__o21ai_1 _15731_ (.A1(_02839_),
    .A2(_02840_),
    .B1(net567),
    .Y(_02841_));
 sky130_fd_sc_hd__o211ai_1 _15732_ (.A1(\core.csr.trapReturnVector[28] ),
    .A2(net1125),
    .B1(net549),
    .C1(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__a21oi_1 _15733_ (.A1(net569),
    .A2(_02838_),
    .B1(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__or2_1 _15734_ (.A(\core.csr.traps.mtvec.csrReadData[28] ),
    .B(\core.csr.traps.mcause.csrReadData[26] ),
    .X(_02844_));
 sky130_fd_sc_hd__nand2_1 _15735_ (.A(\core.csr.traps.mtvec.csrReadData[28] ),
    .B(\core.csr.traps.mcause.csrReadData[26] ),
    .Y(_02845_));
 sky130_fd_sc_hd__nand2_1 _15736_ (.A(_02844_),
    .B(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__a21boi_2 _15737_ (.A1(_02822_),
    .A2(_02825_),
    .B1_N(_02823_),
    .Y(_02847_));
 sky130_fd_sc_hd__xor2_1 _15738_ (.A(_02846_),
    .B(_02847_),
    .X(_02848_));
 sky130_fd_sc_hd__mux2_1 _15739_ (.A0(\core.csr.traps.mtvec.csrReadData[28] ),
    .A1(_02848_),
    .S(net1055),
    .X(_02849_));
 sky130_fd_sc_hd__a21o_1 _15740_ (.A1(net541),
    .A2(_02849_),
    .B1(net537),
    .X(_02850_));
 sky130_fd_sc_hd__o221a_1 _15741_ (.A1(\core.fetchProgramCounter[28] ),
    .A2(net521),
    .B1(_02843_),
    .B2(_02850_),
    .C1(net1808),
    .X(_00832_));
 sky130_fd_sc_hd__o22a_1 _15742_ (.A1(_05217_),
    .A2(net1180),
    .B1(_08575_),
    .B2(_02247_),
    .X(_02851_));
 sky130_fd_sc_hd__o22a_2 _15743_ (.A1(net471),
    .A2(net565),
    .B1(_02851_),
    .B2(net1227),
    .X(_02852_));
 sky130_fd_sc_hd__xnor2_2 _15744_ (.A(net557),
    .B(_02852_),
    .Y(_02853_));
 sky130_fd_sc_hd__o21ba_1 _15745_ (.A1(_02834_),
    .A2(_02837_),
    .B1_N(_02832_),
    .X(_02854_));
 sky130_fd_sc_hd__and3_1 _15746_ (.A(\core.fetchProgramCounter[29] ),
    .B(\core.fetchProgramCounter[28] ),
    .C(_02815_),
    .X(_02855_));
 sky130_fd_sc_hd__o21ai_1 _15747_ (.A1(\core.fetchProgramCounter[29] ),
    .A2(_02839_),
    .B1(net559),
    .Y(_02856_));
 sky130_fd_sc_hd__nor2_1 _15748_ (.A(_02855_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__xnor2_1 _15749_ (.A(_02853_),
    .B(_02854_),
    .Y(_02858_));
 sky130_fd_sc_hd__a21oi_1 _15750_ (.A1(net1299),
    .A2(_02858_),
    .B1(net559),
    .Y(_02859_));
 sky130_fd_sc_hd__or3_1 _15751_ (.A(net1130),
    .B(_02857_),
    .C(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__o21a_1 _15752_ (.A1(\core.csr.trapReturnVector[29] ),
    .A2(net1125),
    .B1(net549),
    .X(_02861_));
 sky130_fd_sc_hd__nor2_1 _15753_ (.A(\core.csr.traps.mtvec.csrReadData[29] ),
    .B(\core.csr.traps.mcause.csrReadData[27] ),
    .Y(_02862_));
 sky130_fd_sc_hd__nand2_1 _15754_ (.A(\core.csr.traps.mtvec.csrReadData[29] ),
    .B(\core.csr.traps.mcause.csrReadData[27] ),
    .Y(_02863_));
 sky130_fd_sc_hd__nand2b_1 _15755_ (.A_N(_02862_),
    .B(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__nand2_1 _15756_ (.A(_02845_),
    .B(_02847_),
    .Y(_02865_));
 sky130_fd_sc_hd__nand2_1 _15757_ (.A(_02844_),
    .B(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__xor2_1 _15758_ (.A(_02864_),
    .B(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__mux2_1 _15759_ (.A0(\core.csr.traps.mtvec.csrReadData[29] ),
    .A1(_02867_),
    .S(net1055),
    .X(_02868_));
 sky130_fd_sc_hd__a221o_1 _15760_ (.A1(_02860_),
    .A2(_02861_),
    .B1(_02868_),
    .B2(net541),
    .C1(net537),
    .X(_02869_));
 sky130_fd_sc_hd__o211a_1 _15761_ (.A1(\core.fetchProgramCounter[29] ),
    .A2(net521),
    .B1(_02869_),
    .C1(net1808),
    .X(_00833_));
 sky130_fd_sc_hd__o2bb2a_1 _15762_ (.A1_N(_08607_),
    .A2_N(_02246_),
    .B1(_05144_),
    .B2(net1180),
    .X(_02870_));
 sky130_fd_sc_hd__o22a_1 _15763_ (.A1(net473),
    .A2(net565),
    .B1(_02870_),
    .B2(net1227),
    .X(_02871_));
 sky130_fd_sc_hd__nand2_1 _15764_ (.A(_02666_),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__or2_1 _15765_ (.A(net558),
    .B(_02871_),
    .X(_02873_));
 sky130_fd_sc_hd__and2_1 _15766_ (.A(_02872_),
    .B(_02873_),
    .X(_02874_));
 sky130_fd_sc_hd__inv_2 _15767_ (.A(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__o21ai_1 _15768_ (.A1(_02830_),
    .A2(_02852_),
    .B1(net558),
    .Y(_02876_));
 sky130_fd_sc_hd__o31a_1 _15769_ (.A1(_02834_),
    .A2(_02837_),
    .A3(_02853_),
    .B1(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__xnor2_1 _15770_ (.A(_02874_),
    .B(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__nand2_1 _15771_ (.A(\core.fetchProgramCounter[30] ),
    .B(_02855_),
    .Y(_02879_));
 sky130_fd_sc_hd__or2_1 _15772_ (.A(\core.fetchProgramCounter[30] ),
    .B(_02855_),
    .X(_02880_));
 sky130_fd_sc_hd__a31o_1 _15773_ (.A1(net559),
    .A2(_02879_),
    .A3(_02880_),
    .B1(net1130),
    .X(_02881_));
 sky130_fd_sc_hd__a21o_1 _15774_ (.A1(net569),
    .A2(_02878_),
    .B1(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__o211a_1 _15775_ (.A1(\core.csr.trapReturnVector[30] ),
    .A2(net1125),
    .B1(net549),
    .C1(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__and2_1 _15776_ (.A(\core.csr.traps.mtvec.csrReadData[30] ),
    .B(\core.csr.traps.mcause.csrReadData[28] ),
    .X(_02884_));
 sky130_fd_sc_hd__or2_1 _15777_ (.A(\core.csr.traps.mtvec.csrReadData[30] ),
    .B(\core.csr.traps.mcause.csrReadData[28] ),
    .X(_02885_));
 sky130_fd_sc_hd__nand2b_1 _15778_ (.A_N(_02884_),
    .B(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__o21ai_2 _15779_ (.A1(_02862_),
    .A2(_02866_),
    .B1(_02863_),
    .Y(_02887_));
 sky130_fd_sc_hd__xnor2_1 _15780_ (.A(_02886_),
    .B(_02887_),
    .Y(_02888_));
 sky130_fd_sc_hd__mux2_1 _15781_ (.A0(\core.csr.traps.mtvec.csrReadData[30] ),
    .A1(_02888_),
    .S(net1055),
    .X(_02889_));
 sky130_fd_sc_hd__a21o_1 _15782_ (.A1(net541),
    .A2(_02889_),
    .B1(net537),
    .X(_02890_));
 sky130_fd_sc_hd__o221a_1 _15783_ (.A1(\core.fetchProgramCounter[30] ),
    .A2(net521),
    .B1(_02883_),
    .B2(_02890_),
    .C1(net1810),
    .X(_00834_));
 sky130_fd_sc_hd__o21ai_1 _15784_ (.A1(_02875_),
    .A2(_02877_),
    .B1(_02872_),
    .Y(_02891_));
 sky130_fd_sc_hd__o22a_1 _15785_ (.A1(_06612_),
    .A2(net1180),
    .B1(_08640_),
    .B2(_02247_),
    .X(_02892_));
 sky130_fd_sc_hd__o22a_1 _15786_ (.A1(_03823_),
    .A2(net566),
    .B1(_02892_),
    .B2(net1228),
    .X(_02893_));
 sky130_fd_sc_hd__xnor2_1 _15787_ (.A(net558),
    .B(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__xnor2_1 _15788_ (.A(_02891_),
    .B(_02894_),
    .Y(_02895_));
 sky130_fd_sc_hd__a21o_1 _15789_ (.A1(net1299),
    .A2(_02895_),
    .B1(net559),
    .X(_02896_));
 sky130_fd_sc_hd__or2_1 _15790_ (.A(\core.fetchProgramCounter[31] ),
    .B(_02879_),
    .X(_02897_));
 sky130_fd_sc_hd__nand2_1 _15791_ (.A(\core.fetchProgramCounter[31] ),
    .B(_02879_),
    .Y(_02898_));
 sky130_fd_sc_hd__a31o_1 _15792_ (.A1(net1125),
    .A2(_02897_),
    .A3(_02898_),
    .B1(net569),
    .X(_02899_));
 sky130_fd_sc_hd__o21ai_1 _15793_ (.A1(\core.csr.trapReturnVector[31] ),
    .A2(net1125),
    .B1(net549),
    .Y(_02900_));
 sky130_fd_sc_hd__a21oi_1 _15794_ (.A1(_02896_),
    .A2(_02899_),
    .B1(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__a21oi_1 _15795_ (.A1(_02885_),
    .A2(_02887_),
    .B1(_02884_),
    .Y(_02902_));
 sky130_fd_sc_hd__xnor2_1 _15796_ (.A(\core.csr.traps.mcause.csrReadData[29] ),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__a21oi_1 _15797_ (.A1(net1055),
    .A2(_02903_),
    .B1(\core.csr.traps.mtvec.csrReadData[31] ),
    .Y(_02904_));
 sky130_fd_sc_hd__a31o_1 _15798_ (.A1(\core.csr.traps.mtvec.csrReadData[31] ),
    .A2(net1055),
    .A3(_02903_),
    .B1(net549),
    .X(_02905_));
 sky130_fd_sc_hd__o21ai_1 _15799_ (.A1(_02904_),
    .A2(_02905_),
    .B1(net521),
    .Y(_02906_));
 sky130_fd_sc_hd__o221a_1 _15800_ (.A1(\core.fetchProgramCounter[31] ),
    .A2(net521),
    .B1(_02901_),
    .B2(_02906_),
    .C1(net1810),
    .X(_00835_));
 sky130_fd_sc_hd__nor2_2 _15801_ (.A(_08760_),
    .B(_08763_),
    .Y(_02907_));
 sky130_fd_sc_hd__mux2_1 _15802_ (.A0(\core.registers[10][0] ),
    .A1(net1077),
    .S(net808),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _15803_ (.A0(\core.registers[10][1] ),
    .A1(net1080),
    .S(net806),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _15804_ (.A0(\core.registers[10][2] ),
    .A1(net1086),
    .S(net808),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _15805_ (.A0(\core.registers[10][3] ),
    .A1(net1090),
    .S(net808),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _15806_ (.A0(\core.registers[10][4] ),
    .A1(net1029),
    .S(net806),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _15807_ (.A0(\core.registers[10][5] ),
    .A1(net1031),
    .S(net806),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _15808_ (.A0(\core.registers[10][6] ),
    .A1(net1036),
    .S(net806),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _15809_ (.A0(\core.registers[10][7] ),
    .A1(net1139),
    .S(net806),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _15810_ (.A0(\core.registers[10][8] ),
    .A1(net897),
    .S(net806),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _15811_ (.A0(\core.registers[10][9] ),
    .A1(net900),
    .S(net807),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _15812_ (.A0(\core.registers[10][10] ),
    .A1(net757),
    .S(net806),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _15813_ (.A0(\core.registers[10][11] ),
    .A1(net761),
    .S(net807),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _15814_ (.A0(\core.registers[10][12] ),
    .A1(net728),
    .S(net807),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _15815_ (.A0(\core.registers[10][13] ),
    .A1(net732),
    .S(net807),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _15816_ (.A0(\core.registers[10][14] ),
    .A1(net736),
    .S(net805),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _15817_ (.A0(\core.registers[10][15] ),
    .A1(net740),
    .S(net808),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _15818_ (.A0(\core.registers[10][16] ),
    .A1(net832),
    .S(net806),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _15819_ (.A0(\core.registers[10][17] ),
    .A1(net834),
    .S(net805),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _15820_ (.A0(\core.registers[10][18] ),
    .A1(net840),
    .S(net807),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _15821_ (.A0(\core.registers[10][19] ),
    .A1(net843),
    .S(net805),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _15822_ (.A0(\core.registers[10][20] ),
    .A1(net847),
    .S(net805),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _15823_ (.A0(\core.registers[10][21] ),
    .A1(net850),
    .S(net805),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _15824_ (.A0(\core.registers[10][22] ),
    .A1(net855),
    .S(net806),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _15825_ (.A0(\core.registers[10][23] ),
    .A1(net860),
    .S(net805),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _15826_ (.A0(\core.registers[10][24] ),
    .A1(net992),
    .S(net805),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _15827_ (.A0(\core.registers[10][25] ),
    .A1(net996),
    .S(net805),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _15828_ (.A0(\core.registers[10][26] ),
    .A1(net1000),
    .S(net805),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _15829_ (.A0(\core.registers[10][27] ),
    .A1(net865),
    .S(net806),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _15830_ (.A0(\core.registers[10][28] ),
    .A1(net869),
    .S(net807),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _15831_ (.A0(\core.registers[10][29] ),
    .A1(net873),
    .S(net807),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _15832_ (.A0(\core.registers[10][30] ),
    .A1(net880),
    .S(net807),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _15833_ (.A0(\core.registers[10][31] ),
    .A1(net1026),
    .S(net805),
    .X(_00867_));
 sky130_fd_sc_hd__nor3_4 _15834_ (.A(_07037_),
    .B(_01915_),
    .C(_01917_),
    .Y(_02908_));
 sky130_fd_sc_hd__and3_1 _15835_ (.A(_06702_),
    .B(_07005_),
    .C(_07008_),
    .X(_02909_));
 sky130_fd_sc_hd__a22oi_4 _15836_ (.A1(\jtag.managementReadData[2] ),
    .A2(net1305),
    .B1(net1197),
    .B2(net237),
    .Y(_02910_));
 sky130_fd_sc_hd__nand2_1 _15837_ (.A(_02908_),
    .B(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__o211a_1 _15838_ (.A1(\core.management_interruptEnable ),
    .A2(_02908_),
    .B1(_02911_),
    .C1(net1846),
    .X(_00900_));
 sky130_fd_sc_hd__a22oi_2 _15839_ (.A1(\jtag.managementReadData[1] ),
    .A2(net1305),
    .B1(net1197),
    .B2(net226),
    .Y(_02912_));
 sky130_fd_sc_hd__nand2_1 _15840_ (.A(_02908_),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__o211a_1 _15841_ (.A1(\coreManagement.control[1] ),
    .A2(_02908_),
    .B1(_02913_),
    .C1(net1839),
    .X(_00901_));
 sky130_fd_sc_hd__a22oi_2 _15842_ (.A1(\jtag.managementReadData[0] ),
    .A2(net1305),
    .B1(net1197),
    .B2(net215),
    .Y(_02914_));
 sky130_fd_sc_hd__nand2_1 _15843_ (.A(_02908_),
    .B(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__o211a_1 _15844_ (.A1(net1724),
    .A2(_02908_),
    .B1(_02915_),
    .C1(net1839),
    .X(_00902_));
 sky130_fd_sc_hd__nor2_8 _15845_ (.A(_03817_),
    .B(_06839_),
    .Y(_02916_));
 sky130_fd_sc_hd__or2_4 _15846_ (.A(\jtag.state[3] ),
    .B(\jtag.state[2] ),
    .X(_02917_));
 sky130_fd_sc_hd__nor2_8 _15847_ (.A(_06834_),
    .B(_02917_),
    .Y(_02918_));
 sky130_fd_sc_hd__or2_4 _15848_ (.A(_06834_),
    .B(_02917_),
    .X(_02919_));
 sky130_fd_sc_hd__or2_4 _15849_ (.A(_06847_),
    .B(_02918_),
    .X(_02920_));
 sky130_fd_sc_hd__and2_1 _15850_ (.A(_02916_),
    .B(_02920_),
    .X(_02921_));
 sky130_fd_sc_hd__nand2_2 _15851_ (.A(_02916_),
    .B(_02920_),
    .Y(_02922_));
 sky130_fd_sc_hd__and2_2 _15852_ (.A(_02916_),
    .B(_02918_),
    .X(_02923_));
 sky130_fd_sc_hd__nand2_4 _15853_ (.A(_02916_),
    .B(_02918_),
    .Y(_02924_));
 sky130_fd_sc_hd__nand2_1 _15854_ (.A(net188),
    .B(_02919_),
    .Y(_02925_));
 sky130_fd_sc_hd__a221o_1 _15855_ (.A1(net188),
    .A2(net1285),
    .B1(net1163),
    .B2(net447),
    .C1(net1167),
    .X(_02926_));
 sky130_fd_sc_hd__o211a_1 _15856_ (.A1(\jtag.dataIDRegister.data[0] ),
    .A2(net1171),
    .B1(_02926_),
    .C1(net1859),
    .X(_00903_));
 sky130_fd_sc_hd__and3_1 _15857_ (.A(net253),
    .B(net1309),
    .C(net1163),
    .X(_02927_));
 sky130_fd_sc_hd__a21o_1 _15858_ (.A1(\jtag.dataIDRegister.data[0] ),
    .A2(_02924_),
    .B1(net1167),
    .X(_02928_));
 sky130_fd_sc_hd__o221a_1 _15859_ (.A1(\jtag.dataIDRegister.data[1] ),
    .A2(net1171),
    .B1(_02927_),
    .B2(_02928_),
    .C1(net1859),
    .X(_00904_));
 sky130_fd_sc_hd__and3_1 _15860_ (.A(net255),
    .B(net1306),
    .C(net1163),
    .X(_02929_));
 sky130_fd_sc_hd__a21o_1 _15861_ (.A1(\jtag.dataIDRegister.data[1] ),
    .A2(_02924_),
    .B1(net1167),
    .X(_02930_));
 sky130_fd_sc_hd__o221a_1 _15862_ (.A1(\jtag.dataIDRegister.data[2] ),
    .A2(net1171),
    .B1(_02929_),
    .B2(_02930_),
    .C1(net1862),
    .X(_00905_));
 sky130_fd_sc_hd__and3_1 _15863_ (.A(net256),
    .B(net1306),
    .C(net1164),
    .X(_02931_));
 sky130_fd_sc_hd__a21o_1 _15864_ (.A1(\jtag.dataIDRegister.data[2] ),
    .A2(_02924_),
    .B1(net1167),
    .X(_02932_));
 sky130_fd_sc_hd__o221a_1 _15865_ (.A1(\jtag.dataIDRegister.data[3] ),
    .A2(net1172),
    .B1(_02931_),
    .B2(_02932_),
    .C1(net1862),
    .X(_00906_));
 sky130_fd_sc_hd__and3_1 _15866_ (.A(net257),
    .B(net1308),
    .C(net1164),
    .X(_02933_));
 sky130_fd_sc_hd__a21o_1 _15867_ (.A1(\jtag.dataIDRegister.data[3] ),
    .A2(_02924_),
    .B1(net1167),
    .X(_02934_));
 sky130_fd_sc_hd__o221a_1 _15868_ (.A1(\jtag.dataIDRegister.data[4] ),
    .A2(net1172),
    .B1(_02933_),
    .B2(_02934_),
    .C1(net1862),
    .X(_00907_));
 sky130_fd_sc_hd__and3_1 _15869_ (.A(net258),
    .B(net1306),
    .C(net1163),
    .X(_02935_));
 sky130_fd_sc_hd__a21o_1 _15870_ (.A1(\jtag.dataIDRegister.data[4] ),
    .A2(_02924_),
    .B1(net1168),
    .X(_02936_));
 sky130_fd_sc_hd__o221a_1 _15871_ (.A1(\jtag.dataIDRegister.data[5] ),
    .A2(net1171),
    .B1(_02935_),
    .B2(_02936_),
    .C1(net1862),
    .X(_00908_));
 sky130_fd_sc_hd__and3_1 _15872_ (.A(net259),
    .B(net1309),
    .C(net1163),
    .X(_02937_));
 sky130_fd_sc_hd__a21o_1 _15873_ (.A1(\jtag.dataIDRegister.data[5] ),
    .A2(_02924_),
    .B1(net1167),
    .X(_02938_));
 sky130_fd_sc_hd__o221a_1 _15874_ (.A1(\jtag.dataIDRegister.data[6] ),
    .A2(net1171),
    .B1(_02937_),
    .B2(_02938_),
    .C1(net1861),
    .X(_00909_));
 sky130_fd_sc_hd__and3_1 _15875_ (.A(net260),
    .B(net1306),
    .C(net1163),
    .X(_02939_));
 sky130_fd_sc_hd__a21o_1 _15876_ (.A1(\jtag.dataIDRegister.data[6] ),
    .A2(_02924_),
    .B1(net1167),
    .X(_02940_));
 sky130_fd_sc_hd__o221a_1 _15877_ (.A1(\jtag.dataIDRegister.data[7] ),
    .A2(net1171),
    .B1(_02939_),
    .B2(_02940_),
    .C1(net1861),
    .X(_00910_));
 sky130_fd_sc_hd__nand2b_1 _15878_ (.A_N(net261),
    .B(net1309),
    .Y(_02941_));
 sky130_fd_sc_hd__a221o_1 _15879_ (.A1(\jtag.dataIDRegister.data[7] ),
    .A2(net1282),
    .B1(net1163),
    .B2(_02941_),
    .C1(net1167),
    .X(_02942_));
 sky130_fd_sc_hd__o211a_1 _15880_ (.A1(\jtag.dataIDRegister.data[8] ),
    .A2(net1171),
    .B1(_02942_),
    .C1(net1861),
    .X(_00911_));
 sky130_fd_sc_hd__and3_1 _15881_ (.A(net262),
    .B(net1309),
    .C(net1163),
    .X(_02943_));
 sky130_fd_sc_hd__a211o_1 _15882_ (.A1(\jtag.dataIDRegister.data[8] ),
    .A2(net1282),
    .B1(net1167),
    .C1(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__o211a_1 _15883_ (.A1(\jtag.dataIDRegister.data[9] ),
    .A2(net1171),
    .B1(_02944_),
    .C1(net1861),
    .X(_00912_));
 sky130_fd_sc_hd__and3_1 _15884_ (.A(net263),
    .B(net1306),
    .C(net1163),
    .X(_02945_));
 sky130_fd_sc_hd__a211o_1 _15885_ (.A1(\jtag.dataIDRegister.data[9] ),
    .A2(net1282),
    .B1(net1170),
    .C1(_02945_),
    .X(_02946_));
 sky130_fd_sc_hd__o211a_1 _15886_ (.A1(\jtag.dataIDRegister.data[10] ),
    .A2(net1171),
    .B1(_02946_),
    .C1(net1861),
    .X(_00913_));
 sky130_fd_sc_hd__and3_1 _15887_ (.A(net254),
    .B(net1306),
    .C(net1165),
    .X(_02947_));
 sky130_fd_sc_hd__a211o_1 _15888_ (.A1(\jtag.dataIDRegister.data[10] ),
    .A2(net1282),
    .B1(net1169),
    .C1(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__o211a_1 _15889_ (.A1(\jtag.dataIDRegister.data[11] ),
    .A2(net1172),
    .B1(_02948_),
    .C1(net1861),
    .X(_00914_));
 sky130_fd_sc_hd__and3_1 _15890_ (.A(net264),
    .B(net1306),
    .C(net1164),
    .X(_02949_));
 sky130_fd_sc_hd__a211o_1 _15891_ (.A1(\jtag.dataIDRegister.data[11] ),
    .A2(net1282),
    .B1(net1168),
    .C1(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__o211a_1 _15892_ (.A1(\jtag.dataIDRegister.data[12] ),
    .A2(net1172),
    .B1(_02950_),
    .C1(net1861),
    .X(_00915_));
 sky130_fd_sc_hd__and3_1 _15893_ (.A(net271),
    .B(net1306),
    .C(net1164),
    .X(_02951_));
 sky130_fd_sc_hd__a211o_1 _15894_ (.A1(\jtag.dataIDRegister.data[12] ),
    .A2(net1282),
    .B1(net1168),
    .C1(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__o211a_1 _15895_ (.A1(\jtag.dataIDRegister.data[13] ),
    .A2(net1172),
    .B1(_02952_),
    .C1(net1861),
    .X(_00916_));
 sky130_fd_sc_hd__nand2b_1 _15896_ (.A_N(net272),
    .B(net1308),
    .Y(_02953_));
 sky130_fd_sc_hd__a221o_1 _15897_ (.A1(\jtag.dataIDRegister.data[13] ),
    .A2(net1282),
    .B1(net1164),
    .B2(_02953_),
    .C1(net1168),
    .X(_02954_));
 sky130_fd_sc_hd__o211a_1 _15898_ (.A1(\jtag.dataIDRegister.data[14] ),
    .A2(net1172),
    .B1(_02954_),
    .C1(net1862),
    .X(_00917_));
 sky130_fd_sc_hd__and3_1 _15899_ (.A(net273),
    .B(net1308),
    .C(net1164),
    .X(_02955_));
 sky130_fd_sc_hd__a211o_1 _15900_ (.A1(\jtag.dataIDRegister.data[14] ),
    .A2(net1282),
    .B1(net1168),
    .C1(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__o211a_1 _15901_ (.A1(\jtag.dataIDRegister.data[15] ),
    .A2(net1172),
    .B1(_02956_),
    .C1(net1861),
    .X(_00918_));
 sky130_fd_sc_hd__and3_1 _15902_ (.A(net274),
    .B(net1306),
    .C(net1164),
    .X(_02957_));
 sky130_fd_sc_hd__a211o_1 _15903_ (.A1(\jtag.dataIDRegister.data[15] ),
    .A2(net1282),
    .B1(net1168),
    .C1(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__o211a_1 _15904_ (.A1(\jtag.dataIDRegister.data[16] ),
    .A2(net1172),
    .B1(_02958_),
    .C1(net1861),
    .X(_00919_));
 sky130_fd_sc_hd__and3_1 _15905_ (.A(net275),
    .B(net1306),
    .C(net1164),
    .X(_02959_));
 sky130_fd_sc_hd__a211o_1 _15906_ (.A1(\jtag.dataIDRegister.data[16] ),
    .A2(net1282),
    .B1(net1167),
    .C1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__o211a_1 _15907_ (.A1(\jtag.dataIDRegister.data[17] ),
    .A2(net1172),
    .B1(_02960_),
    .C1(net1862),
    .X(_00920_));
 sky130_fd_sc_hd__and3_1 _15908_ (.A(net276),
    .B(net1308),
    .C(net1163),
    .X(_02961_));
 sky130_fd_sc_hd__a211o_1 _15909_ (.A1(\jtag.dataIDRegister.data[17] ),
    .A2(net1284),
    .B1(net1169),
    .C1(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__o211a_1 _15910_ (.A1(\jtag.dataIDRegister.data[18] ),
    .A2(net1172),
    .B1(_02962_),
    .C1(net1862),
    .X(_00921_));
 sky130_fd_sc_hd__and3_1 _15911_ (.A(net277),
    .B(net1307),
    .C(net1165),
    .X(_02963_));
 sky130_fd_sc_hd__a211o_1 _15912_ (.A1(\jtag.dataIDRegister.data[18] ),
    .A2(net1284),
    .B1(net1169),
    .C1(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__o211a_1 _15913_ (.A1(\jtag.dataIDRegister.data[19] ),
    .A2(net1173),
    .B1(_02964_),
    .C1(net1867),
    .X(_00922_));
 sky130_fd_sc_hd__and3_1 _15914_ (.A(net278),
    .B(net1307),
    .C(net1165),
    .X(_02965_));
 sky130_fd_sc_hd__a211o_1 _15915_ (.A1(\jtag.dataIDRegister.data[19] ),
    .A2(net1284),
    .B1(net1169),
    .C1(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__o211a_1 _15916_ (.A1(\jtag.dataIDRegister.data[20] ),
    .A2(net1173),
    .B1(_02966_),
    .C1(net1866),
    .X(_00923_));
 sky130_fd_sc_hd__and3_1 _15917_ (.A(net279),
    .B(net1308),
    .C(net1165),
    .X(_02967_));
 sky130_fd_sc_hd__a211o_1 _15918_ (.A1(\jtag.dataIDRegister.data[20] ),
    .A2(net1284),
    .B1(net1170),
    .C1(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__o211a_1 _15919_ (.A1(\jtag.dataIDRegister.data[21] ),
    .A2(net1173),
    .B1(_02968_),
    .C1(net1866),
    .X(_00924_));
 sky130_fd_sc_hd__and3_1 _15920_ (.A(net265),
    .B(net1307),
    .C(net1165),
    .X(_02969_));
 sky130_fd_sc_hd__a211o_1 _15921_ (.A1(\jtag.dataIDRegister.data[21] ),
    .A2(net1283),
    .B1(net1170),
    .C1(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__o211a_1 _15922_ (.A1(\jtag.dataIDRegister.data[22] ),
    .A2(net1173),
    .B1(_02970_),
    .C1(net1866),
    .X(_00925_));
 sky130_fd_sc_hd__and3_1 _15923_ (.A(net266),
    .B(net1308),
    .C(net1165),
    .X(_02971_));
 sky130_fd_sc_hd__a211o_1 _15924_ (.A1(\jtag.dataIDRegister.data[22] ),
    .A2(net1283),
    .B1(net1169),
    .C1(_02971_),
    .X(_02972_));
 sky130_fd_sc_hd__o211a_1 _15925_ (.A1(\jtag.dataIDRegister.data[23] ),
    .A2(net1173),
    .B1(_02972_),
    .C1(net1866),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _15926_ (.A0(net1),
    .A1(net267),
    .S(net1307),
    .X(_02973_));
 sky130_fd_sc_hd__a221o_1 _15927_ (.A1(\jtag.dataIDRegister.data[23] ),
    .A2(net1283),
    .B1(net1165),
    .B2(_02973_),
    .C1(net1169),
    .X(_02974_));
 sky130_fd_sc_hd__o211a_1 _15928_ (.A1(\jtag.dataIDRegister.data[24] ),
    .A2(net1173),
    .B1(_02974_),
    .C1(net1866),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _15929_ (.A0(net2),
    .A1(net268),
    .S(net1307),
    .X(_02975_));
 sky130_fd_sc_hd__a221o_1 _15930_ (.A1(\jtag.dataIDRegister.data[24] ),
    .A2(net1283),
    .B1(net1165),
    .B2(_02975_),
    .C1(net1169),
    .X(_02976_));
 sky130_fd_sc_hd__o211a_1 _15931_ (.A1(\jtag.dataIDRegister.data[25] ),
    .A2(net1173),
    .B1(_02976_),
    .C1(net1867),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _15932_ (.A0(net3),
    .A1(net269),
    .S(net1307),
    .X(_02977_));
 sky130_fd_sc_hd__a221o_1 _15933_ (.A1(\jtag.dataIDRegister.data[25] ),
    .A2(net1283),
    .B1(net1165),
    .B2(_02977_),
    .C1(net1169),
    .X(_02978_));
 sky130_fd_sc_hd__o211a_1 _15934_ (.A1(\jtag.dataIDRegister.data[26] ),
    .A2(net1173),
    .B1(_02978_),
    .C1(net1866),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _15935_ (.A0(net4),
    .A1(net270),
    .S(net1307),
    .X(_02979_));
 sky130_fd_sc_hd__a221o_1 _15936_ (.A1(\jtag.dataIDRegister.data[26] ),
    .A2(net1283),
    .B1(net1166),
    .B2(_02979_),
    .C1(net1169),
    .X(_02980_));
 sky130_fd_sc_hd__o211a_1 _15937_ (.A1(\jtag.dataIDRegister.data[27] ),
    .A2(net1173),
    .B1(_02980_),
    .C1(net1866),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _15938_ (.A0(net5),
    .A1(net280),
    .S(net1307),
    .X(_02981_));
 sky130_fd_sc_hd__a221o_1 _15939_ (.A1(\jtag.dataIDRegister.data[27] ),
    .A2(net1283),
    .B1(net1166),
    .B2(_02981_),
    .C1(net1170),
    .X(_02982_));
 sky130_fd_sc_hd__o211a_1 _15940_ (.A1(\jtag.dataIDRegister.data[28] ),
    .A2(net1174),
    .B1(_02982_),
    .C1(net1866),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _15941_ (.A0(net6),
    .A1(net281),
    .S(net1308),
    .X(_02983_));
 sky130_fd_sc_hd__a221o_1 _15942_ (.A1(\jtag.dataIDRegister.data[28] ),
    .A2(net1283),
    .B1(net1166),
    .B2(_02983_),
    .C1(net1170),
    .X(_02984_));
 sky130_fd_sc_hd__o211a_1 _15943_ (.A1(\jtag.dataIDRegister.data[29] ),
    .A2(net1173),
    .B1(_02984_),
    .C1(net1866),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _15944_ (.A0(net7),
    .A1(net282),
    .S(net1307),
    .X(_02985_));
 sky130_fd_sc_hd__a221o_1 _15945_ (.A1(\jtag.dataIDRegister.data[29] ),
    .A2(net1283),
    .B1(net1165),
    .B2(_02985_),
    .C1(net1169),
    .X(_02986_));
 sky130_fd_sc_hd__o211a_1 _15946_ (.A1(\jtag.dataIDRegister.data[30] ),
    .A2(net1174),
    .B1(_02986_),
    .C1(net1866),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _15947_ (.A0(net8),
    .A1(net283),
    .S(net1307),
    .X(_02987_));
 sky130_fd_sc_hd__a221o_1 _15948_ (.A1(\jtag.dataIDRegister.data[30] ),
    .A2(net1283),
    .B1(net1166),
    .B2(_02987_),
    .C1(net1170),
    .X(_02988_));
 sky130_fd_sc_hd__o211a_1 _15949_ (.A1(\jtag.dataIDRegister.data[31] ),
    .A2(net1171),
    .B1(_02988_),
    .C1(net1859),
    .X(_00934_));
 sky130_fd_sc_hd__a31o_1 _15950_ (.A1(net1723),
    .A2(_06841_),
    .A3(_06847_),
    .B1(\jtag.dataBypassRegister.data ),
    .X(_02989_));
 sky130_fd_sc_hd__a41o_1 _15951_ (.A1(net1723),
    .A2(_06841_),
    .A3(_02920_),
    .A4(_02925_),
    .B1(net1874),
    .X(_02990_));
 sky130_fd_sc_hd__and2b_1 _15952_ (.A_N(_02990_),
    .B(_02989_),
    .X(_00935_));
 sky130_fd_sc_hd__nor2_1 _15953_ (.A(_08703_),
    .B(net1280),
    .Y(_02991_));
 sky130_fd_sc_hd__and3_1 _15954_ (.A(\jtag.tckRisingEdge ),
    .B(_06844_),
    .C(_02920_),
    .X(_02992_));
 sky130_fd_sc_hd__nand2b_1 _15955_ (.A_N(_08703_),
    .B(_02920_),
    .Y(_02993_));
 sky130_fd_sc_hd__a221o_1 _15956_ (.A1(net188),
    .A2(net1286),
    .B1(net1190),
    .B2(\jtag.managementReadData[0] ),
    .C1(net1155),
    .X(_02994_));
 sky130_fd_sc_hd__o211a_1 _15957_ (.A1(\jtag.dataBSRRegister.data[0] ),
    .A2(net1159),
    .B1(_02994_),
    .C1(net1842),
    .X(_00936_));
 sky130_fd_sc_hd__a221o_1 _15958_ (.A1(\jtag.dataBSRRegister.data[0] ),
    .A2(net1286),
    .B1(net1190),
    .B2(\jtag.managementReadData[1] ),
    .C1(net1155),
    .X(_02995_));
 sky130_fd_sc_hd__o211a_1 _15959_ (.A1(\jtag.dataBSRRegister.data[1] ),
    .A2(net1159),
    .B1(_02995_),
    .C1(net1852),
    .X(_00937_));
 sky130_fd_sc_hd__a221o_1 _15960_ (.A1(\jtag.dataBSRRegister.data[1] ),
    .A2(net1286),
    .B1(net1190),
    .B2(\jtag.managementReadData[2] ),
    .C1(net1155),
    .X(_02996_));
 sky130_fd_sc_hd__o211a_1 _15961_ (.A1(\jtag.dataBSRRegister.data[2] ),
    .A2(net1159),
    .B1(_02996_),
    .C1(net1852),
    .X(_00938_));
 sky130_fd_sc_hd__a221o_1 _15962_ (.A1(\jtag.dataBSRRegister.data[2] ),
    .A2(net1286),
    .B1(net1190),
    .B2(\jtag.managementReadData[3] ),
    .C1(net1155),
    .X(_02997_));
 sky130_fd_sc_hd__o211a_1 _15963_ (.A1(\jtag.dataBSRRegister.data[3] ),
    .A2(net1159),
    .B1(_02997_),
    .C1(net1852),
    .X(_00939_));
 sky130_fd_sc_hd__a221o_1 _15964_ (.A1(\jtag.dataBSRRegister.data[3] ),
    .A2(net1286),
    .B1(net1190),
    .B2(\jtag.managementReadData[4] ),
    .C1(net1155),
    .X(_02998_));
 sky130_fd_sc_hd__o211a_1 _15965_ (.A1(\jtag.dataBSRRegister.data[4] ),
    .A2(net1159),
    .B1(_02998_),
    .C1(net1850),
    .X(_00940_));
 sky130_fd_sc_hd__a221o_1 _15966_ (.A1(\jtag.dataBSRRegister.data[4] ),
    .A2(net1286),
    .B1(net1190),
    .B2(\jtag.managementReadData[5] ),
    .C1(net1155),
    .X(_02999_));
 sky130_fd_sc_hd__o211a_1 _15967_ (.A1(\jtag.dataBSRRegister.data[5] ),
    .A2(net1159),
    .B1(_02999_),
    .C1(net1839),
    .X(_00941_));
 sky130_fd_sc_hd__a221o_1 _15968_ (.A1(\jtag.dataBSRRegister.data[5] ),
    .A2(net1286),
    .B1(net1190),
    .B2(\jtag.managementReadData[6] ),
    .C1(net1155),
    .X(_03000_));
 sky130_fd_sc_hd__o211a_1 _15969_ (.A1(\jtag.dataBSRRegister.data[6] ),
    .A2(net1159),
    .B1(_03000_),
    .C1(net1839),
    .X(_00942_));
 sky130_fd_sc_hd__a221o_1 _15970_ (.A1(\jtag.dataBSRRegister.data[6] ),
    .A2(net1286),
    .B1(net1190),
    .B2(\jtag.managementReadData[7] ),
    .C1(net1155),
    .X(_03001_));
 sky130_fd_sc_hd__o211a_1 _15971_ (.A1(\jtag.dataBSRRegister.data[7] ),
    .A2(net1159),
    .B1(_03001_),
    .C1(net1842),
    .X(_00943_));
 sky130_fd_sc_hd__a221o_1 _15972_ (.A1(\jtag.dataBSRRegister.data[7] ),
    .A2(net1280),
    .B1(net1190),
    .B2(\jtag.managementReadData[8] ),
    .C1(net1155),
    .X(_03002_));
 sky130_fd_sc_hd__o211a_1 _15973_ (.A1(\jtag.dataBSRRegister.data[8] ),
    .A2(net1159),
    .B1(_03002_),
    .C1(net1856),
    .X(_00944_));
 sky130_fd_sc_hd__a221o_1 _15974_ (.A1(\jtag.dataBSRRegister.data[8] ),
    .A2(net1280),
    .B1(net1193),
    .B2(\jtag.managementReadData[9] ),
    .C1(net1158),
    .X(_03003_));
 sky130_fd_sc_hd__o211a_1 _15975_ (.A1(\jtag.dataBSRRegister.data[9] ),
    .A2(net1162),
    .B1(_03003_),
    .C1(net1864),
    .X(_00945_));
 sky130_fd_sc_hd__a221o_1 _15976_ (.A1(\jtag.dataBSRRegister.data[9] ),
    .A2(net1280),
    .B1(net1190),
    .B2(\jtag.managementReadData[10] ),
    .C1(net1155),
    .X(_03004_));
 sky130_fd_sc_hd__o211a_1 _15977_ (.A1(\jtag.dataBSRRegister.data[10] ),
    .A2(net1159),
    .B1(_03004_),
    .C1(net1864),
    .X(_00946_));
 sky130_fd_sc_hd__a221o_1 _15978_ (.A1(\jtag.dataBSRRegister.data[10] ),
    .A2(net1280),
    .B1(net1192),
    .B2(\jtag.managementReadData[11] ),
    .C1(net1156),
    .X(_03005_));
 sky130_fd_sc_hd__o211a_1 _15979_ (.A1(\jtag.dataBSRRegister.data[11] ),
    .A2(net1160),
    .B1(_03005_),
    .C1(net1864),
    .X(_00947_));
 sky130_fd_sc_hd__a221o_1 _15980_ (.A1(\jtag.dataBSRRegister.data[11] ),
    .A2(net1280),
    .B1(net1192),
    .B2(\jtag.managementReadData[12] ),
    .C1(net1157),
    .X(_03006_));
 sky130_fd_sc_hd__o211a_1 _15981_ (.A1(\jtag.dataBSRRegister.data[12] ),
    .A2(net1160),
    .B1(_03006_),
    .C1(net1865),
    .X(_00948_));
 sky130_fd_sc_hd__a221o_1 _15982_ (.A1(\jtag.dataBSRRegister.data[12] ),
    .A2(net1281),
    .B1(net1191),
    .B2(\jtag.managementReadData[13] ),
    .C1(net1156),
    .X(_03007_));
 sky130_fd_sc_hd__o211a_1 _15983_ (.A1(\jtag.dataBSRRegister.data[13] ),
    .A2(net1161),
    .B1(_03007_),
    .C1(net1864),
    .X(_00949_));
 sky130_fd_sc_hd__a221o_1 _15984_ (.A1(\jtag.dataBSRRegister.data[13] ),
    .A2(net1281),
    .B1(net1191),
    .B2(\jtag.managementReadData[14] ),
    .C1(net1156),
    .X(_03008_));
 sky130_fd_sc_hd__o211a_1 _15985_ (.A1(\jtag.dataBSRRegister.data[14] ),
    .A2(net1160),
    .B1(_03008_),
    .C1(net1857),
    .X(_00950_));
 sky130_fd_sc_hd__a221o_1 _15986_ (.A1(\jtag.dataBSRRegister.data[14] ),
    .A2(net1281),
    .B1(net1192),
    .B2(\jtag.managementReadData[15] ),
    .C1(net1157),
    .X(_03009_));
 sky130_fd_sc_hd__o211a_1 _15987_ (.A1(\jtag.dataBSRRegister.data[15] ),
    .A2(net1161),
    .B1(_03009_),
    .C1(net1857),
    .X(_00951_));
 sky130_fd_sc_hd__a221o_1 _15988_ (.A1(\jtag.dataBSRRegister.data[15] ),
    .A2(net1281),
    .B1(net1192),
    .B2(\jtag.managementReadData[16] ),
    .C1(net1157),
    .X(_03010_));
 sky130_fd_sc_hd__o211a_1 _15989_ (.A1(\jtag.dataBSRRegister.data[16] ),
    .A2(net1161),
    .B1(_03010_),
    .C1(net1860),
    .X(_00952_));
 sky130_fd_sc_hd__a221o_1 _15990_ (.A1(\jtag.dataBSRRegister.data[16] ),
    .A2(net1285),
    .B1(net1192),
    .B2(\jtag.managementReadData[17] ),
    .C1(net1157),
    .X(_03011_));
 sky130_fd_sc_hd__o211a_1 _15991_ (.A1(\jtag.dataBSRRegister.data[17] ),
    .A2(net1161),
    .B1(_03011_),
    .C1(net1859),
    .X(_00953_));
 sky130_fd_sc_hd__a221o_1 _15992_ (.A1(\jtag.dataBSRRegister.data[17] ),
    .A2(net1285),
    .B1(net1192),
    .B2(\jtag.managementReadData[18] ),
    .C1(net1157),
    .X(_03012_));
 sky130_fd_sc_hd__o211a_1 _15993_ (.A1(\jtag.dataBSRRegister.data[18] ),
    .A2(net1161),
    .B1(_03012_),
    .C1(net1859),
    .X(_00954_));
 sky130_fd_sc_hd__a221o_1 _15994_ (.A1(\jtag.dataBSRRegister.data[18] ),
    .A2(net1285),
    .B1(net1193),
    .B2(\jtag.managementReadData[19] ),
    .C1(net1158),
    .X(_03013_));
 sky130_fd_sc_hd__o211a_1 _15995_ (.A1(\jtag.dataBSRRegister.data[19] ),
    .A2(net1162),
    .B1(_03013_),
    .C1(net1860),
    .X(_00955_));
 sky130_fd_sc_hd__a221o_1 _15996_ (.A1(\jtag.dataBSRRegister.data[19] ),
    .A2(net1285),
    .B1(net1192),
    .B2(\jtag.managementReadData[20] ),
    .C1(net1157),
    .X(_03014_));
 sky130_fd_sc_hd__o211a_1 _15997_ (.A1(\jtag.dataBSRRegister.data[20] ),
    .A2(net1161),
    .B1(_03014_),
    .C1(net1859),
    .X(_00956_));
 sky130_fd_sc_hd__a221o_1 _15998_ (.A1(\jtag.dataBSRRegister.data[20] ),
    .A2(net1285),
    .B1(net1192),
    .B2(\jtag.managementReadData[21] ),
    .C1(net1157),
    .X(_03015_));
 sky130_fd_sc_hd__o211a_1 _15999_ (.A1(\jtag.dataBSRRegister.data[21] ),
    .A2(net1161),
    .B1(_03015_),
    .C1(net1859),
    .X(_00957_));
 sky130_fd_sc_hd__a221o_1 _16000_ (.A1(\jtag.dataBSRRegister.data[21] ),
    .A2(net1285),
    .B1(net1193),
    .B2(\jtag.managementReadData[22] ),
    .C1(net1157),
    .X(_03016_));
 sky130_fd_sc_hd__o211a_1 _16001_ (.A1(\jtag.dataBSRRegister.data[22] ),
    .A2(net1161),
    .B1(_03016_),
    .C1(net1859),
    .X(_00958_));
 sky130_fd_sc_hd__a221o_1 _16002_ (.A1(\jtag.dataBSRRegister.data[22] ),
    .A2(net1285),
    .B1(net1193),
    .B2(\jtag.managementReadData[23] ),
    .C1(net1158),
    .X(_03017_));
 sky130_fd_sc_hd__o211a_1 _16003_ (.A1(\jtag.dataBSRRegister.data[23] ),
    .A2(net1162),
    .B1(_03017_),
    .C1(net1859),
    .X(_00959_));
 sky130_fd_sc_hd__a221o_1 _16004_ (.A1(\jtag.dataBSRRegister.data[23] ),
    .A2(net1281),
    .B1(net1192),
    .B2(\jtag.managementReadData[24] ),
    .C1(net1157),
    .X(_03018_));
 sky130_fd_sc_hd__o211a_1 _16005_ (.A1(\jtag.dataBSRRegister.data[24] ),
    .A2(net1161),
    .B1(_03018_),
    .C1(net1857),
    .X(_00960_));
 sky130_fd_sc_hd__a221o_1 _16006_ (.A1(\jtag.dataBSRRegister.data[24] ),
    .A2(net1281),
    .B1(net1191),
    .B2(\jtag.managementReadData[25] ),
    .C1(net1156),
    .X(_03019_));
 sky130_fd_sc_hd__o211a_1 _16007_ (.A1(\jtag.dataBSRRegister.data[25] ),
    .A2(net1160),
    .B1(_03019_),
    .C1(net1857),
    .X(_00961_));
 sky130_fd_sc_hd__a221o_1 _16008_ (.A1(\jtag.dataBSRRegister.data[25] ),
    .A2(net1280),
    .B1(net1191),
    .B2(\jtag.managementReadData[26] ),
    .C1(net1156),
    .X(_03020_));
 sky130_fd_sc_hd__o211a_1 _16009_ (.A1(\jtag.dataBSRRegister.data[26] ),
    .A2(net1160),
    .B1(_03020_),
    .C1(net1856),
    .X(_00962_));
 sky130_fd_sc_hd__a221o_1 _16010_ (.A1(\jtag.dataBSRRegister.data[26] ),
    .A2(net1280),
    .B1(net1191),
    .B2(\jtag.managementReadData[27] ),
    .C1(net1156),
    .X(_03021_));
 sky130_fd_sc_hd__o211a_1 _16011_ (.A1(\jtag.dataBSRRegister.data[27] ),
    .A2(net1160),
    .B1(_03021_),
    .C1(net1856),
    .X(_00963_));
 sky130_fd_sc_hd__a221o_1 _16012_ (.A1(\jtag.dataBSRRegister.data[27] ),
    .A2(net1280),
    .B1(net1191),
    .B2(\jtag.managementReadData[28] ),
    .C1(net1156),
    .X(_03022_));
 sky130_fd_sc_hd__o211a_1 _16013_ (.A1(\jtag.dataBSRRegister.data[28] ),
    .A2(net1160),
    .B1(_03022_),
    .C1(net1857),
    .X(_00964_));
 sky130_fd_sc_hd__a221o_1 _16014_ (.A1(\jtag.dataBSRRegister.data[28] ),
    .A2(net1281),
    .B1(net1191),
    .B2(\jtag.managementReadData[29] ),
    .C1(net1156),
    .X(_03023_));
 sky130_fd_sc_hd__o211a_1 _16015_ (.A1(\jtag.dataBSRRegister.data[29] ),
    .A2(net1160),
    .B1(_03023_),
    .C1(net1857),
    .X(_00965_));
 sky130_fd_sc_hd__a221o_1 _16016_ (.A1(\jtag.dataBSRRegister.data[29] ),
    .A2(net1281),
    .B1(net1191),
    .B2(\jtag.managementReadData[30] ),
    .C1(net1156),
    .X(_03024_));
 sky130_fd_sc_hd__o211a_1 _16017_ (.A1(\jtag.dataBSRRegister.data[30] ),
    .A2(net1160),
    .B1(_03024_),
    .C1(net1857),
    .X(_00966_));
 sky130_fd_sc_hd__a221o_1 _16018_ (.A1(\jtag.dataBSRRegister.data[30] ),
    .A2(net1280),
    .B1(net1191),
    .B2(\jtag.managementReadData[31] ),
    .C1(net1156),
    .X(_03025_));
 sky130_fd_sc_hd__o211a_1 _16019_ (.A1(\jtag.dataBSRRegister.data[31] ),
    .A2(net1160),
    .B1(_03025_),
    .C1(net1857),
    .X(_00967_));
 sky130_fd_sc_hd__nand2_2 _16020_ (.A(net1722),
    .B(_06835_),
    .Y(_03026_));
 sky130_fd_sc_hd__a21o_1 _16021_ (.A1(net1722),
    .A2(_06835_),
    .B1(\jtag.instructionRegister.data[0] ),
    .X(_03027_));
 sky130_fd_sc_hd__mux2_1 _16022_ (.A0(net445),
    .A1(net188),
    .S(net1721),
    .X(_03028_));
 sky130_fd_sc_hd__o211a_1 _16023_ (.A1(_03026_),
    .A2(_03028_),
    .B1(_03027_),
    .C1(net1803),
    .X(_00968_));
 sky130_fd_sc_hd__a21o_1 _16024_ (.A1(net1722),
    .A2(_06835_),
    .B1(\jtag.instructionRegister.data[1] ),
    .X(_03029_));
 sky130_fd_sc_hd__mux2_1 _16025_ (.A0(net446),
    .A1(\jtag.instructionRegister.data[0] ),
    .S(net1721),
    .X(_03030_));
 sky130_fd_sc_hd__o211a_1 _16026_ (.A1(_03026_),
    .A2(_03030_),
    .B1(_03029_),
    .C1(net1803),
    .X(_00969_));
 sky130_fd_sc_hd__a21o_1 _16027_ (.A1(net1722),
    .A2(_06835_),
    .B1(\jtag.instructionRegister.data[2] ),
    .X(_03031_));
 sky130_fd_sc_hd__mux2_1 _16028_ (.A0(net447),
    .A1(\jtag.instructionRegister.data[1] ),
    .S(net1721),
    .X(_03032_));
 sky130_fd_sc_hd__o211a_1 _16029_ (.A1(_03026_),
    .A2(_03032_),
    .B1(_03031_),
    .C1(net1803),
    .X(_00970_));
 sky130_fd_sc_hd__a21o_1 _16030_ (.A1(net1722),
    .A2(_06835_),
    .B1(\jtag.instructionRegister.data[3] ),
    .X(_03033_));
 sky130_fd_sc_hd__mux2_1 _16031_ (.A0(net448),
    .A1(\jtag.instructionRegister.data[2] ),
    .S(net1721),
    .X(_03034_));
 sky130_fd_sc_hd__o211a_1 _16032_ (.A1(_03026_),
    .A2(_03034_),
    .B1(_03033_),
    .C1(net1803),
    .X(_00971_));
 sky130_fd_sc_hd__a21o_1 _16033_ (.A1(net1722),
    .A2(_06835_),
    .B1(\jtag.instructionRegister.data[4] ),
    .X(_03035_));
 sky130_fd_sc_hd__mux2_1 _16034_ (.A0(net449),
    .A1(\jtag.instructionRegister.data[3] ),
    .S(net1721),
    .X(_03036_));
 sky130_fd_sc_hd__o211a_1 _16035_ (.A1(_03026_),
    .A2(_03036_),
    .B1(_03035_),
    .C1(net1803),
    .X(_00972_));
 sky130_fd_sc_hd__o21ai_1 _16036_ (.A1(_03817_),
    .A2(net187),
    .B1(\jtag.tckState ),
    .Y(_03037_));
 sky130_fd_sc_hd__o211a_1 _16037_ (.A1(net187),
    .A2(\jtag.tckState ),
    .B1(net1802),
    .C1(_03037_),
    .X(_00973_));
 sky130_fd_sc_hd__and2_1 _16038_ (.A(net187),
    .B(net1802),
    .X(_00974_));
 sky130_fd_sc_hd__or3_2 _16039_ (.A(net1720),
    .B(\jtag.state[0] ),
    .C(_02917_),
    .X(_03038_));
 sky130_fd_sc_hd__nand2_2 _16040_ (.A(\jtag.state[3] ),
    .B(\jtag.state[2] ),
    .Y(_03039_));
 sky130_fd_sc_hd__or2_1 _16041_ (.A(_06834_),
    .B(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__a21o_4 _16042_ (.A1(_03038_),
    .A2(_03040_),
    .B1(_03817_),
    .X(_03041_));
 sky130_fd_sc_hd__mux2_1 _16043_ (.A0(\jtag.instructionRegister.data[0] ),
    .A1(net445),
    .S(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__and2_1 _16044_ (.A(net1802),
    .B(_03042_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _16045_ (.A0(\jtag.instructionRegister.data[1] ),
    .A1(net446),
    .S(_03041_),
    .X(_03043_));
 sky130_fd_sc_hd__and2_1 _16046_ (.A(net1802),
    .B(_03043_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _16047_ (.A0(\jtag.instructionRegister.data[2] ),
    .A1(net447),
    .S(_03041_),
    .X(_03044_));
 sky130_fd_sc_hd__or2_1 _16048_ (.A(net1874),
    .B(_03044_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _16049_ (.A0(\jtag.instructionRegister.data[3] ),
    .A1(net448),
    .S(_03041_),
    .X(_03045_));
 sky130_fd_sc_hd__and2_1 _16050_ (.A(net1803),
    .B(_03045_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _16051_ (.A0(\jtag.instructionRegister.data[4] ),
    .A1(net449),
    .S(_03041_),
    .X(_03046_));
 sky130_fd_sc_hd__and2_1 _16052_ (.A(net1803),
    .B(_03046_),
    .X(_00979_));
 sky130_fd_sc_hd__o21ai_1 _16053_ (.A1(\jtag.state[0] ),
    .A2(_06846_),
    .B1(_02919_),
    .Y(_03047_));
 sky130_fd_sc_hd__or2_2 _16054_ (.A(net1720),
    .B(_03819_),
    .X(_03048_));
 sky130_fd_sc_hd__inv_2 _16055_ (.A(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__nor2_1 _16056_ (.A(net189),
    .B(_06835_),
    .Y(_03050_));
 sky130_fd_sc_hd__o211a_1 _16057_ (.A1(_02917_),
    .A2(_03048_),
    .B1(_03040_),
    .C1(_08702_),
    .X(_03051_));
 sky130_fd_sc_hd__o211a_1 _16058_ (.A1(_03039_),
    .A2(_03048_),
    .B1(_03051_),
    .C1(_03038_),
    .X(_03052_));
 sky130_fd_sc_hd__a2bb2o_1 _16059_ (.A1_N(_03853_),
    .A2_N(_03047_),
    .B1(_03050_),
    .B2(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__or3b_2 _16060_ (.A(\jtag.state[0] ),
    .B(_02917_),
    .C_N(\jtag.state[1] ),
    .X(_03054_));
 sky130_fd_sc_hd__o211a_1 _16061_ (.A1(net1721),
    .A2(_03039_),
    .B1(_03054_),
    .C1(net1722),
    .X(_03055_));
 sky130_fd_sc_hd__a221oi_1 _16062_ (.A1(_03817_),
    .A2(_03819_),
    .B1(_03053_),
    .B2(_03055_),
    .C1(net1874),
    .Y(_00980_));
 sky130_fd_sc_hd__nand3_1 _16063_ (.A(_02917_),
    .B(_03039_),
    .C(_03049_),
    .Y(_03056_));
 sky130_fd_sc_hd__o211a_1 _16064_ (.A1(net1720),
    .A2(_03039_),
    .B1(_03051_),
    .C1(net189),
    .X(_03057_));
 sky130_fd_sc_hd__a31oi_1 _16065_ (.A1(_03050_),
    .A2(_03054_),
    .A3(_03056_),
    .B1(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__a31o_1 _16066_ (.A1(\jtag.state[2] ),
    .A2(net1720),
    .A3(_03819_),
    .B1(_03817_),
    .X(_03059_));
 sky130_fd_sc_hd__o221a_1 _16067_ (.A1(net1722),
    .A2(net1720),
    .B1(_03058_),
    .B2(_03059_),
    .C1(net1804),
    .X(_00981_));
 sky130_fd_sc_hd__o211a_1 _16068_ (.A1(_03818_),
    .A2(_03819_),
    .B1(net1720),
    .C1(\jtag.state[3] ),
    .X(_03060_));
 sky130_fd_sc_hd__or2_1 _16069_ (.A(_03819_),
    .B(_06846_),
    .X(_03061_));
 sky130_fd_sc_hd__o21ai_1 _16070_ (.A1(net1720),
    .A2(_03039_),
    .B1(net1723),
    .Y(_03062_));
 sky130_fd_sc_hd__a211oi_1 _16071_ (.A1(net189),
    .A2(_03060_),
    .B1(_03062_),
    .C1(_03047_),
    .Y(_03063_));
 sky130_fd_sc_hd__o21ai_1 _16072_ (.A1(net189),
    .A2(_03061_),
    .B1(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__o211a_1 _16073_ (.A1(net1722),
    .A2(\jtag.state[2] ),
    .B1(net1804),
    .C1(_03064_),
    .X(_00982_));
 sky130_fd_sc_hd__a31o_1 _16074_ (.A1(\jtag.state[3] ),
    .A2(_03818_),
    .A3(_03049_),
    .B1(net189),
    .X(_03065_));
 sky130_fd_sc_hd__nand3_1 _16075_ (.A(net189),
    .B(_03054_),
    .C(_03061_),
    .Y(_03066_));
 sky130_fd_sc_hd__a21o_1 _16076_ (.A1(_03065_),
    .A2(_03066_),
    .B1(_03062_),
    .X(_03067_));
 sky130_fd_sc_hd__o221a_1 _16077_ (.A1(\jtag.state[3] ),
    .A2(net1722),
    .B1(_03060_),
    .B2(_03067_),
    .C1(net1804),
    .X(_00983_));
 sky130_fd_sc_hd__or3_4 _16078_ (.A(_03816_),
    .B(net1610),
    .C(_02103_),
    .X(_03068_));
 sky130_fd_sc_hd__nand2_1 _16079_ (.A(\jtag.managementReadData[0] ),
    .B(net1610),
    .Y(_03069_));
 sky130_fd_sc_hd__a21oi_1 _16080_ (.A1(net575),
    .A2(_03069_),
    .B1(net1886),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _16081_ (.A(\jtag.managementReadData[1] ),
    .B(net1610),
    .Y(_03070_));
 sky130_fd_sc_hd__a21oi_1 _16082_ (.A1(net575),
    .A2(_03070_),
    .B1(net1886),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_1 _16083_ (.A(\jtag.managementReadData[2] ),
    .B(net1610),
    .Y(_03071_));
 sky130_fd_sc_hd__a21oi_1 _16084_ (.A1(net575),
    .A2(_03071_),
    .B1(net1886),
    .Y(_00986_));
 sky130_fd_sc_hd__nand2_1 _16085_ (.A(\jtag.managementReadData[3] ),
    .B(net1610),
    .Y(_03072_));
 sky130_fd_sc_hd__a21oi_1 _16086_ (.A1(net575),
    .A2(_03072_),
    .B1(net1886),
    .Y(_00987_));
 sky130_fd_sc_hd__nand2_1 _16087_ (.A(\jtag.managementReadData[4] ),
    .B(net1610),
    .Y(_03073_));
 sky130_fd_sc_hd__a21oi_1 _16088_ (.A1(net575),
    .A2(_03073_),
    .B1(net1886),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _16089_ (.A(\jtag.managementReadData[5] ),
    .B(net1610),
    .Y(_03074_));
 sky130_fd_sc_hd__a21oi_1 _16090_ (.A1(net575),
    .A2(_03074_),
    .B1(net1886),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2_1 _16091_ (.A(\jtag.managementReadData[6] ),
    .B(net1610),
    .Y(_03075_));
 sky130_fd_sc_hd__a21oi_1 _16092_ (.A1(net575),
    .A2(_03075_),
    .B1(net1886),
    .Y(_00990_));
 sky130_fd_sc_hd__nand2_1 _16093_ (.A(\jtag.managementReadData[7] ),
    .B(net1610),
    .Y(_03076_));
 sky130_fd_sc_hd__a21oi_1 _16094_ (.A1(net575),
    .A2(_03076_),
    .B1(net1886),
    .Y(_00991_));
 sky130_fd_sc_hd__nand2_1 _16095_ (.A(\jtag.managementReadData[8] ),
    .B(_07009_),
    .Y(_03077_));
 sky130_fd_sc_hd__a21oi_1 _16096_ (.A1(net575),
    .A2(_03077_),
    .B1(net1887),
    .Y(_00992_));
 sky130_fd_sc_hd__nand2_1 _16097_ (.A(\jtag.managementReadData[9] ),
    .B(net1611),
    .Y(_03078_));
 sky130_fd_sc_hd__a21oi_1 _16098_ (.A1(net574),
    .A2(_03078_),
    .B1(net1887),
    .Y(_00993_));
 sky130_fd_sc_hd__nand2_1 _16099_ (.A(\jtag.managementReadData[10] ),
    .B(net1611),
    .Y(_03079_));
 sky130_fd_sc_hd__a21oi_1 _16100_ (.A1(net574),
    .A2(_03079_),
    .B1(net1887),
    .Y(_00994_));
 sky130_fd_sc_hd__nand2_1 _16101_ (.A(\jtag.managementReadData[11] ),
    .B(net1611),
    .Y(_03080_));
 sky130_fd_sc_hd__a21oi_1 _16102_ (.A1(net574),
    .A2(_03080_),
    .B1(net1887),
    .Y(_00995_));
 sky130_fd_sc_hd__nand2_1 _16103_ (.A(\jtag.managementReadData[12] ),
    .B(net1611),
    .Y(_03081_));
 sky130_fd_sc_hd__a21oi_1 _16104_ (.A1(net574),
    .A2(_03081_),
    .B1(net1887),
    .Y(_00996_));
 sky130_fd_sc_hd__nand2_1 _16105_ (.A(\jtag.managementReadData[13] ),
    .B(net1613),
    .Y(_03082_));
 sky130_fd_sc_hd__a21oi_1 _16106_ (.A1(net573),
    .A2(_03082_),
    .B1(net1887),
    .Y(_00997_));
 sky130_fd_sc_hd__nand2_1 _16107_ (.A(\jtag.managementReadData[14] ),
    .B(net1613),
    .Y(_03083_));
 sky130_fd_sc_hd__a21oi_1 _16108_ (.A1(net574),
    .A2(_03083_),
    .B1(net1887),
    .Y(_00998_));
 sky130_fd_sc_hd__nand2_1 _16109_ (.A(\jtag.managementReadData[15] ),
    .B(net1612),
    .Y(_03084_));
 sky130_fd_sc_hd__a21oi_1 _16110_ (.A1(_03068_),
    .A2(_03084_),
    .B1(net1904),
    .Y(_00999_));
 sky130_fd_sc_hd__nand2_1 _16111_ (.A(\jtag.managementReadData[16] ),
    .B(net1613),
    .Y(_03085_));
 sky130_fd_sc_hd__a21oi_1 _16112_ (.A1(_03068_),
    .A2(_03085_),
    .B1(net1889),
    .Y(_01000_));
 sky130_fd_sc_hd__nand2_1 _16113_ (.A(\jtag.managementReadData[17] ),
    .B(net1613),
    .Y(_03086_));
 sky130_fd_sc_hd__a21oi_1 _16114_ (.A1(_03068_),
    .A2(_03086_),
    .B1(net1889),
    .Y(_01001_));
 sky130_fd_sc_hd__nand2_1 _16115_ (.A(\jtag.managementReadData[18] ),
    .B(net1612),
    .Y(_03087_));
 sky130_fd_sc_hd__a21oi_1 _16116_ (.A1(net573),
    .A2(_03087_),
    .B1(net1888),
    .Y(_01002_));
 sky130_fd_sc_hd__nand2_1 _16117_ (.A(\jtag.managementReadData[19] ),
    .B(net1612),
    .Y(_03088_));
 sky130_fd_sc_hd__a21oi_1 _16118_ (.A1(net573),
    .A2(_03088_),
    .B1(net1889),
    .Y(_01003_));
 sky130_fd_sc_hd__nand2_1 _16119_ (.A(\jtag.managementReadData[20] ),
    .B(net1612),
    .Y(_03089_));
 sky130_fd_sc_hd__a21oi_1 _16120_ (.A1(net573),
    .A2(_03089_),
    .B1(net1891),
    .Y(_01004_));
 sky130_fd_sc_hd__nand2_1 _16121_ (.A(\jtag.managementReadData[21] ),
    .B(net1612),
    .Y(_03090_));
 sky130_fd_sc_hd__a21oi_1 _16122_ (.A1(net573),
    .A2(_03090_),
    .B1(net1888),
    .Y(_01005_));
 sky130_fd_sc_hd__nand2_1 _16123_ (.A(\jtag.managementReadData[22] ),
    .B(net1612),
    .Y(_03091_));
 sky130_fd_sc_hd__a21oi_1 _16124_ (.A1(net573),
    .A2(_03091_),
    .B1(net1891),
    .Y(_01006_));
 sky130_fd_sc_hd__nand2_1 _16125_ (.A(\jtag.managementReadData[23] ),
    .B(net1612),
    .Y(_03092_));
 sky130_fd_sc_hd__a21oi_1 _16126_ (.A1(net573),
    .A2(_03092_),
    .B1(net1891),
    .Y(_01007_));
 sky130_fd_sc_hd__nand2_1 _16127_ (.A(\jtag.managementReadData[24] ),
    .B(net1612),
    .Y(_03093_));
 sky130_fd_sc_hd__a21oi_1 _16128_ (.A1(net573),
    .A2(_03093_),
    .B1(net1891),
    .Y(_01008_));
 sky130_fd_sc_hd__nand2_1 _16129_ (.A(\jtag.managementReadData[25] ),
    .B(net1612),
    .Y(_03094_));
 sky130_fd_sc_hd__a21oi_1 _16130_ (.A1(net573),
    .A2(_03094_),
    .B1(net1888),
    .Y(_01009_));
 sky130_fd_sc_hd__nand2_1 _16131_ (.A(\jtag.managementReadData[26] ),
    .B(net1611),
    .Y(_03095_));
 sky130_fd_sc_hd__a21oi_1 _16132_ (.A1(net574),
    .A2(_03095_),
    .B1(net1888),
    .Y(_01010_));
 sky130_fd_sc_hd__nand2_1 _16133_ (.A(\jtag.managementReadData[27] ),
    .B(net1611),
    .Y(_03096_));
 sky130_fd_sc_hd__a21oi_1 _16134_ (.A1(net574),
    .A2(_03096_),
    .B1(net1888),
    .Y(_01011_));
 sky130_fd_sc_hd__nand2_1 _16135_ (.A(\jtag.managementReadData[28] ),
    .B(net1611),
    .Y(_03097_));
 sky130_fd_sc_hd__a21oi_1 _16136_ (.A1(net574),
    .A2(_03097_),
    .B1(net1888),
    .Y(_01012_));
 sky130_fd_sc_hd__nand2_1 _16137_ (.A(\jtag.managementReadData[29] ),
    .B(net1613),
    .Y(_03098_));
 sky130_fd_sc_hd__a21oi_1 _16138_ (.A1(_03068_),
    .A2(_03098_),
    .B1(net1888),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _16139_ (.A(\jtag.managementReadData[30] ),
    .B(net1612),
    .Y(_03099_));
 sky130_fd_sc_hd__a21oi_1 _16140_ (.A1(net573),
    .A2(_03099_),
    .B1(net1888),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2_1 _16141_ (.A(\jtag.managementReadData[31] ),
    .B(net1611),
    .Y(_03100_));
 sky130_fd_sc_hd__a21oi_1 _16142_ (.A1(net574),
    .A2(_03100_),
    .B1(net1888),
    .Y(_01015_));
 sky130_fd_sc_hd__or4b_2 _16143_ (.A(\jtag.managementState[2] ),
    .B(_08704_),
    .C(_03816_),
    .D_N(\jtag.managementState[1] ),
    .X(_03101_));
 sky130_fd_sc_hd__nor2_1 _16144_ (.A(\jtag.dataBSRRegister.data[31] ),
    .B(\jtag.dataBSRRegister.data[30] ),
    .Y(_03102_));
 sky130_fd_sc_hd__or3_1 _16145_ (.A(\jtag.managementState[1] ),
    .B(_08705_),
    .C(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__or3b_1 _16146_ (.A(\jtag.managementState[2] ),
    .B(\jtag.managementState[0] ),
    .C_N(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__a21o_1 _16147_ (.A1(\jtag.managementState[1] ),
    .A2(net1191),
    .B1(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__o21a_1 _16148_ (.A1(net1175),
    .A2(_03102_),
    .B1(_03101_),
    .X(_03106_));
 sky130_fd_sc_hd__nor2_1 _16149_ (.A(net1887),
    .B(_03106_),
    .Y(_01016_));
 sky130_fd_sc_hd__a21o_1 _16150_ (.A1(_03816_),
    .A2(\jtag.dataBSRRegister.data[31] ),
    .B1(net1611),
    .X(_03107_));
 sky130_fd_sc_hd__a31o_1 _16151_ (.A1(_03101_),
    .A2(_03105_),
    .A3(_03107_),
    .B1(net1887),
    .X(_03108_));
 sky130_fd_sc_hd__o21ba_1 _16152_ (.A1(\jtag.managementState[1] ),
    .A2(_03104_),
    .B1_N(_03108_),
    .X(_01017_));
 sky130_fd_sc_hd__and4b_1 _16153_ (.A_N(\jtag.managementState[2] ),
    .B(\jtag.managementState[1] ),
    .C(\jtag.managementState[0] ),
    .D(net1856),
    .X(_03109_));
 sky130_fd_sc_hd__and3_1 _16154_ (.A(_03101_),
    .B(_03105_),
    .C(_03109_),
    .X(_01018_));
 sky130_fd_sc_hd__and2_1 _16155_ (.A(_00517_),
    .B(_02261_),
    .X(_03110_));
 sky130_fd_sc_hd__nor2_1 _16156_ (.A(net544),
    .B(_02261_),
    .Y(_03111_));
 sky130_fd_sc_hd__a41o_1 _16157_ (.A1(\core.csr.trapReturnVector[0] ),
    .A2(net1825),
    .A3(net1131),
    .A4(_03111_),
    .B1(_03110_),
    .X(_01019_));
 sky130_fd_sc_hd__o21a_1 _16158_ (.A1(\core.csr.trapReturnVector[1] ),
    .A2(net1128),
    .B1(net1830),
    .X(_03112_));
 sky130_fd_sc_hd__o211a_1 _16159_ (.A1(net1131),
    .A2(_02251_),
    .B1(_03111_),
    .C1(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__a21o_1 _16160_ (.A1(_00518_),
    .A2(_02261_),
    .B1(_03113_),
    .X(_01020_));
 sky130_fd_sc_hd__nand2_2 _16161_ (.A(_06851_),
    .B(_08759_),
    .Y(_03114_));
 sky130_fd_sc_hd__mux2_1 _16162_ (.A0(net1077),
    .A1(\core.registers[27][0] ),
    .S(net804),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _16163_ (.A0(net1080),
    .A1(\core.registers[27][1] ),
    .S(net804),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _16164_ (.A0(net1088),
    .A1(\core.registers[27][2] ),
    .S(net803),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _16165_ (.A0(net1089),
    .A1(\core.registers[27][3] ),
    .S(net804),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _16166_ (.A0(net1029),
    .A1(\core.registers[27][4] ),
    .S(net802),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _16167_ (.A0(net1032),
    .A1(\core.registers[27][5] ),
    .S(net803),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _16168_ (.A0(net1038),
    .A1(\core.registers[27][6] ),
    .S(net803),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _16169_ (.A0(net1138),
    .A1(\core.registers[27][7] ),
    .S(net802),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _16170_ (.A0(net897),
    .A1(\core.registers[27][8] ),
    .S(net803),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _16171_ (.A0(net900),
    .A1(\core.registers[27][9] ),
    .S(net802),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _16172_ (.A0(net757),
    .A1(\core.registers[27][10] ),
    .S(net802),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _16173_ (.A0(net764),
    .A1(\core.registers[27][11] ),
    .S(net802),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _16174_ (.A0(net731),
    .A1(\core.registers[27][12] ),
    .S(net802),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _16175_ (.A0(net735),
    .A1(\core.registers[27][13] ),
    .S(net803),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _16176_ (.A0(net737),
    .A1(\core.registers[27][14] ),
    .S(net801),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _16177_ (.A0(net741),
    .A1(\core.registers[27][15] ),
    .S(net803),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _16178_ (.A0(net831),
    .A1(\core.registers[27][16] ),
    .S(net803),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _16179_ (.A0(net834),
    .A1(\core.registers[27][17] ),
    .S(net801),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _16180_ (.A0(net841),
    .A1(\core.registers[27][18] ),
    .S(net802),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _16181_ (.A0(net842),
    .A1(\core.registers[27][19] ),
    .S(net801),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _16182_ (.A0(net846),
    .A1(\core.registers[27][20] ),
    .S(net801),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _16183_ (.A0(net851),
    .A1(\core.registers[27][21] ),
    .S(net801),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _16184_ (.A0(net855),
    .A1(\core.registers[27][22] ),
    .S(net803),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _16185_ (.A0(net861),
    .A1(\core.registers[27][23] ),
    .S(net801),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _16186_ (.A0(net993),
    .A1(\core.registers[27][24] ),
    .S(net801),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _16187_ (.A0(net997),
    .A1(\core.registers[27][25] ),
    .S(net801),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _16188_ (.A0(net1000),
    .A1(\core.registers[27][26] ),
    .S(net801),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _16189_ (.A0(net864),
    .A1(\core.registers[27][27] ),
    .S(net803),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _16190_ (.A0(net870),
    .A1(\core.registers[27][28] ),
    .S(net802),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _16191_ (.A0(net873),
    .A1(\core.registers[27][29] ),
    .S(net802),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _16192_ (.A0(net877),
    .A1(\core.registers[27][30] ),
    .S(net802),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _16193_ (.A0(net1026),
    .A1(\core.registers[27][31] ),
    .S(net801),
    .X(_01052_));
 sky130_fd_sc_hd__or2_4 _16194_ (.A(_08678_),
    .B(_08763_),
    .X(_03115_));
 sky130_fd_sc_hd__mux2_1 _16195_ (.A0(net1076),
    .A1(\core.registers[9][0] ),
    .S(net927),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _16196_ (.A0(net1080),
    .A1(\core.registers[9][1] ),
    .S(net925),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _16197_ (.A0(net1086),
    .A1(\core.registers[9][2] ),
    .S(net927),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _16198_ (.A0(net1089),
    .A1(\core.registers[9][3] ),
    .S(net924),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _16199_ (.A0(net1029),
    .A1(\core.registers[9][4] ),
    .S(net925),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _16200_ (.A0(net1031),
    .A1(\core.registers[9][5] ),
    .S(net926),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _16201_ (.A0(net1038),
    .A1(\core.registers[9][6] ),
    .S(net926),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _16202_ (.A0(net1137),
    .A1(\core.registers[9][7] ),
    .S(net926),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _16203_ (.A0(net897),
    .A1(\core.registers[9][8] ),
    .S(net926),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _16204_ (.A0(net903),
    .A1(\core.registers[9][9] ),
    .S(net926),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _16205_ (.A0(net760),
    .A1(\core.registers[9][10] ),
    .S(net925),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _16206_ (.A0(net761),
    .A1(\core.registers[9][11] ),
    .S(net925),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _16207_ (.A0(net728),
    .A1(\core.registers[9][12] ),
    .S(net925),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _16208_ (.A0(net732),
    .A1(\core.registers[9][13] ),
    .S(net925),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _16209_ (.A0(net736),
    .A1(\core.registers[9][14] ),
    .S(net924),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _16210_ (.A0(net740),
    .A1(\core.registers[9][15] ),
    .S(net927),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _16211_ (.A0(net831),
    .A1(\core.registers[9][16] ),
    .S(net926),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _16212_ (.A0(net834),
    .A1(\core.registers[9][17] ),
    .S(net927),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _16213_ (.A0(net840),
    .A1(\core.registers[9][18] ),
    .S(net925),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _16214_ (.A0(net843),
    .A1(\core.registers[9][19] ),
    .S(net924),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _16215_ (.A0(net846),
    .A1(\core.registers[9][20] ),
    .S(net924),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _16216_ (.A0(net850),
    .A1(\core.registers[9][21] ),
    .S(net924),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _16217_ (.A0(net856),
    .A1(\core.registers[9][22] ),
    .S(net926),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _16218_ (.A0(net860),
    .A1(\core.registers[9][23] ),
    .S(net924),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _16219_ (.A0(net992),
    .A1(\core.registers[9][24] ),
    .S(net924),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _16220_ (.A0(net996),
    .A1(\core.registers[9][25] ),
    .S(net924),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _16221_ (.A0(net1000),
    .A1(\core.registers[9][26] ),
    .S(net924),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _16222_ (.A0(net864),
    .A1(\core.registers[9][27] ),
    .S(net926),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _16223_ (.A0(net870),
    .A1(\core.registers[9][28] ),
    .S(net925),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _16224_ (.A0(net876),
    .A1(\core.registers[9][29] ),
    .S(net925),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _16225_ (.A0(net877),
    .A1(\core.registers[9][30] ),
    .S(net925),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _16226_ (.A0(net1026),
    .A1(\core.registers[9][31] ),
    .S(net924),
    .X(_01084_));
 sky130_fd_sc_hd__nand2_1 _16227_ (.A(_08680_),
    .B(_08759_),
    .Y(_03116_));
 sky130_fd_sc_hd__mux2_1 _16228_ (.A0(net1077),
    .A1(\core.registers[24][0] ),
    .S(net920),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _16229_ (.A0(net1080),
    .A1(\core.registers[24][1] ),
    .S(net922),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _16230_ (.A0(net1088),
    .A1(\core.registers[24][2] ),
    .S(net922),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _16231_ (.A0(net1091),
    .A1(\core.registers[24][3] ),
    .S(net923),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _16232_ (.A0(net1029),
    .A1(\core.registers[24][4] ),
    .S(net921),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _16233_ (.A0(net1032),
    .A1(\core.registers[24][5] ),
    .S(net922),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _16234_ (.A0(net1038),
    .A1(\core.registers[24][6] ),
    .S(net922),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _16235_ (.A0(net1137),
    .A1(\core.registers[24][7] ),
    .S(net921),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _16236_ (.A0(net896),
    .A1(\core.registers[24][8] ),
    .S(net921),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _16237_ (.A0(net901),
    .A1(\core.registers[24][9] ),
    .S(net922),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _16238_ (.A0(net757),
    .A1(\core.registers[24][10] ),
    .S(net921),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _16239_ (.A0(net764),
    .A1(\core.registers[24][11] ),
    .S(net921),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _16240_ (.A0(net731),
    .A1(\core.registers[24][12] ),
    .S(net922),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _16241_ (.A0(net735),
    .A1(\core.registers[24][13] ),
    .S(net921),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _16242_ (.A0(net736),
    .A1(\core.registers[24][14] ),
    .S(net920),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _16243_ (.A0(net741),
    .A1(\core.registers[24][15] ),
    .S(net923),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _16244_ (.A0(net831),
    .A1(\core.registers[24][16] ),
    .S(net922),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _16245_ (.A0(net835),
    .A1(\core.registers[24][17] ),
    .S(net923),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _16246_ (.A0(net841),
    .A1(\core.registers[24][18] ),
    .S(net921),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _16247_ (.A0(net842),
    .A1(\core.registers[24][19] ),
    .S(net920),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _16248_ (.A0(net846),
    .A1(\core.registers[24][20] ),
    .S(net920),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _16249_ (.A0(net851),
    .A1(\core.registers[24][21] ),
    .S(net920),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _16250_ (.A0(net855),
    .A1(\core.registers[24][22] ),
    .S(net922),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _16251_ (.A0(net860),
    .A1(\core.registers[24][23] ),
    .S(net920),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _16252_ (.A0(net993),
    .A1(\core.registers[24][24] ),
    .S(net920),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _16253_ (.A0(net996),
    .A1(\core.registers[24][25] ),
    .S(net920),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _16254_ (.A0(net1000),
    .A1(\core.registers[24][26] ),
    .S(net920),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _16255_ (.A0(net865),
    .A1(\core.registers[24][27] ),
    .S(net922),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _16256_ (.A0(net870),
    .A1(\core.registers[24][28] ),
    .S(net921),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _16257_ (.A0(net873),
    .A1(\core.registers[24][29] ),
    .S(net921),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _16258_ (.A0(net877),
    .A1(\core.registers[24][30] ),
    .S(net921),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _16259_ (.A0(net1026),
    .A1(\core.registers[24][31] ),
    .S(net920),
    .X(_01116_));
 sky130_fd_sc_hd__nand2_1 _16260_ (.A(_08677_),
    .B(_08759_),
    .Y(_03117_));
 sky130_fd_sc_hd__mux2_1 _16261_ (.A0(net1076),
    .A1(\core.registers[25][0] ),
    .S(net916),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _16262_ (.A0(net1080),
    .A1(\core.registers[25][1] ),
    .S(net918),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _16263_ (.A0(net1088),
    .A1(\core.registers[25][2] ),
    .S(net918),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _16264_ (.A0(net1091),
    .A1(\core.registers[25][3] ),
    .S(net919),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _16265_ (.A0(net1029),
    .A1(\core.registers[25][4] ),
    .S(net917),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _16266_ (.A0(net1032),
    .A1(\core.registers[25][5] ),
    .S(net918),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _16267_ (.A0(net1038),
    .A1(\core.registers[25][6] ),
    .S(net917),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _16268_ (.A0(net1138),
    .A1(\core.registers[25][7] ),
    .S(net917),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _16269_ (.A0(net896),
    .A1(\core.registers[25][8] ),
    .S(net917),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _16270_ (.A0(net901),
    .A1(\core.registers[25][9] ),
    .S(net918),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _16271_ (.A0(net757),
    .A1(\core.registers[25][10] ),
    .S(net917),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _16272_ (.A0(net764),
    .A1(\core.registers[25][11] ),
    .S(net917),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _16273_ (.A0(net731),
    .A1(\core.registers[25][12] ),
    .S(net918),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _16274_ (.A0(net735),
    .A1(\core.registers[25][13] ),
    .S(net917),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _16275_ (.A0(net736),
    .A1(\core.registers[25][14] ),
    .S(net916),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _16276_ (.A0(net743),
    .A1(\core.registers[25][15] ),
    .S(net919),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _16277_ (.A0(net831),
    .A1(\core.registers[25][16] ),
    .S(net918),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _16278_ (.A0(net835),
    .A1(\core.registers[25][17] ),
    .S(net919),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _16279_ (.A0(net841),
    .A1(\core.registers[25][18] ),
    .S(net918),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _16280_ (.A0(net842),
    .A1(\core.registers[25][19] ),
    .S(net916),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _16281_ (.A0(net846),
    .A1(\core.registers[25][20] ),
    .S(net916),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _16282_ (.A0(net851),
    .A1(\core.registers[25][21] ),
    .S(net916),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _16283_ (.A0(net855),
    .A1(\core.registers[25][22] ),
    .S(net918),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _16284_ (.A0(net860),
    .A1(\core.registers[25][23] ),
    .S(net916),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _16285_ (.A0(net993),
    .A1(\core.registers[25][24] ),
    .S(net916),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _16286_ (.A0(net996),
    .A1(\core.registers[25][25] ),
    .S(net916),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _16287_ (.A0(net1000),
    .A1(\core.registers[25][26] ),
    .S(net916),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _16288_ (.A0(net865),
    .A1(\core.registers[25][27] ),
    .S(net918),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _16289_ (.A0(net870),
    .A1(\core.registers[25][28] ),
    .S(net917),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _16290_ (.A0(net873),
    .A1(\core.registers[25][29] ),
    .S(net917),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _16291_ (.A0(net877),
    .A1(\core.registers[25][30] ),
    .S(net917),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _16292_ (.A0(net1026),
    .A1(\core.registers[25][31] ),
    .S(net916),
    .X(_01148_));
 sky130_fd_sc_hd__nand2_2 _16293_ (.A(_06851_),
    .B(_08770_),
    .Y(_03118_));
 sky130_fd_sc_hd__mux2_1 _16294_ (.A0(net1076),
    .A1(\core.registers[15][0] ),
    .S(net800),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _16295_ (.A0(net1080),
    .A1(\core.registers[15][1] ),
    .S(net798),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _16296_ (.A0(net1085),
    .A1(\core.registers[15][2] ),
    .S(net800),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _16297_ (.A0(net1089),
    .A1(\core.registers[15][3] ),
    .S(net797),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _16298_ (.A0(net1027),
    .A1(\core.registers[15][4] ),
    .S(net798),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _16299_ (.A0(net1031),
    .A1(\core.registers[15][5] ),
    .S(net798),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _16300_ (.A0(net1038),
    .A1(\core.registers[15][6] ),
    .S(net798),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _16301_ (.A0(net1137),
    .A1(\core.registers[15][7] ),
    .S(net798),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _16302_ (.A0(net896),
    .A1(\core.registers[15][8] ),
    .S(net799),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _16303_ (.A0(net900),
    .A1(\core.registers[15][9] ),
    .S(net799),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _16304_ (.A0(net758),
    .A1(\core.registers[15][10] ),
    .S(net798),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _16305_ (.A0(net762),
    .A1(\core.registers[15][11] ),
    .S(net799),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _16306_ (.A0(net728),
    .A1(\core.registers[15][12] ),
    .S(net799),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _16307_ (.A0(net732),
    .A1(\core.registers[15][13] ),
    .S(net799),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _16308_ (.A0(net737),
    .A1(\core.registers[15][14] ),
    .S(net797),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _16309_ (.A0(net740),
    .A1(\core.registers[15][15] ),
    .S(net797),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _16310_ (.A0(net830),
    .A1(\core.registers[15][16] ),
    .S(net798),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _16311_ (.A0(net834),
    .A1(\core.registers[15][17] ),
    .S(net800),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _16312_ (.A0(net840),
    .A1(\core.registers[15][18] ),
    .S(net799),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _16313_ (.A0(net844),
    .A1(\core.registers[15][19] ),
    .S(net797),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _16314_ (.A0(net847),
    .A1(\core.registers[15][20] ),
    .S(net797),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _16315_ (.A0(net850),
    .A1(\core.registers[15][21] ),
    .S(net797),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _16316_ (.A0(net855),
    .A1(\core.registers[15][22] ),
    .S(net798),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _16317_ (.A0(net860),
    .A1(\core.registers[15][23] ),
    .S(net797),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _16318_ (.A0(net992),
    .A1(\core.registers[15][24] ),
    .S(net797),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _16319_ (.A0(net996),
    .A1(\core.registers[15][25] ),
    .S(net797),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _16320_ (.A0(net1000),
    .A1(\core.registers[15][26] ),
    .S(net797),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _16321_ (.A0(net865),
    .A1(\core.registers[15][27] ),
    .S(net798),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _16322_ (.A0(net869),
    .A1(\core.registers[15][28] ),
    .S(net799),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _16323_ (.A0(net876),
    .A1(\core.registers[15][29] ),
    .S(net798),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _16324_ (.A0(net878),
    .A1(\core.registers[15][30] ),
    .S(net799),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _16325_ (.A0(net1025),
    .A1(\core.registers[15][31] ),
    .S(net800),
    .X(_01180_));
 sky130_fd_sc_hd__nor2_8 _16326_ (.A(_08760_),
    .B(_08766_),
    .Y(_03119_));
 sky130_fd_sc_hd__mux2_1 _16327_ (.A0(\core.registers[6][0] ),
    .A1(net1078),
    .S(net793),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _16328_ (.A0(\core.registers[6][1] ),
    .A1(net1081),
    .S(net796),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _16329_ (.A0(\core.registers[6][2] ),
    .A1(net1086),
    .S(net794),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _16330_ (.A0(\core.registers[6][3] ),
    .A1(net1092),
    .S(net793),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _16331_ (.A0(\core.registers[6][4] ),
    .A1(net1028),
    .S(net796),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _16332_ (.A0(\core.registers[6][5] ),
    .A1(net1033),
    .S(net794),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _16333_ (.A0(\core.registers[6][6] ),
    .A1(net1035),
    .S(net794),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _16334_ (.A0(\core.registers[6][7] ),
    .A1(net1140),
    .S(net796),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _16335_ (.A0(\core.registers[6][8] ),
    .A1(net898),
    .S(net795),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _16336_ (.A0(\core.registers[6][9] ),
    .A1(net902),
    .S(net795),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _16337_ (.A0(\core.registers[6][10] ),
    .A1(net759),
    .S(net795),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _16338_ (.A0(\core.registers[6][11] ),
    .A1(net762),
    .S(net795),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _16339_ (.A0(\core.registers[6][12] ),
    .A1(net729),
    .S(net795),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _16340_ (.A0(\core.registers[6][13] ),
    .A1(net733),
    .S(net795),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _16341_ (.A0(\core.registers[6][14] ),
    .A1(net738),
    .S(net793),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _16342_ (.A0(\core.registers[6][15] ),
    .A1(net742),
    .S(net794),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _16343_ (.A0(\core.registers[6][16] ),
    .A1(net832),
    .S(net794),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _16344_ (.A0(\core.registers[6][17] ),
    .A1(net837),
    .S(net793),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _16345_ (.A0(\core.registers[6][18] ),
    .A1(net839),
    .S(net796),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _16346_ (.A0(\core.registers[6][19] ),
    .A1(net845),
    .S(net793),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _16347_ (.A0(\core.registers[6][20] ),
    .A1(net848),
    .S(net793),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _16348_ (.A0(\core.registers[6][21] ),
    .A1(net852),
    .S(net793),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _16349_ (.A0(\core.registers[6][22] ),
    .A1(net857),
    .S(net794),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _16350_ (.A0(\core.registers[6][23] ),
    .A1(net862),
    .S(net793),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _16351_ (.A0(\core.registers[6][24] ),
    .A1(net995),
    .S(net793),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _16352_ (.A0(\core.registers[6][25] ),
    .A1(net998),
    .S(net794),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _16353_ (.A0(\core.registers[6][26] ),
    .A1(net1002),
    .S(net795),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _16354_ (.A0(\core.registers[6][27] ),
    .A1(net866),
    .S(net795),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _16355_ (.A0(\core.registers[6][28] ),
    .A1(net871),
    .S(net796),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _16356_ (.A0(\core.registers[6][29] ),
    .A1(net874),
    .S(net795),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _16357_ (.A0(\core.registers[6][30] ),
    .A1(net879),
    .S(net795),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _16358_ (.A0(\core.registers[6][31] ),
    .A1(net1024),
    .S(net793),
    .X(_01212_));
 sky130_fd_sc_hd__or2_4 _16359_ (.A(_08678_),
    .B(_08766_),
    .X(_03120_));
 sky130_fd_sc_hd__mux2_1 _16360_ (.A0(net1077),
    .A1(\core.registers[5][0] ),
    .S(net912),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _16361_ (.A0(net1081),
    .A1(\core.registers[5][1] ),
    .S(net915),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _16362_ (.A0(net1087),
    .A1(\core.registers[5][2] ),
    .S(net913),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _16363_ (.A0(net1092),
    .A1(\core.registers[5][3] ),
    .S(net912),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _16364_ (.A0(net1028),
    .A1(\core.registers[5][4] ),
    .S(net913),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _16365_ (.A0(net1034),
    .A1(\core.registers[5][5] ),
    .S(net913),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _16366_ (.A0(net1035),
    .A1(\core.registers[5][6] ),
    .S(net913),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _16367_ (.A0(net1139),
    .A1(\core.registers[5][7] ),
    .S(net915),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _16368_ (.A0(net898),
    .A1(\core.registers[5][8] ),
    .S(net914),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _16369_ (.A0(net902),
    .A1(\core.registers[5][9] ),
    .S(net914),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _16370_ (.A0(net760),
    .A1(\core.registers[5][10] ),
    .S(net914),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _16371_ (.A0(net763),
    .A1(\core.registers[5][11] ),
    .S(net914),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _16372_ (.A0(net728),
    .A1(\core.registers[5][12] ),
    .S(net914),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _16373_ (.A0(net732),
    .A1(\core.registers[5][13] ),
    .S(net914),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _16374_ (.A0(net739),
    .A1(\core.registers[5][14] ),
    .S(net912),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _16375_ (.A0(net742),
    .A1(\core.registers[5][15] ),
    .S(net913),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _16376_ (.A0(net833),
    .A1(\core.registers[5][16] ),
    .S(net913),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _16377_ (.A0(net837),
    .A1(\core.registers[5][17] ),
    .S(net912),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _16378_ (.A0(net838),
    .A1(\core.registers[5][18] ),
    .S(net914),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _16379_ (.A0(net844),
    .A1(\core.registers[5][19] ),
    .S(net912),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _16380_ (.A0(net848),
    .A1(\core.registers[5][20] ),
    .S(net912),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _16381_ (.A0(net853),
    .A1(\core.registers[5][21] ),
    .S(net912),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _16382_ (.A0(net857),
    .A1(\core.registers[5][22] ),
    .S(net913),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _16383_ (.A0(net863),
    .A1(\core.registers[5][23] ),
    .S(net912),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _16384_ (.A0(net995),
    .A1(\core.registers[5][24] ),
    .S(net912),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _16385_ (.A0(net999),
    .A1(\core.registers[5][25] ),
    .S(net913),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _16386_ (.A0(net1003),
    .A1(\core.registers[5][26] ),
    .S(net915),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _16387_ (.A0(net866),
    .A1(\core.registers[5][27] ),
    .S(net914),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _16388_ (.A0(net871),
    .A1(\core.registers[5][28] ),
    .S(net915),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _16389_ (.A0(net875),
    .A1(\core.registers[5][29] ),
    .S(net914),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _16390_ (.A0(net879),
    .A1(\core.registers[5][30] ),
    .S(net914),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _16391_ (.A0(net1023),
    .A1(\core.registers[5][31] ),
    .S(net912),
    .X(_01244_));
 sky130_fd_sc_hd__and3_2 _16392_ (.A(\core.csr.currentInstruction[10] ),
    .B(net1801),
    .C(_03904_),
    .X(_03121_));
 sky130_fd_sc_hd__nand2_2 _16393_ (.A(_08677_),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__mux2_1 _16394_ (.A0(net1076),
    .A1(\core.registers[29][0] ),
    .S(net911),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _16395_ (.A0(net1082),
    .A1(\core.registers[29][1] ),
    .S(net909),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _16396_ (.A0(net1088),
    .A1(\core.registers[29][2] ),
    .S(net911),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _16397_ (.A0(net1090),
    .A1(\core.registers[29][3] ),
    .S(net911),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _16398_ (.A0(net1029),
    .A1(\core.registers[29][4] ),
    .S(net910),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _16399_ (.A0(net1031),
    .A1(\core.registers[29][5] ),
    .S(net910),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _16400_ (.A0(net1037),
    .A1(\core.registers[29][6] ),
    .S(net910),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _16401_ (.A0(net1138),
    .A1(\core.registers[29][7] ),
    .S(net909),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _16402_ (.A0(net899),
    .A1(\core.registers[29][8] ),
    .S(net909),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _16403_ (.A0(net901),
    .A1(\core.registers[29][9] ),
    .S(net909),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _16404_ (.A0(net757),
    .A1(\core.registers[29][10] ),
    .S(net909),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _16405_ (.A0(net764),
    .A1(\core.registers[29][11] ),
    .S(net909),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _16406_ (.A0(net731),
    .A1(\core.registers[29][12] ),
    .S(net910),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _16407_ (.A0(net735),
    .A1(\core.registers[29][13] ),
    .S(net910),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _16408_ (.A0(net737),
    .A1(\core.registers[29][14] ),
    .S(net908),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _16409_ (.A0(net741),
    .A1(\core.registers[29][15] ),
    .S(net908),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _16410_ (.A0(net831),
    .A1(\core.registers[29][16] ),
    .S(net910),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _16411_ (.A0(net836),
    .A1(\core.registers[29][17] ),
    .S(net908),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _16412_ (.A0(net841),
    .A1(\core.registers[29][18] ),
    .S(net909),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _16413_ (.A0(net842),
    .A1(\core.registers[29][19] ),
    .S(net908),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _16414_ (.A0(net846),
    .A1(\core.registers[29][20] ),
    .S(net908),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _16415_ (.A0(net851),
    .A1(\core.registers[29][21] ),
    .S(net908),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _16416_ (.A0(net856),
    .A1(\core.registers[29][22] ),
    .S(net910),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _16417_ (.A0(net861),
    .A1(\core.registers[29][23] ),
    .S(net908),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _16418_ (.A0(net993),
    .A1(\core.registers[29][24] ),
    .S(net908),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _16419_ (.A0(net997),
    .A1(\core.registers[29][25] ),
    .S(net908),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _16420_ (.A0(net1001),
    .A1(\core.registers[29][26] ),
    .S(net908),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _16421_ (.A0(net864),
    .A1(\core.registers[29][27] ),
    .S(net910),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _16422_ (.A0(net870),
    .A1(\core.registers[29][28] ),
    .S(net909),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _16423_ (.A0(net873),
    .A1(\core.registers[29][29] ),
    .S(net909),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _16424_ (.A0(net879),
    .A1(\core.registers[29][30] ),
    .S(net909),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _16425_ (.A0(net1025),
    .A1(\core.registers[29][31] ),
    .S(net911),
    .X(_01276_));
 sky130_fd_sc_hd__and2_1 _16426_ (.A(_08680_),
    .B(_03121_),
    .X(_03123_));
 sky130_fd_sc_hd__mux2_1 _16427_ (.A0(\core.registers[28][0] ),
    .A1(net1076),
    .S(net907),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _16428_ (.A0(\core.registers[28][1] ),
    .A1(net1082),
    .S(net905),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _16429_ (.A0(\core.registers[28][2] ),
    .A1(_04813_),
    .S(net906),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _16430_ (.A0(\core.registers[28][3] ),
    .A1(net1089),
    .S(net904),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _16431_ (.A0(\core.registers[28][4] ),
    .A1(net1029),
    .S(net906),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _16432_ (.A0(\core.registers[28][5] ),
    .A1(net1032),
    .S(net906),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _16433_ (.A0(\core.registers[28][6] ),
    .A1(net1037),
    .S(net906),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _16434_ (.A0(\core.registers[28][7] ),
    .A1(net1138),
    .S(net905),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _16435_ (.A0(\core.registers[28][8] ),
    .A1(net899),
    .S(net905),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _16436_ (.A0(\core.registers[28][9] ),
    .A1(net901),
    .S(net905),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _16437_ (.A0(\core.registers[28][10] ),
    .A1(net757),
    .S(net905),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _16438_ (.A0(\core.registers[28][11] ),
    .A1(net764),
    .S(net905),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _16439_ (.A0(\core.registers[28][12] ),
    .A1(net731),
    .S(net906),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _16440_ (.A0(\core.registers[28][13] ),
    .A1(net735),
    .S(net906),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _16441_ (.A0(\core.registers[28][14] ),
    .A1(net737),
    .S(net904),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _16442_ (.A0(\core.registers[28][15] ),
    .A1(net741),
    .S(net907),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _16443_ (.A0(\core.registers[28][16] ),
    .A1(net832),
    .S(net906),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _16444_ (.A0(\core.registers[28][17] ),
    .A1(net836),
    .S(net904),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _16445_ (.A0(\core.registers[28][18] ),
    .A1(net841),
    .S(net905),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _16446_ (.A0(\core.registers[28][19] ),
    .A1(net842),
    .S(net904),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _16447_ (.A0(\core.registers[28][20] ),
    .A1(net846),
    .S(net904),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _16448_ (.A0(\core.registers[28][21] ),
    .A1(net851),
    .S(net904),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _16449_ (.A0(\core.registers[28][22] ),
    .A1(net856),
    .S(net906),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _16450_ (.A0(\core.registers[28][23] ),
    .A1(net861),
    .S(net904),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _16451_ (.A0(\core.registers[28][24] ),
    .A1(net992),
    .S(net904),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _16452_ (.A0(\core.registers[28][25] ),
    .A1(net997),
    .S(net904),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _16453_ (.A0(\core.registers[28][26] ),
    .A1(net1001),
    .S(net904),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _16454_ (.A0(\core.registers[28][27] ),
    .A1(net864),
    .S(net906),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _16455_ (.A0(\core.registers[28][28] ),
    .A1(net870),
    .S(net905),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _16456_ (.A0(\core.registers[28][29] ),
    .A1(net873),
    .S(net905),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _16457_ (.A0(\core.registers[28][30] ),
    .A1(net879),
    .S(net905),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _16458_ (.A0(\core.registers[28][31] ),
    .A1(net1025),
    .S(net907),
    .X(_01308_));
 sky130_fd_sc_hd__or4b_4 _16459_ (.A(_03909_),
    .B(_06849_),
    .C(_08766_),
    .D_N(_03911_),
    .X(_03124_));
 sky130_fd_sc_hd__mux2_1 _16460_ (.A0(net1076),
    .A1(\core.registers[4][0] ),
    .S(net1007),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _16461_ (.A0(net1081),
    .A1(\core.registers[4][1] ),
    .S(net1010),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _16462_ (.A0(net1087),
    .A1(\core.registers[4][2] ),
    .S(net1008),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _16463_ (.A0(net1092),
    .A1(\core.registers[4][3] ),
    .S(net1007),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _16464_ (.A0(net1028),
    .A1(\core.registers[4][4] ),
    .S(net1008),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _16465_ (.A0(net1034),
    .A1(\core.registers[4][5] ),
    .S(net1008),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _16466_ (.A0(net1035),
    .A1(\core.registers[4][6] ),
    .S(net1008),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _16467_ (.A0(net1139),
    .A1(\core.registers[4][7] ),
    .S(net1010),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _16468_ (.A0(net898),
    .A1(\core.registers[4][8] ),
    .S(net1009),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _16469_ (.A0(net902),
    .A1(\core.registers[4][9] ),
    .S(net1009),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _16470_ (.A0(net760),
    .A1(\core.registers[4][10] ),
    .S(net1009),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _16471_ (.A0(net763),
    .A1(\core.registers[4][11] ),
    .S(net1009),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _16472_ (.A0(net730),
    .A1(\core.registers[4][12] ),
    .S(net1009),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _16473_ (.A0(net732),
    .A1(\core.registers[4][13] ),
    .S(net1009),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _16474_ (.A0(net739),
    .A1(\core.registers[4][14] ),
    .S(net1007),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _16475_ (.A0(net742),
    .A1(\core.registers[4][15] ),
    .S(net1008),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _16476_ (.A0(net833),
    .A1(\core.registers[4][16] ),
    .S(net1008),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _16477_ (.A0(net837),
    .A1(\core.registers[4][17] ),
    .S(net1007),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _16478_ (.A0(net838),
    .A1(\core.registers[4][18] ),
    .S(net1009),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _16479_ (.A0(net844),
    .A1(\core.registers[4][19] ),
    .S(net1007),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _16480_ (.A0(net848),
    .A1(\core.registers[4][20] ),
    .S(net1007),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _16481_ (.A0(net853),
    .A1(\core.registers[4][21] ),
    .S(net1007),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _16482_ (.A0(net857),
    .A1(\core.registers[4][22] ),
    .S(net1008),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _16483_ (.A0(net863),
    .A1(\core.registers[4][23] ),
    .S(net1007),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _16484_ (.A0(net995),
    .A1(\core.registers[4][24] ),
    .S(net1007),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _16485_ (.A0(net999),
    .A1(\core.registers[4][25] ),
    .S(net1008),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _16486_ (.A0(net1003),
    .A1(\core.registers[4][26] ),
    .S(net1010),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _16487_ (.A0(net866),
    .A1(\core.registers[4][27] ),
    .S(net1009),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _16488_ (.A0(net871),
    .A1(\core.registers[4][28] ),
    .S(net1010),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _16489_ (.A0(net875),
    .A1(\core.registers[4][29] ),
    .S(net1009),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _16490_ (.A0(net879),
    .A1(\core.registers[4][30] ),
    .S(net1009),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _16491_ (.A0(net1024),
    .A1(\core.registers[4][31] ),
    .S(net1007),
    .X(_01340_));
 sky130_fd_sc_hd__nand2_8 _16492_ (.A(_03908_),
    .B(_08761_),
    .Y(_03125_));
 sky130_fd_sc_hd__mux2_1 _16493_ (.A0(net1078),
    .A1(\core.registers[2][0] ),
    .S(net790),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _16494_ (.A0(net1083),
    .A1(\core.registers[2][1] ),
    .S(net792),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _16495_ (.A0(net1088),
    .A1(\core.registers[2][2] ),
    .S(net790),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _16496_ (.A0(net1092),
    .A1(\core.registers[2][3] ),
    .S(net789),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _16497_ (.A0(net1030),
    .A1(\core.registers[2][4] ),
    .S(net792),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _16498_ (.A0(net1033),
    .A1(\core.registers[2][5] ),
    .S(net790),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _16499_ (.A0(net1035),
    .A1(\core.registers[2][6] ),
    .S(net790),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _16500_ (.A0(net1139),
    .A1(\core.registers[2][7] ),
    .S(net792),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _16501_ (.A0(net898),
    .A1(\core.registers[2][8] ),
    .S(net791),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _16502_ (.A0(net902),
    .A1(\core.registers[2][9] ),
    .S(net791),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _16503_ (.A0(net759),
    .A1(\core.registers[2][10] ),
    .S(net791),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _16504_ (.A0(net762),
    .A1(\core.registers[2][11] ),
    .S(net791),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _16505_ (.A0(net730),
    .A1(\core.registers[2][12] ),
    .S(net791),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _16506_ (.A0(net734),
    .A1(\core.registers[2][13] ),
    .S(net791),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _16507_ (.A0(net739),
    .A1(\core.registers[2][14] ),
    .S(net789),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _16508_ (.A0(net742),
    .A1(\core.registers[2][15] ),
    .S(net790),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _16509_ (.A0(net832),
    .A1(\core.registers[2][16] ),
    .S(net790),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _16510_ (.A0(net837),
    .A1(\core.registers[2][17] ),
    .S(net789),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _16511_ (.A0(net839),
    .A1(\core.registers[2][18] ),
    .S(net791),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _16512_ (.A0(net845),
    .A1(\core.registers[2][19] ),
    .S(net789),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _16513_ (.A0(net848),
    .A1(\core.registers[2][20] ),
    .S(net789),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _16514_ (.A0(net853),
    .A1(\core.registers[2][21] ),
    .S(net789),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _16515_ (.A0(net857),
    .A1(\core.registers[2][22] ),
    .S(net790),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _16516_ (.A0(net863),
    .A1(\core.registers[2][23] ),
    .S(net789),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _16517_ (.A0(net995),
    .A1(\core.registers[2][24] ),
    .S(net789),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _16518_ (.A0(net998),
    .A1(\core.registers[2][25] ),
    .S(net789),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _16519_ (.A0(net1002),
    .A1(\core.registers[2][26] ),
    .S(net792),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _16520_ (.A0(net866),
    .A1(\core.registers[2][27] ),
    .S(net791),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _16521_ (.A0(net872),
    .A1(\core.registers[2][28] ),
    .S(net792),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _16522_ (.A0(net875),
    .A1(\core.registers[2][29] ),
    .S(net791),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _16523_ (.A0(net877),
    .A1(\core.registers[2][30] ),
    .S(net791),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _16524_ (.A0(net1024),
    .A1(\core.registers[2][31] ),
    .S(net789),
    .X(_01372_));
 sky130_fd_sc_hd__nand2_8 _16525_ (.A(_03908_),
    .B(_06851_),
    .Y(_03126_));
 sky130_fd_sc_hd__mux2_1 _16526_ (.A0(net1078),
    .A1(\core.registers[3][0] ),
    .S(net786),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _16527_ (.A0(net1083),
    .A1(\core.registers[3][1] ),
    .S(net788),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _16528_ (.A0(net1088),
    .A1(\core.registers[3][2] ),
    .S(net786),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _16529_ (.A0(net1092),
    .A1(\core.registers[3][3] ),
    .S(net785),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _16530_ (.A0(net1030),
    .A1(\core.registers[3][4] ),
    .S(net788),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _16531_ (.A0(net1033),
    .A1(\core.registers[3][5] ),
    .S(net786),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _16532_ (.A0(net1035),
    .A1(\core.registers[3][6] ),
    .S(net786),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _16533_ (.A0(net1140),
    .A1(\core.registers[3][7] ),
    .S(net788),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _16534_ (.A0(net899),
    .A1(\core.registers[3][8] ),
    .S(net787),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _16535_ (.A0(net902),
    .A1(\core.registers[3][9] ),
    .S(net787),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _16536_ (.A0(net759),
    .A1(\core.registers[3][10] ),
    .S(net787),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _16537_ (.A0(net762),
    .A1(\core.registers[3][11] ),
    .S(net787),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _16538_ (.A0(net730),
    .A1(\core.registers[3][12] ),
    .S(net787),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _16539_ (.A0(net734),
    .A1(\core.registers[3][13] ),
    .S(net787),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _16540_ (.A0(net738),
    .A1(\core.registers[3][14] ),
    .S(net785),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _16541_ (.A0(net742),
    .A1(\core.registers[3][15] ),
    .S(net786),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _16542_ (.A0(net832),
    .A1(\core.registers[3][16] ),
    .S(net786),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _16543_ (.A0(net837),
    .A1(\core.registers[3][17] ),
    .S(net785),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _16544_ (.A0(net839),
    .A1(\core.registers[3][18] ),
    .S(net787),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _16545_ (.A0(net845),
    .A1(\core.registers[3][19] ),
    .S(net785),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _16546_ (.A0(net848),
    .A1(\core.registers[3][20] ),
    .S(net785),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _16547_ (.A0(net853),
    .A1(\core.registers[3][21] ),
    .S(net785),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _16548_ (.A0(net857),
    .A1(\core.registers[3][22] ),
    .S(net786),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _16549_ (.A0(net863),
    .A1(\core.registers[3][23] ),
    .S(net785),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _16550_ (.A0(net995),
    .A1(\core.registers[3][24] ),
    .S(net785),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _16551_ (.A0(net998),
    .A1(\core.registers[3][25] ),
    .S(net785),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _16552_ (.A0(net1002),
    .A1(\core.registers[3][26] ),
    .S(net788),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _16553_ (.A0(net866),
    .A1(\core.registers[3][27] ),
    .S(net787),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _16554_ (.A0(net872),
    .A1(\core.registers[3][28] ),
    .S(net788),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _16555_ (.A0(net874),
    .A1(\core.registers[3][29] ),
    .S(net787),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _16556_ (.A0(net877),
    .A1(\core.registers[3][30] ),
    .S(net787),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _16557_ (.A0(net1024),
    .A1(\core.registers[3][31] ),
    .S(net785),
    .X(_01404_));
 sky130_fd_sc_hd__nand2_2 _16558_ (.A(_06851_),
    .B(_03121_),
    .Y(_03127_));
 sky130_fd_sc_hd__mux2_1 _16559_ (.A0(net1077),
    .A1(\core.registers[31][0] ),
    .S(net784),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _16560_ (.A0(net1082),
    .A1(\core.registers[31][1] ),
    .S(net782),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _16561_ (.A0(net1088),
    .A1(\core.registers[31][2] ),
    .S(net783),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _16562_ (.A0(net1089),
    .A1(\core.registers[31][3] ),
    .S(net784),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _16563_ (.A0(net1027),
    .A1(\core.registers[31][4] ),
    .S(net783),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _16564_ (.A0(net1031),
    .A1(\core.registers[31][5] ),
    .S(net783),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _16565_ (.A0(net1037),
    .A1(\core.registers[31][6] ),
    .S(net783),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _16566_ (.A0(net1137),
    .A1(\core.registers[31][7] ),
    .S(net782),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _16567_ (.A0(net896),
    .A1(\core.registers[31][8] ),
    .S(net782),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _16568_ (.A0(net901),
    .A1(\core.registers[31][9] ),
    .S(net782),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _16569_ (.A0(net757),
    .A1(\core.registers[31][10] ),
    .S(net782),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _16570_ (.A0(net764),
    .A1(\core.registers[31][11] ),
    .S(net782),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _16571_ (.A0(net731),
    .A1(\core.registers[31][12] ),
    .S(net783),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _16572_ (.A0(net735),
    .A1(\core.registers[31][13] ),
    .S(net783),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _16573_ (.A0(net736),
    .A1(\core.registers[31][14] ),
    .S(net781),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _16574_ (.A0(net741),
    .A1(\core.registers[31][15] ),
    .S(net781),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _16575_ (.A0(net831),
    .A1(\core.registers[31][16] ),
    .S(net783),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _16576_ (.A0(net835),
    .A1(\core.registers[31][17] ),
    .S(net781),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _16577_ (.A0(net841),
    .A1(\core.registers[31][18] ),
    .S(net782),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _16578_ (.A0(net842),
    .A1(\core.registers[31][19] ),
    .S(net781),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _16579_ (.A0(net846),
    .A1(\core.registers[31][20] ),
    .S(net781),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _16580_ (.A0(net851),
    .A1(\core.registers[31][21] ),
    .S(net781),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _16581_ (.A0(net856),
    .A1(\core.registers[31][22] ),
    .S(net783),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _16582_ (.A0(net861),
    .A1(\core.registers[31][23] ),
    .S(net781),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _16583_ (.A0(net994),
    .A1(\core.registers[31][24] ),
    .S(net781),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _16584_ (.A0(net997),
    .A1(\core.registers[31][25] ),
    .S(net781),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _16585_ (.A0(net1001),
    .A1(\core.registers[31][26] ),
    .S(net781),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _16586_ (.A0(net864),
    .A1(\core.registers[31][27] ),
    .S(net783),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _16587_ (.A0(net869),
    .A1(\core.registers[31][28] ),
    .S(net782),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _16588_ (.A0(net873),
    .A1(\core.registers[31][29] ),
    .S(net782),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _16589_ (.A0(net877),
    .A1(\core.registers[31][30] ),
    .S(net782),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _16590_ (.A0(net1025),
    .A1(\core.registers[31][31] ),
    .S(net784),
    .X(_01436_));
 sky130_fd_sc_hd__nand2_2 _16591_ (.A(_08761_),
    .B(_03121_),
    .Y(_03128_));
 sky130_fd_sc_hd__mux2_1 _16592_ (.A0(net1077),
    .A1(\core.registers[30][0] ),
    .S(net780),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _16593_ (.A0(net1082),
    .A1(\core.registers[30][1] ),
    .S(net778),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _16594_ (.A0(net1088),
    .A1(\core.registers[30][2] ),
    .S(net779),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _16595_ (.A0(net1090),
    .A1(\core.registers[30][3] ),
    .S(net780),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _16596_ (.A0(net1027),
    .A1(\core.registers[30][4] ),
    .S(net779),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _16597_ (.A0(net1032),
    .A1(\core.registers[30][5] ),
    .S(net779),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _16598_ (.A0(net1037),
    .A1(\core.registers[30][6] ),
    .S(net779),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _16599_ (.A0(net1137),
    .A1(\core.registers[30][7] ),
    .S(net778),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _16600_ (.A0(net896),
    .A1(\core.registers[30][8] ),
    .S(net778),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _16601_ (.A0(net901),
    .A1(\core.registers[30][9] ),
    .S(net778),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _16602_ (.A0(net757),
    .A1(\core.registers[30][10] ),
    .S(net778),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _16603_ (.A0(net764),
    .A1(\core.registers[30][11] ),
    .S(net778),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _16604_ (.A0(net731),
    .A1(\core.registers[30][12] ),
    .S(net779),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _16605_ (.A0(net735),
    .A1(\core.registers[30][13] ),
    .S(net779),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _16606_ (.A0(net736),
    .A1(\core.registers[30][14] ),
    .S(net777),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _16607_ (.A0(net741),
    .A1(\core.registers[30][15] ),
    .S(net777),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _16608_ (.A0(net831),
    .A1(\core.registers[30][16] ),
    .S(net779),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _16609_ (.A0(net836),
    .A1(\core.registers[30][17] ),
    .S(net777),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _16610_ (.A0(net841),
    .A1(\core.registers[30][18] ),
    .S(net778),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _16611_ (.A0(net842),
    .A1(\core.registers[30][19] ),
    .S(net777),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _16612_ (.A0(net846),
    .A1(\core.registers[30][20] ),
    .S(net777),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _16613_ (.A0(net850),
    .A1(\core.registers[30][21] ),
    .S(net777),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _16614_ (.A0(net856),
    .A1(\core.registers[30][22] ),
    .S(net779),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _16615_ (.A0(net861),
    .A1(\core.registers[30][23] ),
    .S(net777),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _16616_ (.A0(net994),
    .A1(\core.registers[30][24] ),
    .S(net777),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _16617_ (.A0(net997),
    .A1(\core.registers[30][25] ),
    .S(net777),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _16618_ (.A0(net1001),
    .A1(\core.registers[30][26] ),
    .S(net777),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _16619_ (.A0(net864),
    .A1(\core.registers[30][27] ),
    .S(net779),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _16620_ (.A0(net869),
    .A1(\core.registers[30][28] ),
    .S(net778),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _16621_ (.A0(net873),
    .A1(\core.registers[30][29] ),
    .S(net778),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _16622_ (.A0(net877),
    .A1(\core.registers[30][30] ),
    .S(net778),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _16623_ (.A0(net1025),
    .A1(\core.registers[30][31] ),
    .S(net780),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _16624_ (.A0(\wbSRAMInterface.currentByteSelect[0] ),
    .A1(net247),
    .S(net1287),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _16625_ (.A0(\wbSRAMInterface.currentByteSelect[1] ),
    .A1(net248),
    .S(net1287),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _16626_ (.A0(\wbSRAMInterface.currentByteSelect[2] ),
    .A1(net249),
    .S(net1287),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _16627_ (.A0(\wbSRAMInterface.currentByteSelect[3] ),
    .A1(net250),
    .S(net1287),
    .X(_01472_));
 sky130_fd_sc_hd__a41o_1 _16628_ (.A1(\core.pipe2_stall ),
    .A2(net1797),
    .A3(\core.pipe0_fetch.currentPipeStall ),
    .A4(net602),
    .B1(_03828_),
    .X(_03129_));
 sky130_fd_sc_hd__a21oi_1 _16629_ (.A1(_07046_),
    .A2(_03129_),
    .B1(net1886),
    .Y(_01473_));
 sky130_fd_sc_hd__a21oi_1 _16630_ (.A1(_03807_),
    .A2(\core.csr.instretTimer.currentValue[0] ),
    .B1(net1898),
    .Y(_03130_));
 sky130_fd_sc_hd__o21a_1 _16631_ (.A1(_03807_),
    .A2(\core.csr.instretTimer.currentValue[0] ),
    .B1(_03130_),
    .X(_01474_));
 sky130_fd_sc_hd__a21oi_1 _16632_ (.A1(_03807_),
    .A2(\core.csr.instretTimer.currentValue[0] ),
    .B1(\core.csr.instretTimer.currentValue[1] ),
    .Y(_03131_));
 sky130_fd_sc_hd__and3_2 _16633_ (.A(_03807_),
    .B(\core.csr.instretTimer.currentValue[1] ),
    .C(\core.csr.instretTimer.currentValue[0] ),
    .X(_03132_));
 sky130_fd_sc_hd__nor3_1 _16634_ (.A(net1898),
    .B(_03131_),
    .C(_03132_),
    .Y(_01475_));
 sky130_fd_sc_hd__a21oi_1 _16635_ (.A1(\core.csr.instretTimer.currentValue[2] ),
    .A2(_03132_),
    .B1(net1898),
    .Y(_03133_));
 sky130_fd_sc_hd__o21a_1 _16636_ (.A1(\core.csr.instretTimer.currentValue[2] ),
    .A2(_03132_),
    .B1(_03133_),
    .X(_01476_));
 sky130_fd_sc_hd__a21oi_1 _16637_ (.A1(\core.csr.instretTimer.currentValue[2] ),
    .A2(_03132_),
    .B1(\core.csr.instretTimer.currentValue[3] ),
    .Y(_03134_));
 sky130_fd_sc_hd__and3_1 _16638_ (.A(\core.csr.instretTimer.currentValue[3] ),
    .B(\core.csr.instretTimer.currentValue[2] ),
    .C(_03132_),
    .X(_03135_));
 sky130_fd_sc_hd__nor3_1 _16639_ (.A(net1898),
    .B(_03134_),
    .C(_03135_),
    .Y(_01477_));
 sky130_fd_sc_hd__and2_1 _16640_ (.A(\core.csr.instretTimer.currentValue[4] ),
    .B(_03135_),
    .X(_03136_));
 sky130_fd_sc_hd__nor2_1 _16641_ (.A(net1898),
    .B(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__o21a_1 _16642_ (.A1(\core.csr.instretTimer.currentValue[4] ),
    .A2(_03135_),
    .B1(_03137_),
    .X(_01478_));
 sky130_fd_sc_hd__and3_1 _16643_ (.A(\core.csr.instretTimer.currentValue[5] ),
    .B(\core.csr.instretTimer.currentValue[4] ),
    .C(_03135_),
    .X(_03138_));
 sky130_fd_sc_hd__nor2_1 _16644_ (.A(net1901),
    .B(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__o21a_1 _16645_ (.A1(\core.csr.instretTimer.currentValue[5] ),
    .A2(_03136_),
    .B1(_03139_),
    .X(_01479_));
 sky130_fd_sc_hd__and2_1 _16646_ (.A(\core.csr.instretTimer.currentValue[6] ),
    .B(_03138_),
    .X(_03140_));
 sky130_fd_sc_hd__o21ai_1 _16647_ (.A1(\core.csr.instretTimer.currentValue[6] ),
    .A2(_03138_),
    .B1(net1868),
    .Y(_03141_));
 sky130_fd_sc_hd__nor2_1 _16648_ (.A(_03140_),
    .B(_03141_),
    .Y(_01480_));
 sky130_fd_sc_hd__and3_1 _16649_ (.A(\core.csr.instretTimer.currentValue[7] ),
    .B(\core.csr.instretTimer.currentValue[6] ),
    .C(_03138_),
    .X(_03142_));
 sky130_fd_sc_hd__o21ai_1 _16650_ (.A1(\core.csr.instretTimer.currentValue[7] ),
    .A2(_03140_),
    .B1(net1868),
    .Y(_03143_));
 sky130_fd_sc_hd__nor2_1 _16651_ (.A(_03142_),
    .B(_03143_),
    .Y(_01481_));
 sky130_fd_sc_hd__and4_1 _16652_ (.A(\core.csr.instretTimer.currentValue[8] ),
    .B(\core.csr.instretTimer.currentValue[7] ),
    .C(\core.csr.instretTimer.currentValue[4] ),
    .D(\core.csr.instretTimer.currentValue[3] ),
    .X(_03144_));
 sky130_fd_sc_hd__and4_1 _16653_ (.A(\core.csr.instretTimer.currentValue[6] ),
    .B(\core.csr.instretTimer.currentValue[5] ),
    .C(\core.csr.instretTimer.currentValue[2] ),
    .D(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__and2_1 _16654_ (.A(\core.csr.instretTimer.currentValue[8] ),
    .B(_03142_),
    .X(_03146_));
 sky130_fd_sc_hd__nor2_1 _16655_ (.A(net1899),
    .B(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__o21a_1 _16656_ (.A1(\core.csr.instretTimer.currentValue[8] ),
    .A2(_03142_),
    .B1(_03147_),
    .X(_01482_));
 sky130_fd_sc_hd__nor2_1 _16657_ (.A(\core.csr.instretTimer.currentValue[9] ),
    .B(_03146_),
    .Y(_03148_));
 sky130_fd_sc_hd__and3_1 _16658_ (.A(\core.csr.instretTimer.currentValue[9] ),
    .B(\core.csr.instretTimer.currentValue[8] ),
    .C(_03142_),
    .X(_03149_));
 sky130_fd_sc_hd__nor3_1 _16659_ (.A(net1899),
    .B(_03148_),
    .C(_03149_),
    .Y(_01483_));
 sky130_fd_sc_hd__nor2_1 _16660_ (.A(\core.csr.instretTimer.currentValue[10] ),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__and3_1 _16661_ (.A(\core.csr.instretTimer.currentValue[10] ),
    .B(\core.csr.instretTimer.currentValue[9] ),
    .C(_03146_),
    .X(_03151_));
 sky130_fd_sc_hd__nor3_1 _16662_ (.A(net1899),
    .B(_03150_),
    .C(_03151_),
    .Y(_01484_));
 sky130_fd_sc_hd__nor2_1 _16663_ (.A(\core.csr.instretTimer.currentValue[11] ),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__and3_1 _16664_ (.A(\core.csr.instretTimer.currentValue[11] ),
    .B(\core.csr.instretTimer.currentValue[10] ),
    .C(_03149_),
    .X(_03153_));
 sky130_fd_sc_hd__nor3_1 _16665_ (.A(net1899),
    .B(_03152_),
    .C(_03153_),
    .Y(_01485_));
 sky130_fd_sc_hd__and4_1 _16666_ (.A(\core.csr.instretTimer.currentValue[12] ),
    .B(\core.csr.instretTimer.currentValue[11] ),
    .C(\core.csr.instretTimer.currentValue[10] ),
    .D(\core.csr.instretTimer.currentValue[9] ),
    .X(_03154_));
 sky130_fd_sc_hd__and3_1 _16667_ (.A(\core.csr.instretTimer.currentValue[12] ),
    .B(\core.csr.instretTimer.currentValue[11] ),
    .C(_03151_),
    .X(_03155_));
 sky130_fd_sc_hd__nor2_1 _16668_ (.A(net1899),
    .B(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__o21a_1 _16669_ (.A1(\core.csr.instretTimer.currentValue[12] ),
    .A2(_03153_),
    .B1(_03156_),
    .X(_01486_));
 sky130_fd_sc_hd__and3_1 _16670_ (.A(\core.csr.instretTimer.currentValue[13] ),
    .B(\core.csr.instretTimer.currentValue[12] ),
    .C(_03153_),
    .X(_03157_));
 sky130_fd_sc_hd__nor2_1 _16671_ (.A(net1900),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__o21a_1 _16672_ (.A1(\core.csr.instretTimer.currentValue[13] ),
    .A2(_03155_),
    .B1(_03158_),
    .X(_01487_));
 sky130_fd_sc_hd__nor2_1 _16673_ (.A(\core.csr.instretTimer.currentValue[14] ),
    .B(_03157_),
    .Y(_03159_));
 sky130_fd_sc_hd__and3_1 _16674_ (.A(\core.csr.instretTimer.currentValue[14] ),
    .B(\core.csr.instretTimer.currentValue[13] ),
    .C(_03155_),
    .X(_03160_));
 sky130_fd_sc_hd__nor3_1 _16675_ (.A(net1900),
    .B(_03159_),
    .C(_03160_),
    .Y(_01488_));
 sky130_fd_sc_hd__and3_1 _16676_ (.A(\core.csr.instretTimer.currentValue[15] ),
    .B(\core.csr.instretTimer.currentValue[14] ),
    .C(\core.csr.instretTimer.currentValue[13] ),
    .X(_03161_));
 sky130_fd_sc_hd__and4_2 _16677_ (.A(_03132_),
    .B(_03145_),
    .C(_03154_),
    .D(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__nor2_1 _16678_ (.A(net1900),
    .B(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__and4_1 _16679_ (.A(_03807_),
    .B(\core.csr.instretTimer.currentValue[14] ),
    .C(\core.csr.instretTimer.currentValue[10] ),
    .D(\core.csr.instretTimer.currentValue[6] ),
    .X(_03164_));
 sky130_fd_sc_hd__and4_1 _16680_ (.A(\core.csr.instretTimer.currentValue[3] ),
    .B(\core.csr.instretTimer.currentValue[1] ),
    .C(\core.csr.instretTimer.currentValue[0] ),
    .D(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__and4_1 _16681_ (.A(\core.csr.instretTimer.currentValue[13] ),
    .B(\core.csr.instretTimer.currentValue[12] ),
    .C(\core.csr.instretTimer.currentValue[9] ),
    .D(\core.csr.instretTimer.currentValue[4] ),
    .X(_03166_));
 sky130_fd_sc_hd__and4_1 _16682_ (.A(\core.csr.instretTimer.currentValue[15] ),
    .B(\core.csr.instretTimer.currentValue[11] ),
    .C(\core.csr.instretTimer.currentValue[7] ),
    .D(\core.csr.instretTimer.currentValue[2] ),
    .X(_03167_));
 sky130_fd_sc_hd__and4_1 _16683_ (.A(\core.csr.instretTimer.currentValue[8] ),
    .B(\core.csr.instretTimer.currentValue[5] ),
    .C(_03166_),
    .D(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__o21a_1 _16684_ (.A1(\core.csr.instretTimer.currentValue[15] ),
    .A2(_03160_),
    .B1(_03163_),
    .X(_01489_));
 sky130_fd_sc_hd__and2_1 _16685_ (.A(\core.csr.instretTimer.currentValue[16] ),
    .B(_03162_),
    .X(_03169_));
 sky130_fd_sc_hd__nor2_1 _16686_ (.A(net1901),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__o21a_1 _16687_ (.A1(\core.csr.instretTimer.currentValue[16] ),
    .A2(_03162_),
    .B1(_03170_),
    .X(_01490_));
 sky130_fd_sc_hd__and3_1 _16688_ (.A(\core.csr.instretTimer.currentValue[17] ),
    .B(\core.csr.instretTimer.currentValue[16] ),
    .C(_03162_),
    .X(_03171_));
 sky130_fd_sc_hd__nor2_1 _16689_ (.A(net1901),
    .B(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__and4_1 _16690_ (.A(\core.csr.instretTimer.currentValue[17] ),
    .B(\core.csr.instretTimer.currentValue[16] ),
    .C(_03165_),
    .D(_03168_),
    .X(_03173_));
 sky130_fd_sc_hd__o21a_1 _16691_ (.A1(\core.csr.instretTimer.currentValue[17] ),
    .A2(_03169_),
    .B1(_03172_),
    .X(_01491_));
 sky130_fd_sc_hd__a21oi_1 _16692_ (.A1(\core.csr.instretTimer.currentValue[18] ),
    .A2(_03171_),
    .B1(net1892),
    .Y(_03174_));
 sky130_fd_sc_hd__o21a_1 _16693_ (.A1(\core.csr.instretTimer.currentValue[18] ),
    .A2(_03173_),
    .B1(_03174_),
    .X(_01492_));
 sky130_fd_sc_hd__a21oi_1 _16694_ (.A1(\core.csr.instretTimer.currentValue[18] ),
    .A2(_03173_),
    .B1(\core.csr.instretTimer.currentValue[19] ),
    .Y(_03175_));
 sky130_fd_sc_hd__and3_1 _16695_ (.A(\core.csr.instretTimer.currentValue[19] ),
    .B(\core.csr.instretTimer.currentValue[18] ),
    .C(_03171_),
    .X(_03176_));
 sky130_fd_sc_hd__nor3_1 _16696_ (.A(net1895),
    .B(_03175_),
    .C(_03176_),
    .Y(_01493_));
 sky130_fd_sc_hd__and2_1 _16697_ (.A(\core.csr.instretTimer.currentValue[20] ),
    .B(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__nor2_1 _16698_ (.A(net1895),
    .B(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__and4_1 _16699_ (.A(\core.csr.instretTimer.currentValue[20] ),
    .B(\core.csr.instretTimer.currentValue[19] ),
    .C(\core.csr.instretTimer.currentValue[18] ),
    .D(_03173_),
    .X(_03179_));
 sky130_fd_sc_hd__o21a_1 _16700_ (.A1(\core.csr.instretTimer.currentValue[20] ),
    .A2(_03176_),
    .B1(_03178_),
    .X(_01494_));
 sky130_fd_sc_hd__nand2_1 _16701_ (.A(\core.csr.instretTimer.currentValue[21] ),
    .B(_03177_),
    .Y(_03180_));
 sky130_fd_sc_hd__o211a_1 _16702_ (.A1(\core.csr.instretTimer.currentValue[21] ),
    .A2(_03179_),
    .B1(_03180_),
    .C1(net1865),
    .X(_01495_));
 sky130_fd_sc_hd__a21oi_1 _16703_ (.A1(\core.csr.instretTimer.currentValue[21] ),
    .A2(_03179_),
    .B1(\core.csr.instretTimer.currentValue[22] ),
    .Y(_03181_));
 sky130_fd_sc_hd__and3_1 _16704_ (.A(\core.csr.instretTimer.currentValue[22] ),
    .B(\core.csr.instretTimer.currentValue[21] ),
    .C(_03177_),
    .X(_03182_));
 sky130_fd_sc_hd__nor3_1 _16705_ (.A(net1895),
    .B(_03181_),
    .C(_03182_),
    .Y(_01496_));
 sky130_fd_sc_hd__and2_1 _16706_ (.A(\core.csr.instretTimer.currentValue[23] ),
    .B(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__nor2_1 _16707_ (.A(net1895),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__and4_2 _16708_ (.A(\core.csr.instretTimer.currentValue[23] ),
    .B(\core.csr.instretTimer.currentValue[22] ),
    .C(\core.csr.instretTimer.currentValue[21] ),
    .D(_03179_),
    .X(_03185_));
 sky130_fd_sc_hd__o21a_1 _16709_ (.A1(\core.csr.instretTimer.currentValue[23] ),
    .A2(_03182_),
    .B1(_03184_),
    .X(_01497_));
 sky130_fd_sc_hd__a21oi_1 _16710_ (.A1(\core.csr.instretTimer.currentValue[24] ),
    .A2(_03185_),
    .B1(net1894),
    .Y(_03186_));
 sky130_fd_sc_hd__o21a_1 _16711_ (.A1(\core.csr.instretTimer.currentValue[24] ),
    .A2(_03185_),
    .B1(_03186_),
    .X(_01498_));
 sky130_fd_sc_hd__a21oi_1 _16712_ (.A1(\core.csr.instretTimer.currentValue[24] ),
    .A2(_03185_),
    .B1(\core.csr.instretTimer.currentValue[25] ),
    .Y(_03187_));
 sky130_fd_sc_hd__and3_1 _16713_ (.A(\core.csr.instretTimer.currentValue[25] ),
    .B(\core.csr.instretTimer.currentValue[24] ),
    .C(_03183_),
    .X(_03188_));
 sky130_fd_sc_hd__nor3_1 _16714_ (.A(net1894),
    .B(_03187_),
    .C(_03188_),
    .Y(_01499_));
 sky130_fd_sc_hd__and2_1 _16715_ (.A(\core.csr.instretTimer.currentValue[26] ),
    .B(_03188_),
    .X(_03189_));
 sky130_fd_sc_hd__nor2_1 _16716_ (.A(net1894),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__and4_2 _16717_ (.A(\core.csr.instretTimer.currentValue[26] ),
    .B(\core.csr.instretTimer.currentValue[25] ),
    .C(\core.csr.instretTimer.currentValue[24] ),
    .D(_03185_),
    .X(_03191_));
 sky130_fd_sc_hd__o21a_1 _16718_ (.A1(\core.csr.instretTimer.currentValue[26] ),
    .A2(_03188_),
    .B1(_03190_),
    .X(_01500_));
 sky130_fd_sc_hd__o21ai_1 _16719_ (.A1(\core.csr.instretTimer.currentValue[27] ),
    .A2(_03191_),
    .B1(net1865),
    .Y(_03192_));
 sky130_fd_sc_hd__a21oi_1 _16720_ (.A1(\core.csr.instretTimer.currentValue[27] ),
    .A2(_03191_),
    .B1(_03192_),
    .Y(_01501_));
 sky130_fd_sc_hd__a21oi_1 _16721_ (.A1(\core.csr.instretTimer.currentValue[27] ),
    .A2(_03191_),
    .B1(\core.csr.instretTimer.currentValue[28] ),
    .Y(_03193_));
 sky130_fd_sc_hd__and3_1 _16722_ (.A(\core.csr.instretTimer.currentValue[28] ),
    .B(\core.csr.instretTimer.currentValue[27] ),
    .C(_03189_),
    .X(_03194_));
 sky130_fd_sc_hd__and3_1 _16723_ (.A(\core.csr.instretTimer.currentValue[28] ),
    .B(\core.csr.instretTimer.currentValue[27] ),
    .C(_03191_),
    .X(_03195_));
 sky130_fd_sc_hd__nor3_1 _16724_ (.A(net1895),
    .B(_03193_),
    .C(_03195_),
    .Y(_01502_));
 sky130_fd_sc_hd__a21oi_1 _16725_ (.A1(\core.csr.instretTimer.currentValue[29] ),
    .A2(_03194_),
    .B1(net1892),
    .Y(_03196_));
 sky130_fd_sc_hd__o21a_1 _16726_ (.A1(\core.csr.instretTimer.currentValue[29] ),
    .A2(_03194_),
    .B1(_03196_),
    .X(_01503_));
 sky130_fd_sc_hd__a21oi_1 _16727_ (.A1(\core.csr.instretTimer.currentValue[29] ),
    .A2(_03195_),
    .B1(\core.csr.instretTimer.currentValue[30] ),
    .Y(_03197_));
 sky130_fd_sc_hd__and3_1 _16728_ (.A(\core.csr.instretTimer.currentValue[30] ),
    .B(\core.csr.instretTimer.currentValue[29] ),
    .C(_03194_),
    .X(_03198_));
 sky130_fd_sc_hd__and3_1 _16729_ (.A(\core.csr.instretTimer.currentValue[30] ),
    .B(\core.csr.instretTimer.currentValue[29] ),
    .C(_03195_),
    .X(_03199_));
 sky130_fd_sc_hd__nor3_1 _16730_ (.A(net1897),
    .B(_03197_),
    .C(_03199_),
    .Y(_01504_));
 sky130_fd_sc_hd__a21o_1 _16731_ (.A1(\core.csr.instretTimer.currentValue[31] ),
    .A2(_03198_),
    .B1(net1897),
    .X(_03200_));
 sky130_fd_sc_hd__o21ba_1 _16732_ (.A1(\core.csr.instretTimer.currentValue[31] ),
    .A2(_03198_),
    .B1_N(_03200_),
    .X(_01505_));
 sky130_fd_sc_hd__a21oi_1 _16733_ (.A1(\core.csr.instretTimer.currentValue[31] ),
    .A2(_03199_),
    .B1(\core.csr.instretTimer.currentValue[32] ),
    .Y(_03201_));
 sky130_fd_sc_hd__and3_1 _16734_ (.A(\core.csr.instretTimer.currentValue[32] ),
    .B(\core.csr.instretTimer.currentValue[31] ),
    .C(_03198_),
    .X(_03202_));
 sky130_fd_sc_hd__nor3_1 _16735_ (.A(net1897),
    .B(_03201_),
    .C(_03202_),
    .Y(_01506_));
 sky130_fd_sc_hd__and4_1 _16736_ (.A(\core.csr.instretTimer.currentValue[33] ),
    .B(\core.csr.instretTimer.currentValue[32] ),
    .C(\core.csr.instretTimer.currentValue[31] ),
    .D(_03199_),
    .X(_03203_));
 sky130_fd_sc_hd__nor2_1 _16737_ (.A(net1897),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__o21a_1 _16738_ (.A1(\core.csr.instretTimer.currentValue[33] ),
    .A2(_03202_),
    .B1(_03204_),
    .X(_01507_));
 sky130_fd_sc_hd__and3_1 _16739_ (.A(\core.csr.instretTimer.currentValue[34] ),
    .B(\core.csr.instretTimer.currentValue[33] ),
    .C(_03202_),
    .X(_03205_));
 sky130_fd_sc_hd__nor2_1 _16740_ (.A(net1901),
    .B(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__o21a_1 _16741_ (.A1(\core.csr.instretTimer.currentValue[34] ),
    .A2(_03203_),
    .B1(_03206_),
    .X(_01508_));
 sky130_fd_sc_hd__nor2_1 _16742_ (.A(\core.csr.instretTimer.currentValue[35] ),
    .B(_03205_),
    .Y(_03207_));
 sky130_fd_sc_hd__and3_1 _16743_ (.A(\core.csr.instretTimer.currentValue[35] ),
    .B(\core.csr.instretTimer.currentValue[34] ),
    .C(_03203_),
    .X(_03208_));
 sky130_fd_sc_hd__nor3_1 _16744_ (.A(net1898),
    .B(_03207_),
    .C(_03208_),
    .Y(_01509_));
 sky130_fd_sc_hd__nor2_1 _16745_ (.A(\core.csr.instretTimer.currentValue[36] ),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__and2_2 _16746_ (.A(\core.csr.instretTimer.currentValue[36] ),
    .B(_03208_),
    .X(_03210_));
 sky130_fd_sc_hd__nor3_1 _16747_ (.A(net1898),
    .B(_03209_),
    .C(_03210_),
    .Y(_01510_));
 sky130_fd_sc_hd__o21ai_1 _16748_ (.A1(\core.csr.instretTimer.currentValue[37] ),
    .A2(_03210_),
    .B1(net1868),
    .Y(_03211_));
 sky130_fd_sc_hd__a21oi_1 _16749_ (.A1(\core.csr.instretTimer.currentValue[37] ),
    .A2(_03210_),
    .B1(_03211_),
    .Y(_01511_));
 sky130_fd_sc_hd__a21oi_1 _16750_ (.A1(\core.csr.instretTimer.currentValue[37] ),
    .A2(_03210_),
    .B1(\core.csr.instretTimer.currentValue[38] ),
    .Y(_03212_));
 sky130_fd_sc_hd__and3_1 _16751_ (.A(\core.csr.instretTimer.currentValue[38] ),
    .B(\core.csr.instretTimer.currentValue[37] ),
    .C(_03210_),
    .X(_03213_));
 sky130_fd_sc_hd__nor3_1 _16752_ (.A(net1898),
    .B(_03212_),
    .C(_03213_),
    .Y(_01512_));
 sky130_fd_sc_hd__nor2_1 _16753_ (.A(\core.csr.instretTimer.currentValue[39] ),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__and2_2 _16754_ (.A(\core.csr.instretTimer.currentValue[39] ),
    .B(_03213_),
    .X(_03215_));
 sky130_fd_sc_hd__nor3_1 _16755_ (.A(net1899),
    .B(_03214_),
    .C(_03215_),
    .Y(_01513_));
 sky130_fd_sc_hd__o21ai_1 _16756_ (.A1(\core.csr.instretTimer.currentValue[40] ),
    .A2(_03215_),
    .B1(net1867),
    .Y(_03216_));
 sky130_fd_sc_hd__a21oi_1 _16757_ (.A1(\core.csr.instretTimer.currentValue[40] ),
    .A2(_03215_),
    .B1(_03216_),
    .Y(_01514_));
 sky130_fd_sc_hd__a21oi_1 _16758_ (.A1(\core.csr.instretTimer.currentValue[40] ),
    .A2(_03215_),
    .B1(\core.csr.instretTimer.currentValue[41] ),
    .Y(_03217_));
 sky130_fd_sc_hd__and3_1 _16759_ (.A(\core.csr.instretTimer.currentValue[41] ),
    .B(\core.csr.instretTimer.currentValue[40] ),
    .C(_03215_),
    .X(_03218_));
 sky130_fd_sc_hd__nor3_1 _16760_ (.A(net1899),
    .B(_03217_),
    .C(_03218_),
    .Y(_01515_));
 sky130_fd_sc_hd__nor2_1 _16761_ (.A(\core.csr.instretTimer.currentValue[42] ),
    .B(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__and2_2 _16762_ (.A(\core.csr.instretTimer.currentValue[42] ),
    .B(_03218_),
    .X(_03220_));
 sky130_fd_sc_hd__nor3_1 _16763_ (.A(net1899),
    .B(_03219_),
    .C(_03220_),
    .Y(_01516_));
 sky130_fd_sc_hd__o21ai_1 _16764_ (.A1(\core.csr.instretTimer.currentValue[43] ),
    .A2(_03220_),
    .B1(net1867),
    .Y(_03221_));
 sky130_fd_sc_hd__a21oi_1 _16765_ (.A1(\core.csr.instretTimer.currentValue[43] ),
    .A2(_03220_),
    .B1(_03221_),
    .Y(_01517_));
 sky130_fd_sc_hd__a21oi_1 _16766_ (.A1(\core.csr.instretTimer.currentValue[43] ),
    .A2(_03220_),
    .B1(\core.csr.instretTimer.currentValue[44] ),
    .Y(_03222_));
 sky130_fd_sc_hd__and3_1 _16767_ (.A(\core.csr.instretTimer.currentValue[44] ),
    .B(\core.csr.instretTimer.currentValue[43] ),
    .C(_03220_),
    .X(_03223_));
 sky130_fd_sc_hd__nor3_1 _16768_ (.A(net1899),
    .B(_03222_),
    .C(_03223_),
    .Y(_01518_));
 sky130_fd_sc_hd__nor2_1 _16769_ (.A(\core.csr.instretTimer.currentValue[45] ),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__and2_2 _16770_ (.A(\core.csr.instretTimer.currentValue[45] ),
    .B(_03223_),
    .X(_03225_));
 sky130_fd_sc_hd__nor3_1 _16771_ (.A(net1900),
    .B(_03224_),
    .C(_03225_),
    .Y(_01519_));
 sky130_fd_sc_hd__o21ai_1 _16772_ (.A1(\core.csr.instretTimer.currentValue[46] ),
    .A2(_03225_),
    .B1(net1868),
    .Y(_03226_));
 sky130_fd_sc_hd__a21oi_1 _16773_ (.A1(\core.csr.instretTimer.currentValue[46] ),
    .A2(_03225_),
    .B1(_03226_),
    .Y(_01520_));
 sky130_fd_sc_hd__a21oi_1 _16774_ (.A1(\core.csr.instretTimer.currentValue[46] ),
    .A2(_03225_),
    .B1(\core.csr.instretTimer.currentValue[47] ),
    .Y(_03227_));
 sky130_fd_sc_hd__and3_1 _16775_ (.A(\core.csr.instretTimer.currentValue[47] ),
    .B(\core.csr.instretTimer.currentValue[46] ),
    .C(_03225_),
    .X(_03228_));
 sky130_fd_sc_hd__nor3_1 _16776_ (.A(net1900),
    .B(_03227_),
    .C(_03228_),
    .Y(_01521_));
 sky130_fd_sc_hd__nor2_1 _16777_ (.A(\core.csr.instretTimer.currentValue[48] ),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__and2_2 _16778_ (.A(\core.csr.instretTimer.currentValue[48] ),
    .B(_03228_),
    .X(_03230_));
 sky130_fd_sc_hd__nor3_1 _16779_ (.A(net1902),
    .B(_03229_),
    .C(_03230_),
    .Y(_01522_));
 sky130_fd_sc_hd__o21ai_1 _16780_ (.A1(\core.csr.instretTimer.currentValue[49] ),
    .A2(_03230_),
    .B1(net1868),
    .Y(_03231_));
 sky130_fd_sc_hd__a21oi_1 _16781_ (.A1(\core.csr.instretTimer.currentValue[49] ),
    .A2(_03230_),
    .B1(_03231_),
    .Y(_01523_));
 sky130_fd_sc_hd__a21oi_1 _16782_ (.A1(\core.csr.instretTimer.currentValue[49] ),
    .A2(_03230_),
    .B1(\core.csr.instretTimer.currentValue[50] ),
    .Y(_03232_));
 sky130_fd_sc_hd__and3_1 _16783_ (.A(\core.csr.instretTimer.currentValue[50] ),
    .B(\core.csr.instretTimer.currentValue[49] ),
    .C(_03230_),
    .X(_03233_));
 sky130_fd_sc_hd__nor3_1 _16784_ (.A(net1902),
    .B(_03232_),
    .C(_03233_),
    .Y(_01524_));
 sky130_fd_sc_hd__nor2_1 _16785_ (.A(\core.csr.instretTimer.currentValue[51] ),
    .B(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__and2_2 _16786_ (.A(\core.csr.instretTimer.currentValue[51] ),
    .B(_03233_),
    .X(_03235_));
 sky130_fd_sc_hd__nor3_1 _16787_ (.A(net1902),
    .B(_03234_),
    .C(_03235_),
    .Y(_01525_));
 sky130_fd_sc_hd__o21ai_1 _16788_ (.A1(\core.csr.instretTimer.currentValue[52] ),
    .A2(_03235_),
    .B1(net1865),
    .Y(_03236_));
 sky130_fd_sc_hd__a21oi_1 _16789_ (.A1(\core.csr.instretTimer.currentValue[52] ),
    .A2(_03235_),
    .B1(_03236_),
    .Y(_01526_));
 sky130_fd_sc_hd__a21oi_1 _16790_ (.A1(\core.csr.instretTimer.currentValue[52] ),
    .A2(_03235_),
    .B1(\core.csr.instretTimer.currentValue[53] ),
    .Y(_03237_));
 sky130_fd_sc_hd__and3_1 _16791_ (.A(\core.csr.instretTimer.currentValue[53] ),
    .B(\core.csr.instretTimer.currentValue[52] ),
    .C(_03235_),
    .X(_03238_));
 sky130_fd_sc_hd__nor3_1 _16792_ (.A(net1895),
    .B(_03237_),
    .C(_03238_),
    .Y(_01527_));
 sky130_fd_sc_hd__nor2_1 _16793_ (.A(\core.csr.instretTimer.currentValue[54] ),
    .B(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__and2_2 _16794_ (.A(\core.csr.instretTimer.currentValue[54] ),
    .B(_03238_),
    .X(_03240_));
 sky130_fd_sc_hd__nor3_1 _16795_ (.A(net1895),
    .B(_03239_),
    .C(_03240_),
    .Y(_01528_));
 sky130_fd_sc_hd__o21ai_1 _16796_ (.A1(\core.csr.instretTimer.currentValue[55] ),
    .A2(_03240_),
    .B1(net1869),
    .Y(_03241_));
 sky130_fd_sc_hd__a21oi_1 _16797_ (.A1(\core.csr.instretTimer.currentValue[55] ),
    .A2(_03240_),
    .B1(_03241_),
    .Y(_01529_));
 sky130_fd_sc_hd__a21oi_1 _16798_ (.A1(\core.csr.instretTimer.currentValue[55] ),
    .A2(_03240_),
    .B1(\core.csr.instretTimer.currentValue[56] ),
    .Y(_03242_));
 sky130_fd_sc_hd__and3_1 _16799_ (.A(\core.csr.instretTimer.currentValue[56] ),
    .B(\core.csr.instretTimer.currentValue[55] ),
    .C(_03240_),
    .X(_03243_));
 sky130_fd_sc_hd__nor3_1 _16800_ (.A(net1896),
    .B(_03242_),
    .C(_03243_),
    .Y(_01530_));
 sky130_fd_sc_hd__nor2_1 _16801_ (.A(\core.csr.instretTimer.currentValue[57] ),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__and2_2 _16802_ (.A(\core.csr.instretTimer.currentValue[57] ),
    .B(_03243_),
    .X(_03245_));
 sky130_fd_sc_hd__nor3_1 _16803_ (.A(net1896),
    .B(_03244_),
    .C(_03245_),
    .Y(_01531_));
 sky130_fd_sc_hd__o21ai_1 _16804_ (.A1(\core.csr.instretTimer.currentValue[58] ),
    .A2(_03245_),
    .B1(net1869),
    .Y(_03246_));
 sky130_fd_sc_hd__a21oi_1 _16805_ (.A1(\core.csr.instretTimer.currentValue[58] ),
    .A2(_03245_),
    .B1(_03246_),
    .Y(_01532_));
 sky130_fd_sc_hd__a21oi_1 _16806_ (.A1(\core.csr.instretTimer.currentValue[58] ),
    .A2(_03245_),
    .B1(\core.csr.instretTimer.currentValue[59] ),
    .Y(_03247_));
 sky130_fd_sc_hd__and3_2 _16807_ (.A(\core.csr.instretTimer.currentValue[59] ),
    .B(\core.csr.instretTimer.currentValue[58] ),
    .C(_03245_),
    .X(_03248_));
 sky130_fd_sc_hd__nor3_1 _16808_ (.A(net1894),
    .B(_03247_),
    .C(_03248_),
    .Y(_01533_));
 sky130_fd_sc_hd__nor2_1 _16809_ (.A(\core.csr.instretTimer.currentValue[60] ),
    .B(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hd__and2_2 _16810_ (.A(\core.csr.instretTimer.currentValue[60] ),
    .B(_03248_),
    .X(_03250_));
 sky130_fd_sc_hd__nor3_1 _16811_ (.A(net1893),
    .B(_03249_),
    .C(_03250_),
    .Y(_01534_));
 sky130_fd_sc_hd__o21ai_1 _16812_ (.A1(\core.csr.instretTimer.currentValue[61] ),
    .A2(_03250_),
    .B1(net1869),
    .Y(_03251_));
 sky130_fd_sc_hd__a21oi_1 _16813_ (.A1(\core.csr.instretTimer.currentValue[61] ),
    .A2(_03250_),
    .B1(_03251_),
    .Y(_01535_));
 sky130_fd_sc_hd__a31o_1 _16814_ (.A1(\core.csr.instretTimer.currentValue[61] ),
    .A2(\core.csr.instretTimer.currentValue[60] ),
    .A3(_03248_),
    .B1(\core.csr.instretTimer.currentValue[62] ),
    .X(_03252_));
 sky130_fd_sc_hd__nand3_2 _16815_ (.A(\core.csr.instretTimer.currentValue[62] ),
    .B(\core.csr.instretTimer.currentValue[61] ),
    .C(_03250_),
    .Y(_03253_));
 sky130_fd_sc_hd__and3_1 _16816_ (.A(net1865),
    .B(_03252_),
    .C(_03253_),
    .X(_01536_));
 sky130_fd_sc_hd__o21ai_1 _16817_ (.A1(_03813_),
    .A2(_03253_),
    .B1(net1865),
    .Y(_03254_));
 sky130_fd_sc_hd__a21oi_1 _16818_ (.A1(_03813_),
    .A2(_03253_),
    .B1(_03254_),
    .Y(_01537_));
 sky130_fd_sc_hd__nor3_1 _16819_ (.A(_07037_),
    .B(_07041_),
    .C(_07159_),
    .Y(_03255_));
 sky130_fd_sc_hd__a31o_1 _16820_ (.A1(net1726),
    .A2(net1719),
    .A3(net1248),
    .B1(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__nand2_1 _16821_ (.A(net1726),
    .B(\core.csr.currentInstruction[23] ),
    .Y(_03257_));
 sky130_fd_sc_hd__and3_1 _16822_ (.A(_07166_),
    .B(_03256_),
    .C(_03257_),
    .X(_03258_));
 sky130_fd_sc_hd__mux2_2 _16823_ (.A0(\core.csr.currentInstruction[22] ),
    .A1(_07029_),
    .S(net1713),
    .X(_03259_));
 sky130_fd_sc_hd__nand2_1 _16824_ (.A(_03258_),
    .B(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__o21ba_4 _16825_ (.A1(net1713),
    .A2(\core.csr.currentInstruction[26] ),
    .B1_N(_07180_),
    .X(_03261_));
 sky130_fd_sc_hd__mux2_2 _16826_ (.A0(\core.csr.currentInstruction[20] ),
    .A1(_07033_),
    .S(net1713),
    .X(_03262_));
 sky130_fd_sc_hd__mux2_2 _16827_ (.A0(\core.csr.currentInstruction[21] ),
    .A1(_07032_),
    .S(net1713),
    .X(_03263_));
 sky130_fd_sc_hd__nand2b_1 _16828_ (.A_N(_03263_),
    .B(_03262_),
    .Y(_03264_));
 sky130_fd_sc_hd__a21o_1 _16829_ (.A1(net1726),
    .A2(\core.csr.currentInstruction[29] ),
    .B1(_07178_),
    .X(_03265_));
 sky130_fd_sc_hd__a21o_1 _16830_ (.A1(net1726),
    .A2(\core.csr.currentInstruction[28] ),
    .B1(_07176_),
    .X(_03266_));
 sky130_fd_sc_hd__nand2_1 _16831_ (.A(_03265_),
    .B(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__a21o_1 _16832_ (.A1(net1726),
    .A2(\core.csr.currentInstruction[25] ),
    .B1(_07188_),
    .X(_03268_));
 sky130_fd_sc_hd__a21o_1 _16833_ (.A1(net1726),
    .A2(\core.csr.currentInstruction[27] ),
    .B1(_07194_),
    .X(_03269_));
 sky130_fd_sc_hd__or2_1 _16834_ (.A(_03268_),
    .B(_03269_),
    .X(_03270_));
 sky130_fd_sc_hd__mux2_1 _16835_ (.A0(\core.csr.currentInstruction[24] ),
    .A1(_07024_),
    .S(net1713),
    .X(_03271_));
 sky130_fd_sc_hd__mux2_1 _16836_ (.A0(\core.csr.currentInstruction[31] ),
    .A1(_07016_),
    .S(net1713),
    .X(_03272_));
 sky130_fd_sc_hd__a21o_1 _16837_ (.A1(net1726),
    .A2(\core.csr.currentInstruction[30] ),
    .B1(_07185_),
    .X(_03273_));
 sky130_fd_sc_hd__and4bb_1 _16838_ (.A_N(_03261_),
    .B_N(_03270_),
    .C(_03271_),
    .D(_03273_),
    .X(_03274_));
 sky130_fd_sc_hd__nand2_1 _16839_ (.A(_07166_),
    .B(_03256_),
    .Y(_03275_));
 sky130_fd_sc_hd__nand3b_1 _16840_ (.A_N(_03275_),
    .B(_03257_),
    .C(_03259_),
    .Y(_03276_));
 sky130_fd_sc_hd__or2_4 _16841_ (.A(_03260_),
    .B(_03264_),
    .X(_03277_));
 sky130_fd_sc_hd__inv_2 _16842_ (.A(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__and4b_4 _16843_ (.A_N(_03267_),
    .B(_03272_),
    .C(_03274_),
    .D(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__mux2_2 _16844_ (.A0(_03830_),
    .A1(_02914_),
    .S(net1715),
    .X(_03280_));
 sky130_fd_sc_hd__inv_2 _16845_ (.A(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__nand2_1 _16846_ (.A(net626),
    .B(_03280_),
    .Y(_03282_));
 sky130_fd_sc_hd__o211a_1 _16847_ (.A1(\core.csr.mconfigptr.currentValue[0] ),
    .A2(net626),
    .B1(_03282_),
    .C1(net1850),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_4 _16848_ (.A0(_03829_),
    .A1(_02912_),
    .S(net1715),
    .X(_03283_));
 sky130_fd_sc_hd__clkinv_4 _16849_ (.A(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__nand2_1 _16850_ (.A(net626),
    .B(_03283_),
    .Y(_03285_));
 sky130_fd_sc_hd__o211a_1 _16851_ (.A1(\core.csr.mconfigptr.currentValue[1] ),
    .A2(net626),
    .B1(_03285_),
    .C1(net1850),
    .X(_01539_));
 sky130_fd_sc_hd__nand2_1 _16852_ (.A(net1725),
    .B(\core.pipe1_resultRegister[2] ),
    .Y(_03286_));
 sky130_fd_sc_hd__o21ai_4 _16853_ (.A1(net1725),
    .A2(_02910_),
    .B1(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__mux2_1 _16854_ (.A0(\core.csr.mconfigptr.currentValue[2] ),
    .A1(_03287_),
    .S(net626),
    .X(_03288_));
 sky130_fd_sc_hd__and2_1 _16855_ (.A(net1851),
    .B(_03288_),
    .X(_01540_));
 sky130_fd_sc_hd__a221o_2 _16856_ (.A1(\jtag.managementReadData[3] ),
    .A2(net1305),
    .B1(net1197),
    .B2(net240),
    .C1(net1724),
    .X(_03289_));
 sky130_fd_sc_hd__o21ai_4 _16857_ (.A1(net1713),
    .A2(\core.pipe1_resultRegister[3] ),
    .B1(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__nand2_1 _16858_ (.A(net626),
    .B(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__o211a_1 _16859_ (.A1(\core.csr.mconfigptr.currentValue[3] ),
    .A2(net626),
    .B1(_03291_),
    .C1(net1850),
    .X(_01541_));
 sky130_fd_sc_hd__a221o_1 _16860_ (.A1(\jtag.managementReadData[4] ),
    .A2(net1305),
    .B1(net1197),
    .B2(net241),
    .C1(net1724),
    .X(_03292_));
 sky130_fd_sc_hd__o21a_4 _16861_ (.A1(net1716),
    .A2(\core.pipe1_resultRegister[4] ),
    .B1(_03292_),
    .X(_03293_));
 sky130_fd_sc_hd__mux2_1 _16862_ (.A0(\core.csr.mconfigptr.currentValue[4] ),
    .A1(_03293_),
    .S(net629),
    .X(_03294_));
 sky130_fd_sc_hd__and2_1 _16863_ (.A(net1852),
    .B(_03294_),
    .X(_01542_));
 sky130_fd_sc_hd__a221o_1 _16864_ (.A1(\jtag.managementReadData[5] ),
    .A2(net1305),
    .B1(net1197),
    .B2(net242),
    .C1(net1730),
    .X(_03295_));
 sky130_fd_sc_hd__o21a_4 _16865_ (.A1(net1714),
    .A2(\core.pipe1_resultRegister[5] ),
    .B1(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__mux2_1 _16866_ (.A0(\core.csr.mconfigptr.currentValue[5] ),
    .A1(_03296_),
    .S(net629),
    .X(_03297_));
 sky130_fd_sc_hd__and2_1 _16867_ (.A(net1852),
    .B(_03297_),
    .X(_01543_));
 sky130_fd_sc_hd__a221o_1 _16868_ (.A1(\jtag.managementReadData[6] ),
    .A2(net1305),
    .B1(net1197),
    .B2(net243),
    .C1(net1730),
    .X(_03298_));
 sky130_fd_sc_hd__o21a_4 _16869_ (.A1(net1715),
    .A2(\core.pipe1_resultRegister[6] ),
    .B1(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__inv_2 _16870_ (.A(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__mux2_1 _16871_ (.A0(\core.csr.mconfigptr.currentValue[6] ),
    .A1(_03299_),
    .S(net627),
    .X(_03301_));
 sky130_fd_sc_hd__and2_1 _16872_ (.A(net1851),
    .B(_03301_),
    .X(_01544_));
 sky130_fd_sc_hd__a221o_1 _16873_ (.A1(\jtag.managementReadData[7] ),
    .A2(net1305),
    .B1(net1197),
    .B2(net244),
    .C1(net1729),
    .X(_03302_));
 sky130_fd_sc_hd__o21a_4 _16874_ (.A1(net1715),
    .A2(\core.pipe1_resultRegister[7] ),
    .B1(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__mux2_1 _16875_ (.A0(\core.csr.mconfigptr.currentValue[7] ),
    .A1(_03303_),
    .S(net629),
    .X(_03304_));
 sky130_fd_sc_hd__and2_1 _16876_ (.A(net1852),
    .B(_03304_),
    .X(_01545_));
 sky130_fd_sc_hd__a221o_1 _16877_ (.A1(\jtag.managementReadData[8] ),
    .A2(net1305),
    .B1(net1197),
    .B2(net245),
    .C1(net1729),
    .X(_03305_));
 sky130_fd_sc_hd__o21a_4 _16878_ (.A1(net1716),
    .A2(\core.pipe1_resultRegister[8] ),
    .B1(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__mux2_1 _16879_ (.A0(\core.csr.mconfigptr.currentValue[8] ),
    .A1(_03306_),
    .S(net626),
    .X(_03307_));
 sky130_fd_sc_hd__and2_1 _16880_ (.A(net1850),
    .B(_03307_),
    .X(_01546_));
 sky130_fd_sc_hd__a221o_1 _16881_ (.A1(\jtag.managementReadData[9] ),
    .A2(net1304),
    .B1(net1196),
    .B2(net246),
    .C1(net1729),
    .X(_03308_));
 sky130_fd_sc_hd__o21a_4 _16882_ (.A1(net1718),
    .A2(\core.pipe1_resultRegister[9] ),
    .B1(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__mux2_1 _16883_ (.A0(\core.csr.mconfigptr.currentValue[9] ),
    .A1(_03309_),
    .S(net629),
    .X(_03310_));
 sky130_fd_sc_hd__and2_1 _16884_ (.A(net1864),
    .B(_03310_),
    .X(_01547_));
 sky130_fd_sc_hd__a221o_1 _16885_ (.A1(\jtag.managementReadData[10] ),
    .A2(net1304),
    .B1(net1196),
    .B2(net216),
    .C1(net1729),
    .X(_03311_));
 sky130_fd_sc_hd__o21a_4 _16886_ (.A1(net1718),
    .A2(\core.pipe1_resultRegister[10] ),
    .B1(_03311_),
    .X(_03312_));
 sky130_fd_sc_hd__mux2_1 _16887_ (.A0(\core.csr.mconfigptr.currentValue[10] ),
    .A1(_03312_),
    .S(net629),
    .X(_03313_));
 sky130_fd_sc_hd__and2_1 _16888_ (.A(net1864),
    .B(_03313_),
    .X(_01548_));
 sky130_fd_sc_hd__a221o_1 _16889_ (.A1(\jtag.managementReadData[11] ),
    .A2(net1304),
    .B1(net1196),
    .B2(net217),
    .C1(net1729),
    .X(_03314_));
 sky130_fd_sc_hd__o21a_4 _16890_ (.A1(net1717),
    .A2(\core.pipe1_resultRegister[11] ),
    .B1(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__mux2_1 _16891_ (.A0(\core.csr.mconfigptr.currentValue[11] ),
    .A1(_03315_),
    .S(net629),
    .X(_03316_));
 sky130_fd_sc_hd__and2_1 _16892_ (.A(net1852),
    .B(_03316_),
    .X(_01549_));
 sky130_fd_sc_hd__a221o_1 _16893_ (.A1(\jtag.managementReadData[12] ),
    .A2(net1304),
    .B1(net1196),
    .B2(net218),
    .C1(net1729),
    .X(_03317_));
 sky130_fd_sc_hd__o21a_4 _16894_ (.A1(net1717),
    .A2(\core.pipe1_resultRegister[12] ),
    .B1(_03317_),
    .X(_03318_));
 sky130_fd_sc_hd__mux2_1 _16895_ (.A0(\core.csr.mconfigptr.currentValue[12] ),
    .A1(_03318_),
    .S(net629),
    .X(_03319_));
 sky130_fd_sc_hd__and2_1 _16896_ (.A(net1853),
    .B(_03319_),
    .X(_01550_));
 sky130_fd_sc_hd__a221o_1 _16897_ (.A1(\jtag.managementReadData[13] ),
    .A2(net1303),
    .B1(net1195),
    .B2(net219),
    .C1(net1730),
    .X(_03320_));
 sky130_fd_sc_hd__o21a_4 _16898_ (.A1(net1718),
    .A2(\core.pipe1_resultRegister[13] ),
    .B1(_03320_),
    .X(_03321_));
 sky130_fd_sc_hd__mux2_1 _16899_ (.A0(\core.csr.mconfigptr.currentValue[13] ),
    .A1(_03321_),
    .S(net630),
    .X(_03322_));
 sky130_fd_sc_hd__and2_1 _16900_ (.A(net1854),
    .B(_03322_),
    .X(_01551_));
 sky130_fd_sc_hd__a221o_1 _16901_ (.A1(\jtag.managementReadData[14] ),
    .A2(net1303),
    .B1(net1195),
    .B2(net220),
    .C1(net1728),
    .X(_03323_));
 sky130_fd_sc_hd__o21a_4 _16902_ (.A1(net1717),
    .A2(\core.pipe1_resultRegister[14] ),
    .B1(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__mux2_1 _16903_ (.A0(\core.csr.mconfigptr.currentValue[14] ),
    .A1(_03324_),
    .S(net629),
    .X(_03325_));
 sky130_fd_sc_hd__and2_1 _16904_ (.A(net1853),
    .B(_03325_),
    .X(_01552_));
 sky130_fd_sc_hd__a221o_2 _16905_ (.A1(\jtag.managementReadData[15] ),
    .A2(net1303),
    .B1(net1195),
    .B2(net221),
    .C1(net1728),
    .X(_03326_));
 sky130_fd_sc_hd__o21a_4 _16906_ (.A1(net1715),
    .A2(\core.pipe1_resultRegister[15] ),
    .B1(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__mux2_1 _16907_ (.A0(\core.csr.mconfigptr.currentValue[15] ),
    .A1(_03327_),
    .S(net630),
    .X(_03328_));
 sky130_fd_sc_hd__and2_1 _16908_ (.A(net1854),
    .B(_03328_),
    .X(_01553_));
 sky130_fd_sc_hd__a221o_2 _16909_ (.A1(\jtag.managementReadData[16] ),
    .A2(net1303),
    .B1(net1195),
    .B2(net222),
    .C1(net1728),
    .X(_03329_));
 sky130_fd_sc_hd__o21a_4 _16910_ (.A1(net1715),
    .A2(\core.pipe1_resultRegister[16] ),
    .B1(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__mux2_1 _16911_ (.A0(\core.csr.mconfigptr.currentValue[16] ),
    .A1(_03330_),
    .S(net628),
    .X(_03331_));
 sky130_fd_sc_hd__and2_1 _16912_ (.A(net1854),
    .B(_03331_),
    .X(_01554_));
 sky130_fd_sc_hd__a221o_2 _16913_ (.A1(\jtag.managementReadData[17] ),
    .A2(net1302),
    .B1(net1195),
    .B2(net223),
    .C1(net1728),
    .X(_03332_));
 sky130_fd_sc_hd__o21a_4 _16914_ (.A1(net1715),
    .A2(\core.pipe1_resultRegister[17] ),
    .B1(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_1 _16915_ (.A0(\core.csr.mconfigptr.currentValue[17] ),
    .A1(_03333_),
    .S(net626),
    .X(_03334_));
 sky130_fd_sc_hd__and2_1 _16916_ (.A(net1851),
    .B(_03334_),
    .X(_01555_));
 sky130_fd_sc_hd__a221o_1 _16917_ (.A1(\jtag.managementReadData[18] ),
    .A2(net1301),
    .B1(net1194),
    .B2(net224),
    .C1(net1728),
    .X(_03335_));
 sky130_fd_sc_hd__o21a_4 _16918_ (.A1(net1717),
    .A2(\core.pipe1_resultRegister[18] ),
    .B1(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__mux2_1 _16919_ (.A0(\core.csr.mconfigptr.currentValue[18] ),
    .A1(_03336_),
    .S(net627),
    .X(_03337_));
 sky130_fd_sc_hd__and2_1 _16920_ (.A(net1850),
    .B(_03337_),
    .X(_01556_));
 sky130_fd_sc_hd__a221o_2 _16921_ (.A1(\jtag.managementReadData[19] ),
    .A2(net1302),
    .B1(net1195),
    .B2(net225),
    .C1(net1727),
    .X(_03338_));
 sky130_fd_sc_hd__o21a_4 _16922_ (.A1(net1714),
    .A2(\core.pipe1_resultRegister[19] ),
    .B1(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_1 _16923_ (.A0(\core.csr.mconfigptr.currentValue[19] ),
    .A1(_03339_),
    .S(net627),
    .X(_03340_));
 sky130_fd_sc_hd__and2_1 _16924_ (.A(net1851),
    .B(_03340_),
    .X(_01557_));
 sky130_fd_sc_hd__a221o_2 _16925_ (.A1(\jtag.managementReadData[20] ),
    .A2(net1301),
    .B1(net1194),
    .B2(net227),
    .C1(net1727),
    .X(_03341_));
 sky130_fd_sc_hd__o21a_4 _16926_ (.A1(net1715),
    .A2(\core.pipe1_resultRegister[20] ),
    .B1(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_1 _16927_ (.A0(\core.csr.mconfigptr.currentValue[20] ),
    .A1(_03342_),
    .S(net627),
    .X(_03343_));
 sky130_fd_sc_hd__and2_1 _16928_ (.A(net1851),
    .B(_03343_),
    .X(_01558_));
 sky130_fd_sc_hd__a221o_4 _16929_ (.A1(\jtag.managementReadData[21] ),
    .A2(net1302),
    .B1(net1195),
    .B2(net228),
    .C1(net1728),
    .X(_03344_));
 sky130_fd_sc_hd__o21a_4 _16930_ (.A1(net1713),
    .A2(\core.pipe1_resultRegister[21] ),
    .B1(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _16931_ (.A0(\core.csr.mconfigptr.currentValue[21] ),
    .A1(_03345_),
    .S(net628),
    .X(_03346_));
 sky130_fd_sc_hd__and2_1 _16932_ (.A(net1848),
    .B(_03346_),
    .X(_01559_));
 sky130_fd_sc_hd__a221o_4 _16933_ (.A1(\jtag.managementReadData[22] ),
    .A2(net1301),
    .B1(net1194),
    .B2(net229),
    .C1(net1727),
    .X(_03347_));
 sky130_fd_sc_hd__o21a_4 _16934_ (.A1(net1714),
    .A2(\core.pipe1_resultRegister[22] ),
    .B1(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_1 _16935_ (.A0(\core.csr.mconfigptr.currentValue[22] ),
    .A1(_03348_),
    .S(net628),
    .X(_03349_));
 sky130_fd_sc_hd__and2_1 _16936_ (.A(net1849),
    .B(_03349_),
    .X(_01560_));
 sky130_fd_sc_hd__a221o_4 _16937_ (.A1(\jtag.managementReadData[23] ),
    .A2(net1301),
    .B1(net1194),
    .B2(net230),
    .C1(net1727),
    .X(_03350_));
 sky130_fd_sc_hd__o21a_4 _16938_ (.A1(net1714),
    .A2(\core.pipe1_resultRegister[23] ),
    .B1(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__mux2_1 _16939_ (.A0(\core.csr.mconfigptr.currentValue[23] ),
    .A1(_03351_),
    .S(net628),
    .X(_03352_));
 sky130_fd_sc_hd__and2_1 _16940_ (.A(net1848),
    .B(_03352_),
    .X(_01561_));
 sky130_fd_sc_hd__a221o_2 _16941_ (.A1(\jtag.managementReadData[24] ),
    .A2(net1301),
    .B1(net1194),
    .B2(net231),
    .C1(net1727),
    .X(_03353_));
 sky130_fd_sc_hd__o21a_4 _16942_ (.A1(net1715),
    .A2(\core.pipe1_resultRegister[24] ),
    .B1(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__mux2_1 _16943_ (.A0(\core.csr.mconfigptr.currentValue[24] ),
    .A1(_03354_),
    .S(net628),
    .X(_03355_));
 sky130_fd_sc_hd__and2_1 _16944_ (.A(net1854),
    .B(_03355_),
    .X(_01562_));
 sky130_fd_sc_hd__a221o_2 _16945_ (.A1(\jtag.managementReadData[25] ),
    .A2(net1301),
    .B1(net1194),
    .B2(net232),
    .C1(net1727),
    .X(_03356_));
 sky130_fd_sc_hd__o21a_4 _16946_ (.A1(net1715),
    .A2(\core.pipe1_resultRegister[25] ),
    .B1(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__mux2_1 _16947_ (.A0(\core.csr.mconfigptr.currentValue[25] ),
    .A1(_03357_),
    .S(net628),
    .X(_03358_));
 sky130_fd_sc_hd__and2_1 _16948_ (.A(net1854),
    .B(_03358_),
    .X(_01563_));
 sky130_fd_sc_hd__a221o_2 _16949_ (.A1(\jtag.managementReadData[26] ),
    .A2(net1301),
    .B1(net1194),
    .B2(net233),
    .C1(net1727),
    .X(_03359_));
 sky130_fd_sc_hd__o21a_4 _16950_ (.A1(net1717),
    .A2(\core.pipe1_resultRegister[26] ),
    .B1(_03359_),
    .X(_03360_));
 sky130_fd_sc_hd__mux2_1 _16951_ (.A0(\core.csr.mconfigptr.currentValue[26] ),
    .A1(_03360_),
    .S(net629),
    .X(_03361_));
 sky130_fd_sc_hd__and2_1 _16952_ (.A(net1854),
    .B(_03361_),
    .X(_01564_));
 sky130_fd_sc_hd__a221o_1 _16953_ (.A1(\jtag.managementReadData[27] ),
    .A2(net1301),
    .B1(net1194),
    .B2(net234),
    .C1(net1727),
    .X(_03362_));
 sky130_fd_sc_hd__o21a_4 _16954_ (.A1(net1717),
    .A2(\core.pipe1_resultRegister[27] ),
    .B1(_03362_),
    .X(_03363_));
 sky130_fd_sc_hd__mux2_1 _16955_ (.A0(\core.csr.mconfigptr.currentValue[27] ),
    .A1(_03363_),
    .S(net630),
    .X(_03364_));
 sky130_fd_sc_hd__and2_1 _16956_ (.A(net1854),
    .B(_03364_),
    .X(_01565_));
 sky130_fd_sc_hd__a221o_1 _16957_ (.A1(\jtag.managementReadData[28] ),
    .A2(net1301),
    .B1(net1194),
    .B2(net235),
    .C1(net1727),
    .X(_03365_));
 sky130_fd_sc_hd__o21a_4 _16958_ (.A1(net1717),
    .A2(\core.pipe1_resultRegister[28] ),
    .B1(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__mux2_1 _16959_ (.A0(\core.csr.mconfigptr.currentValue[28] ),
    .A1(_03366_),
    .S(net630),
    .X(_03367_));
 sky130_fd_sc_hd__and2_1 _16960_ (.A(net1854),
    .B(_03367_),
    .X(_01566_));
 sky130_fd_sc_hd__a221o_1 _16961_ (.A1(\jtag.managementReadData[29] ),
    .A2(net1303),
    .B1(net1195),
    .B2(net236),
    .C1(net1728),
    .X(_03368_));
 sky130_fd_sc_hd__o21a_4 _16962_ (.A1(net1717),
    .A2(\core.pipe1_resultRegister[29] ),
    .B1(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__mux2_1 _16963_ (.A0(\core.csr.mconfigptr.currentValue[29] ),
    .A1(_03369_),
    .S(net630),
    .X(_03370_));
 sky130_fd_sc_hd__and2_1 _16964_ (.A(net1865),
    .B(_03370_),
    .X(_01567_));
 sky130_fd_sc_hd__a221o_1 _16965_ (.A1(\jtag.managementReadData[30] ),
    .A2(net1301),
    .B1(net1194),
    .B2(net238),
    .C1(net1727),
    .X(_03371_));
 sky130_fd_sc_hd__o21a_4 _16966_ (.A1(net1717),
    .A2(\core.pipe1_resultRegister[30] ),
    .B1(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__mux2_1 _16967_ (.A0(\core.csr.mconfigptr.currentValue[30] ),
    .A1(_03372_),
    .S(net626),
    .X(_03373_));
 sky130_fd_sc_hd__and2_1 _16968_ (.A(net1850),
    .B(_03373_),
    .X(_01568_));
 sky130_fd_sc_hd__a221o_1 _16969_ (.A1(\jtag.managementReadData[31] ),
    .A2(net1302),
    .B1(net1195),
    .B2(net239),
    .C1(net1728),
    .X(_03374_));
 sky130_fd_sc_hd__o21a_4 _16970_ (.A1(net1717),
    .A2(\core.pipe1_resultRegister[31] ),
    .B1(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__mux2_1 _16971_ (.A0(\core.csr.mconfigptr.currentValue[31] ),
    .A1(_03375_),
    .S(net629),
    .X(_03376_));
 sky130_fd_sc_hd__and2_1 _16972_ (.A(net1864),
    .B(_03376_),
    .X(_01569_));
 sky130_fd_sc_hd__or2_4 _16973_ (.A(_03262_),
    .B(_03263_),
    .X(_03377_));
 sky130_fd_sc_hd__or3_1 _16974_ (.A(_03271_),
    .B(_03272_),
    .C(_03273_),
    .X(_03378_));
 sky130_fd_sc_hd__or3_2 _16975_ (.A(_03267_),
    .B(_03270_),
    .C(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__clkinv_2 _16976_ (.A(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand2_8 _16977_ (.A(_03261_),
    .B(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__or3b_4 _16978_ (.A(_03259_),
    .B(_03381_),
    .C_N(_03258_),
    .X(_03382_));
 sky130_fd_sc_hd__inv_2 _16979_ (.A(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__or2_4 _16980_ (.A(_03377_),
    .B(_03382_),
    .X(_03384_));
 sky130_fd_sc_hd__or3b_4 _16981_ (.A(_03275_),
    .B(_03259_),
    .C_N(_03257_),
    .X(_03385_));
 sky130_fd_sc_hd__nor3_4 _16982_ (.A(_03377_),
    .B(_03381_),
    .C(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__or2_1 _16983_ (.A(\core.csr.traps.mscratch.currentValue[0] ),
    .B(net652),
    .X(_03387_));
 sky130_fd_sc_hd__o211a_1 _16984_ (.A1(_03281_),
    .A2(net624),
    .B1(_03387_),
    .C1(net1845),
    .X(_01570_));
 sky130_fd_sc_hd__or2_1 _16985_ (.A(\core.csr.traps.mscratch.currentValue[1] ),
    .B(net652),
    .X(_03388_));
 sky130_fd_sc_hd__o211a_1 _16986_ (.A1(_03284_),
    .A2(net624),
    .B1(_03388_),
    .C1(net1844),
    .X(_01571_));
 sky130_fd_sc_hd__or2_1 _16987_ (.A(\core.csr.traps.mscratch.currentValue[2] ),
    .B(net652),
    .X(_03389_));
 sky130_fd_sc_hd__o211a_1 _16988_ (.A1(_03287_),
    .A2(net624),
    .B1(_03389_),
    .C1(net1845),
    .X(_01572_));
 sky130_fd_sc_hd__nand2_1 _16989_ (.A(_03290_),
    .B(net652),
    .Y(_03390_));
 sky130_fd_sc_hd__o211a_1 _16990_ (.A1(\core.csr.traps.mscratch.currentValue[3] ),
    .A2(net652),
    .B1(_03390_),
    .C1(net1845),
    .X(_01573_));
 sky130_fd_sc_hd__or2_1 _16991_ (.A(\core.csr.traps.mscratch.currentValue[4] ),
    .B(net653),
    .X(_03391_));
 sky130_fd_sc_hd__o211a_1 _16992_ (.A1(_03293_),
    .A2(net625),
    .B1(_03391_),
    .C1(net1829),
    .X(_01574_));
 sky130_fd_sc_hd__or2_1 _16993_ (.A(\core.csr.traps.mscratch.currentValue[5] ),
    .B(net652),
    .X(_03392_));
 sky130_fd_sc_hd__o211a_1 _16994_ (.A1(_03296_),
    .A2(net624),
    .B1(_03392_),
    .C1(net1846),
    .X(_01575_));
 sky130_fd_sc_hd__or2_1 _16995_ (.A(\core.csr.traps.mscratch.currentValue[6] ),
    .B(net652),
    .X(_03393_));
 sky130_fd_sc_hd__o211a_1 _16996_ (.A1(_03299_),
    .A2(net624),
    .B1(_03393_),
    .C1(net1847),
    .X(_01576_));
 sky130_fd_sc_hd__or2_1 _16997_ (.A(\core.csr.traps.mscratch.currentValue[7] ),
    .B(net652),
    .X(_03394_));
 sky130_fd_sc_hd__o211a_1 _16998_ (.A1(_03303_),
    .A2(net624),
    .B1(_03394_),
    .C1(net1847),
    .X(_01577_));
 sky130_fd_sc_hd__or2_1 _16999_ (.A(\core.csr.traps.mscratch.currentValue[8] ),
    .B(net653),
    .X(_03395_));
 sky130_fd_sc_hd__o211a_1 _17000_ (.A1(_03306_),
    .A2(net625),
    .B1(_03395_),
    .C1(net1847),
    .X(_01578_));
 sky130_fd_sc_hd__or2_1 _17001_ (.A(\core.csr.traps.mscratch.currentValue[9] ),
    .B(net651),
    .X(_03396_));
 sky130_fd_sc_hd__o211a_1 _17002_ (.A1(_03309_),
    .A2(net623),
    .B1(_03396_),
    .C1(net1827),
    .X(_01579_));
 sky130_fd_sc_hd__or2_1 _17003_ (.A(\core.csr.traps.mscratch.currentValue[10] ),
    .B(_03386_),
    .X(_03397_));
 sky130_fd_sc_hd__o211a_1 _17004_ (.A1(_03312_),
    .A2(net625),
    .B1(_03397_),
    .C1(net1831),
    .X(_01580_));
 sky130_fd_sc_hd__or2_1 _17005_ (.A(\core.csr.traps.mscratch.currentValue[11] ),
    .B(net653),
    .X(_03398_));
 sky130_fd_sc_hd__o211a_1 _17006_ (.A1(_03315_),
    .A2(net624),
    .B1(_03398_),
    .C1(net1848),
    .X(_01581_));
 sky130_fd_sc_hd__or2_1 _17007_ (.A(\core.csr.traps.mscratch.currentValue[12] ),
    .B(net653),
    .X(_03399_));
 sky130_fd_sc_hd__o211a_1 _17008_ (.A1(_03318_),
    .A2(net625),
    .B1(_03399_),
    .C1(net1849),
    .X(_01582_));
 sky130_fd_sc_hd__or2_1 _17009_ (.A(\core.csr.traps.mscratch.currentValue[13] ),
    .B(net653),
    .X(_03400_));
 sky130_fd_sc_hd__o211a_1 _17010_ (.A1(_03321_),
    .A2(net624),
    .B1(_03400_),
    .C1(net1847),
    .X(_01583_));
 sky130_fd_sc_hd__or2_1 _17011_ (.A(\core.csr.traps.mscratch.currentValue[14] ),
    .B(net652),
    .X(_03401_));
 sky130_fd_sc_hd__o211a_1 _17012_ (.A1(_03324_),
    .A2(net624),
    .B1(_03401_),
    .C1(net1848),
    .X(_01584_));
 sky130_fd_sc_hd__or2_1 _17013_ (.A(\core.csr.traps.mscratch.currentValue[15] ),
    .B(net651),
    .X(_03402_));
 sky130_fd_sc_hd__o211a_1 _17014_ (.A1(_03327_),
    .A2(net623),
    .B1(_03402_),
    .C1(net1828),
    .X(_01585_));
 sky130_fd_sc_hd__or2_1 _17015_ (.A(\core.csr.traps.mscratch.currentValue[16] ),
    .B(net651),
    .X(_03403_));
 sky130_fd_sc_hd__o211a_1 _17016_ (.A1(_03330_),
    .A2(net623),
    .B1(_03403_),
    .C1(net1828),
    .X(_01586_));
 sky130_fd_sc_hd__or2_1 _17017_ (.A(\core.csr.traps.mscratch.currentValue[17] ),
    .B(net651),
    .X(_03404_));
 sky130_fd_sc_hd__o211a_1 _17018_ (.A1(_03333_),
    .A2(net623),
    .B1(_03404_),
    .C1(net1825),
    .X(_01587_));
 sky130_fd_sc_hd__or2_1 _17019_ (.A(\core.csr.traps.mscratch.currentValue[18] ),
    .B(net650),
    .X(_03405_));
 sky130_fd_sc_hd__o211a_1 _17020_ (.A1(_03336_),
    .A2(net622),
    .B1(_03405_),
    .C1(net1815),
    .X(_01588_));
 sky130_fd_sc_hd__or2_1 _17021_ (.A(\core.csr.traps.mscratch.currentValue[19] ),
    .B(net650),
    .X(_03406_));
 sky130_fd_sc_hd__o211a_1 _17022_ (.A1(_03339_),
    .A2(net622),
    .B1(_03406_),
    .C1(net1815),
    .X(_01589_));
 sky130_fd_sc_hd__or2_1 _17023_ (.A(\core.csr.traps.mscratch.currentValue[20] ),
    .B(net650),
    .X(_03407_));
 sky130_fd_sc_hd__o211a_1 _17024_ (.A1(_03342_),
    .A2(net622),
    .B1(_03407_),
    .C1(net1810),
    .X(_01590_));
 sky130_fd_sc_hd__or2_1 _17025_ (.A(\core.csr.traps.mscratch.currentValue[21] ),
    .B(net651),
    .X(_03408_));
 sky130_fd_sc_hd__o211a_1 _17026_ (.A1(_03345_),
    .A2(net623),
    .B1(_03408_),
    .C1(net1828),
    .X(_01591_));
 sky130_fd_sc_hd__or2_1 _17027_ (.A(\core.csr.traps.mscratch.currentValue[22] ),
    .B(net651),
    .X(_03409_));
 sky130_fd_sc_hd__o211a_1 _17028_ (.A1(_03348_),
    .A2(net623),
    .B1(_03409_),
    .C1(net1818),
    .X(_01592_));
 sky130_fd_sc_hd__or2_1 _17029_ (.A(\core.csr.traps.mscratch.currentValue[23] ),
    .B(net650),
    .X(_03410_));
 sky130_fd_sc_hd__o211a_1 _17030_ (.A1(_03351_),
    .A2(net622),
    .B1(_03410_),
    .C1(net1817),
    .X(_01593_));
 sky130_fd_sc_hd__or2_1 _17031_ (.A(\core.csr.traps.mscratch.currentValue[24] ),
    .B(net650),
    .X(_03411_));
 sky130_fd_sc_hd__o211a_1 _17032_ (.A1(_03354_),
    .A2(net623),
    .B1(_03411_),
    .C1(net1819),
    .X(_01594_));
 sky130_fd_sc_hd__or2_1 _17033_ (.A(\core.csr.traps.mscratch.currentValue[25] ),
    .B(net650),
    .X(_03412_));
 sky130_fd_sc_hd__o211a_1 _17034_ (.A1(_03357_),
    .A2(net622),
    .B1(_03412_),
    .C1(net1817),
    .X(_01595_));
 sky130_fd_sc_hd__or2_1 _17035_ (.A(\core.csr.traps.mscratch.currentValue[26] ),
    .B(net650),
    .X(_03413_));
 sky130_fd_sc_hd__o211a_1 _17036_ (.A1(_03360_),
    .A2(net622),
    .B1(_03413_),
    .C1(net1817),
    .X(_01596_));
 sky130_fd_sc_hd__or2_1 _17037_ (.A(\core.csr.traps.mscratch.currentValue[27] ),
    .B(net650),
    .X(_03414_));
 sky130_fd_sc_hd__o211a_1 _17038_ (.A1(_03363_),
    .A2(net622),
    .B1(_03414_),
    .C1(net1818),
    .X(_01597_));
 sky130_fd_sc_hd__or2_1 _17039_ (.A(\core.csr.traps.mscratch.currentValue[28] ),
    .B(net650),
    .X(_03415_));
 sky130_fd_sc_hd__o211a_1 _17040_ (.A1(_03366_),
    .A2(net622),
    .B1(_03415_),
    .C1(net1813),
    .X(_01598_));
 sky130_fd_sc_hd__or2_1 _17041_ (.A(\core.csr.traps.mscratch.currentValue[29] ),
    .B(net650),
    .X(_03416_));
 sky130_fd_sc_hd__o211a_1 _17042_ (.A1(_03369_),
    .A2(net622),
    .B1(_03416_),
    .C1(net1813),
    .X(_01599_));
 sky130_fd_sc_hd__or2_1 _17043_ (.A(\core.csr.traps.mscratch.currentValue[30] ),
    .B(net652),
    .X(_03417_));
 sky130_fd_sc_hd__o211a_1 _17044_ (.A1(_03372_),
    .A2(net624),
    .B1(_03417_),
    .C1(net1845),
    .X(_01600_));
 sky130_fd_sc_hd__or2_1 _17045_ (.A(\core.csr.traps.mscratch.currentValue[31] ),
    .B(net651),
    .X(_03418_));
 sky130_fd_sc_hd__o211a_1 _17046_ (.A1(_03375_),
    .A2(net622),
    .B1(_03418_),
    .C1(net1815),
    .X(_01601_));
 sky130_fd_sc_hd__or2_4 _17047_ (.A(_03261_),
    .B(_03379_),
    .X(_03419_));
 sky130_fd_sc_hd__or2_4 _17048_ (.A(_03260_),
    .B(_03377_),
    .X(_03420_));
 sky130_fd_sc_hd__nor2_8 _17049_ (.A(_03419_),
    .B(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hd__or2_4 _17050_ (.A(_03419_),
    .B(_03420_),
    .X(_03422_));
 sky130_fd_sc_hd__or4_1 _17051_ (.A(_03261_),
    .B(_03268_),
    .C(_03269_),
    .D(_03271_),
    .X(_03423_));
 sky130_fd_sc_hd__or4_4 _17052_ (.A(_03267_),
    .B(_03272_),
    .C(_03273_),
    .D(_03423_),
    .X(_03424_));
 sky130_fd_sc_hd__or2_1 _17053_ (.A(\core.csr.traps.mie.currentValue[0] ),
    .B(net648),
    .X(_03425_));
 sky130_fd_sc_hd__o211a_1 _17054_ (.A1(_03281_),
    .A2(net644),
    .B1(_03425_),
    .C1(net1845),
    .X(_01602_));
 sky130_fd_sc_hd__or2_1 _17055_ (.A(\core.csr.traps.mie.currentValue[1] ),
    .B(net648),
    .X(_03426_));
 sky130_fd_sc_hd__o211a_1 _17056_ (.A1(_03284_),
    .A2(net645),
    .B1(_03426_),
    .C1(net1845),
    .X(_01603_));
 sky130_fd_sc_hd__or2_1 _17057_ (.A(\core.csr.traps.mie.currentValue[2] ),
    .B(net648),
    .X(_03427_));
 sky130_fd_sc_hd__o211a_1 _17058_ (.A1(_03287_),
    .A2(net644),
    .B1(_03427_),
    .C1(net1845),
    .X(_01604_));
 sky130_fd_sc_hd__nand2_1 _17059_ (.A(_03290_),
    .B(net648),
    .Y(_03428_));
 sky130_fd_sc_hd__o211a_1 _17060_ (.A1(\core.csr.traps.mie.currentValue[3] ),
    .A2(net648),
    .B1(_03428_),
    .C1(net1850),
    .X(_01605_));
 sky130_fd_sc_hd__or2_1 _17061_ (.A(\core.csr.traps.mie.currentValue[4] ),
    .B(_03421_),
    .X(_03429_));
 sky130_fd_sc_hd__o211a_1 _17062_ (.A1(_03293_),
    .A2(net645),
    .B1(_03429_),
    .C1(net1846),
    .X(_01606_));
 sky130_fd_sc_hd__or2_1 _17063_ (.A(\core.csr.traps.mie.currentValue[5] ),
    .B(net648),
    .X(_03430_));
 sky130_fd_sc_hd__o211a_1 _17064_ (.A1(_03296_),
    .A2(net644),
    .B1(_03430_),
    .C1(net1845),
    .X(_01607_));
 sky130_fd_sc_hd__or2_1 _17065_ (.A(\core.csr.traps.mie.currentValue[6] ),
    .B(net649),
    .X(_03431_));
 sky130_fd_sc_hd__o211a_1 _17066_ (.A1(_03299_),
    .A2(net645),
    .B1(_03431_),
    .C1(net1848),
    .X(_01608_));
 sky130_fd_sc_hd__or2_1 _17067_ (.A(\core.csr.traps.mie.currentValue[7] ),
    .B(net649),
    .X(_03432_));
 sky130_fd_sc_hd__o211a_1 _17068_ (.A1(_03303_),
    .A2(net644),
    .B1(_03432_),
    .C1(net1847),
    .X(_01609_));
 sky130_fd_sc_hd__or2_1 _17069_ (.A(\core.csr.traps.mie.currentValue[8] ),
    .B(net649),
    .X(_03433_));
 sky130_fd_sc_hd__o211a_1 _17070_ (.A1(_03306_),
    .A2(net644),
    .B1(_03433_),
    .C1(net1847),
    .X(_01610_));
 sky130_fd_sc_hd__or2_1 _17071_ (.A(\core.csr.traps.mie.currentValue[9] ),
    .B(net647),
    .X(_03434_));
 sky130_fd_sc_hd__o211a_1 _17072_ (.A1(_03309_),
    .A2(net643),
    .B1(_03434_),
    .C1(net1827),
    .X(_01611_));
 sky130_fd_sc_hd__or2_1 _17073_ (.A(\core.csr.traps.mie.currentValue[10] ),
    .B(_03421_),
    .X(_03435_));
 sky130_fd_sc_hd__o211a_1 _17074_ (.A1(_03312_),
    .A2(net645),
    .B1(_03435_),
    .C1(net1831),
    .X(_01612_));
 sky130_fd_sc_hd__or2_1 _17075_ (.A(\core.csr.traps.mie.currentValue[11] ),
    .B(net648),
    .X(_03436_));
 sky130_fd_sc_hd__o211a_1 _17076_ (.A1(_03315_),
    .A2(net644),
    .B1(_03436_),
    .C1(net1848),
    .X(_01613_));
 sky130_fd_sc_hd__or2_1 _17077_ (.A(\core.csr.traps.mie.currentValue[12] ),
    .B(net649),
    .X(_03437_));
 sky130_fd_sc_hd__o211a_1 _17078_ (.A1(_03318_),
    .A2(net644),
    .B1(_03437_),
    .C1(net1848),
    .X(_01614_));
 sky130_fd_sc_hd__or2_1 _17079_ (.A(\core.csr.traps.mie.currentValue[13] ),
    .B(net648),
    .X(_03438_));
 sky130_fd_sc_hd__o211a_1 _17080_ (.A1(_03321_),
    .A2(net644),
    .B1(_03438_),
    .C1(net1848),
    .X(_01615_));
 sky130_fd_sc_hd__or2_1 _17081_ (.A(\core.csr.traps.mie.currentValue[14] ),
    .B(net648),
    .X(_03439_));
 sky130_fd_sc_hd__o211a_1 _17082_ (.A1(_03324_),
    .A2(net644),
    .B1(_03439_),
    .C1(net1848),
    .X(_01616_));
 sky130_fd_sc_hd__or2_1 _17083_ (.A(\core.csr.traps.mie.currentValue[15] ),
    .B(net647),
    .X(_03440_));
 sky130_fd_sc_hd__o211a_1 _17084_ (.A1(_03327_),
    .A2(net643),
    .B1(_03440_),
    .C1(net1828),
    .X(_01617_));
 sky130_fd_sc_hd__or2_1 _17085_ (.A(\core.csr.traps.mie.currentValue[16] ),
    .B(net646),
    .X(_03441_));
 sky130_fd_sc_hd__o211a_1 _17086_ (.A1(_03330_),
    .A2(net643),
    .B1(_03441_),
    .C1(net1828),
    .X(_01618_));
 sky130_fd_sc_hd__or2_1 _17087_ (.A(\core.csr.traps.mie.currentValue[17] ),
    .B(net647),
    .X(_03442_));
 sky130_fd_sc_hd__o211a_1 _17088_ (.A1(_03333_),
    .A2(net643),
    .B1(_03442_),
    .C1(net1826),
    .X(_01619_));
 sky130_fd_sc_hd__or2_1 _17089_ (.A(\core.csr.traps.mie.currentValue[18] ),
    .B(net646),
    .X(_03443_));
 sky130_fd_sc_hd__o211a_1 _17090_ (.A1(_03336_),
    .A2(net642),
    .B1(_03443_),
    .C1(net1815),
    .X(_01620_));
 sky130_fd_sc_hd__or2_1 _17091_ (.A(\core.csr.traps.mie.currentValue[19] ),
    .B(net646),
    .X(_03444_));
 sky130_fd_sc_hd__o211a_1 _17092_ (.A1(_03339_),
    .A2(net642),
    .B1(_03444_),
    .C1(net1814),
    .X(_01621_));
 sky130_fd_sc_hd__or2_1 _17093_ (.A(\core.csr.traps.mie.currentValue[20] ),
    .B(net646),
    .X(_03445_));
 sky130_fd_sc_hd__o211a_1 _17094_ (.A1(_03342_),
    .A2(net642),
    .B1(_03445_),
    .C1(net1814),
    .X(_01622_));
 sky130_fd_sc_hd__or2_1 _17095_ (.A(\core.csr.traps.mie.currentValue[21] ),
    .B(net647),
    .X(_03446_));
 sky130_fd_sc_hd__o211a_1 _17096_ (.A1(_03345_),
    .A2(net643),
    .B1(_03446_),
    .C1(net1828),
    .X(_01623_));
 sky130_fd_sc_hd__or2_1 _17097_ (.A(\core.csr.traps.mie.currentValue[22] ),
    .B(net647),
    .X(_03447_));
 sky130_fd_sc_hd__o211a_1 _17098_ (.A1(_03348_),
    .A2(net642),
    .B1(_03447_),
    .C1(net1818),
    .X(_01624_));
 sky130_fd_sc_hd__or2_1 _17099_ (.A(\core.csr.traps.mie.currentValue[23] ),
    .B(net646),
    .X(_03448_));
 sky130_fd_sc_hd__o211a_1 _17100_ (.A1(_03351_),
    .A2(net642),
    .B1(_03448_),
    .C1(net1817),
    .X(_01625_));
 sky130_fd_sc_hd__or2_1 _17101_ (.A(\core.csr.traps.mie.currentValue[24] ),
    .B(net647),
    .X(_03449_));
 sky130_fd_sc_hd__o211a_1 _17102_ (.A1(_03354_),
    .A2(net643),
    .B1(_03449_),
    .C1(net1819),
    .X(_01626_));
 sky130_fd_sc_hd__or2_1 _17103_ (.A(\core.csr.traps.mie.currentValue[25] ),
    .B(net646),
    .X(_03450_));
 sky130_fd_sc_hd__o211a_1 _17104_ (.A1(_03357_),
    .A2(net642),
    .B1(_03450_),
    .C1(net1816),
    .X(_01627_));
 sky130_fd_sc_hd__or2_1 _17105_ (.A(\core.csr.traps.mie.currentValue[26] ),
    .B(net646),
    .X(_03451_));
 sky130_fd_sc_hd__o211a_1 _17106_ (.A1(_03360_),
    .A2(net642),
    .B1(_03451_),
    .C1(net1817),
    .X(_01628_));
 sky130_fd_sc_hd__or2_1 _17107_ (.A(\core.csr.traps.mie.currentValue[27] ),
    .B(net647),
    .X(_03452_));
 sky130_fd_sc_hd__o211a_1 _17108_ (.A1(_03363_),
    .A2(net643),
    .B1(_03452_),
    .C1(net1819),
    .X(_01629_));
 sky130_fd_sc_hd__or2_1 _17109_ (.A(\core.csr.traps.mie.currentValue[28] ),
    .B(net646),
    .X(_03453_));
 sky130_fd_sc_hd__o211a_1 _17110_ (.A1(_03366_),
    .A2(net642),
    .B1(_03453_),
    .C1(net1816),
    .X(_01630_));
 sky130_fd_sc_hd__or2_1 _17111_ (.A(\core.csr.traps.mie.currentValue[29] ),
    .B(net646),
    .X(_03454_));
 sky130_fd_sc_hd__o211a_1 _17112_ (.A1(_03369_),
    .A2(net642),
    .B1(_03454_),
    .C1(net1816),
    .X(_01631_));
 sky130_fd_sc_hd__or2_1 _17113_ (.A(\core.csr.traps.mie.currentValue[30] ),
    .B(net648),
    .X(_03455_));
 sky130_fd_sc_hd__o211a_1 _17114_ (.A1(_03372_),
    .A2(net644),
    .B1(_03455_),
    .C1(net1846),
    .X(_01632_));
 sky130_fd_sc_hd__or2_1 _17115_ (.A(\core.csr.traps.mie.currentValue[31] ),
    .B(net646),
    .X(_03456_));
 sky130_fd_sc_hd__o211a_1 _17116_ (.A1(_03375_),
    .A2(net642),
    .B1(_03456_),
    .C1(net1815),
    .X(_01633_));
 sky130_fd_sc_hd__nand2_1 _17117_ (.A(net555),
    .B(_03281_),
    .Y(_03457_));
 sky130_fd_sc_hd__or3b_2 _17118_ (.A(_03382_),
    .B(_03262_),
    .C_N(_03263_),
    .X(_03458_));
 sky130_fd_sc_hd__and2_1 _17119_ (.A(net550),
    .B(net618),
    .X(_03459_));
 sky130_fd_sc_hd__nand2_8 _17120_ (.A(net551),
    .B(net619),
    .Y(_03460_));
 sky130_fd_sc_hd__a31o_1 _17121_ (.A1(_02255_),
    .A2(_03457_),
    .A3(_03460_),
    .B1(net1877),
    .X(_03461_));
 sky130_fd_sc_hd__o21ba_1 _17122_ (.A1(\core.csr.traps.mcause.csrReadData[0] ),
    .A2(_03460_),
    .B1_N(_03461_),
    .X(_01634_));
 sky130_fd_sc_hd__nand2_1 _17123_ (.A(net555),
    .B(_03284_),
    .Y(_03462_));
 sky130_fd_sc_hd__or3b_1 _17124_ (.A(_02257_),
    .B(net535),
    .C_N(_03462_),
    .X(_03463_));
 sky130_fd_sc_hd__o211a_1 _17125_ (.A1(\core.csr.traps.mcause.csrReadData[1] ),
    .A2(_03460_),
    .B1(_03463_),
    .C1(net1830),
    .X(_01635_));
 sky130_fd_sc_hd__nand2_1 _17126_ (.A(net555),
    .B(_03287_),
    .Y(_03464_));
 sky130_fd_sc_hd__a31o_1 _17127_ (.A1(_02254_),
    .A2(_03460_),
    .A3(_03464_),
    .B1(net1877),
    .X(_03465_));
 sky130_fd_sc_hd__o21ba_1 _17128_ (.A1(\core.csr.traps.mcause.csrReadData[2] ),
    .A2(_03460_),
    .B1_N(_03465_),
    .X(_01636_));
 sky130_fd_sc_hd__nor2_2 _17129_ (.A(net545),
    .B(_03290_),
    .Y(_03466_));
 sky130_fd_sc_hd__a21oi_1 _17130_ (.A1(net444),
    .A2(_02253_),
    .B1(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__a31o_1 _17131_ (.A1(net1103),
    .A2(_03460_),
    .A3(_03467_),
    .B1(net1875),
    .X(_03468_));
 sky130_fd_sc_hd__o21ba_1 _17132_ (.A1(\core.csr.traps.mcause.csrReadData[3] ),
    .A2(_03460_),
    .B1_N(_03468_),
    .X(_01637_));
 sky130_fd_sc_hd__nand2_1 _17133_ (.A(net555),
    .B(_03293_),
    .Y(_03469_));
 sky130_fd_sc_hd__o2bb2a_1 _17134_ (.A1_N(\core.csr.traps.mcause.csrReadData[4] ),
    .A2_N(net534),
    .B1(_03469_),
    .B2(net620),
    .X(_03470_));
 sky130_fd_sc_hd__nor2_1 _17135_ (.A(net1877),
    .B(_03470_),
    .Y(_01638_));
 sky130_fd_sc_hd__nand2_1 _17136_ (.A(net555),
    .B(_03296_),
    .Y(_03471_));
 sky130_fd_sc_hd__o2bb2a_1 _17137_ (.A1_N(\core.csr.traps.mcause.csrReadData[5] ),
    .A2_N(net534),
    .B1(_03471_),
    .B2(net620),
    .X(_03472_));
 sky130_fd_sc_hd__nor2_1 _17138_ (.A(net1877),
    .B(_03472_),
    .Y(_01639_));
 sky130_fd_sc_hd__nand2_1 _17139_ (.A(net555),
    .B(_03299_),
    .Y(_03473_));
 sky130_fd_sc_hd__o2bb2a_1 _17140_ (.A1_N(\core.csr.traps.mcause.csrReadData[6] ),
    .A2_N(net534),
    .B1(_03473_),
    .B2(net621),
    .X(_03474_));
 sky130_fd_sc_hd__nor2_1 _17141_ (.A(net1877),
    .B(_03474_),
    .Y(_01640_));
 sky130_fd_sc_hd__nand2_2 _17142_ (.A(net556),
    .B(_03303_),
    .Y(_03475_));
 sky130_fd_sc_hd__o2bb2a_1 _17143_ (.A1_N(\core.csr.traps.mcause.csrReadData[7] ),
    .A2_N(net535),
    .B1(_03475_),
    .B2(net621),
    .X(_03476_));
 sky130_fd_sc_hd__nor2_1 _17144_ (.A(net1878),
    .B(_03476_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_1 _17145_ (.A(net556),
    .B(_03306_),
    .Y(_03477_));
 sky130_fd_sc_hd__o2bb2a_1 _17146_ (.A1_N(\core.csr.traps.mcause.csrReadData[8] ),
    .A2_N(net534),
    .B1(_03477_),
    .B2(net620),
    .X(_03478_));
 sky130_fd_sc_hd__nor2_1 _17147_ (.A(net1878),
    .B(_03478_),
    .Y(_01642_));
 sky130_fd_sc_hd__nand2_1 _17148_ (.A(net553),
    .B(_03309_),
    .Y(_03479_));
 sky130_fd_sc_hd__o2bb2a_1 _17149_ (.A1_N(\core.csr.traps.mcause.csrReadData[9] ),
    .A2_N(net534),
    .B1(_03479_),
    .B2(net620),
    .X(_03480_));
 sky130_fd_sc_hd__nor2_1 _17150_ (.A(net1876),
    .B(_03480_),
    .Y(_01643_));
 sky130_fd_sc_hd__nand2_1 _17151_ (.A(net556),
    .B(_03312_),
    .Y(_03481_));
 sky130_fd_sc_hd__o2bb2a_1 _17152_ (.A1_N(\core.csr.traps.mcause.csrReadData[10] ),
    .A2_N(net535),
    .B1(_03481_),
    .B2(net621),
    .X(_03482_));
 sky130_fd_sc_hd__nor2_1 _17153_ (.A(net1878),
    .B(_03482_),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _17154_ (.A(net555),
    .B(_03315_),
    .Y(_03483_));
 sky130_fd_sc_hd__o2bb2a_1 _17155_ (.A1_N(\core.csr.traps.mcause.csrReadData[11] ),
    .A2_N(net535),
    .B1(_03483_),
    .B2(net620),
    .X(_03484_));
 sky130_fd_sc_hd__nor2_1 _17156_ (.A(net1878),
    .B(_03484_),
    .Y(_01645_));
 sky130_fd_sc_hd__nand2_1 _17157_ (.A(net555),
    .B(_03318_),
    .Y(_03485_));
 sky130_fd_sc_hd__o2bb2a_1 _17158_ (.A1_N(\core.csr.traps.mcause.csrReadData[12] ),
    .A2_N(net535),
    .B1(_03485_),
    .B2(net621),
    .X(_03486_));
 sky130_fd_sc_hd__nor2_1 _17159_ (.A(net1880),
    .B(_03486_),
    .Y(_01646_));
 sky130_fd_sc_hd__nand2_1 _17160_ (.A(net553),
    .B(_03321_),
    .Y(_03487_));
 sky130_fd_sc_hd__o2bb2a_1 _17161_ (.A1_N(\core.csr.traps.mcause.csrReadData[13] ),
    .A2_N(net534),
    .B1(_03487_),
    .B2(net620),
    .X(_03488_));
 sky130_fd_sc_hd__nor2_1 _17162_ (.A(net1875),
    .B(_03488_),
    .Y(_01647_));
 sky130_fd_sc_hd__nand2_1 _17163_ (.A(net554),
    .B(_03324_),
    .Y(_03489_));
 sky130_fd_sc_hd__o2bb2a_1 _17164_ (.A1_N(\core.csr.traps.mcause.csrReadData[14] ),
    .A2_N(net534),
    .B1(_03489_),
    .B2(net620),
    .X(_03490_));
 sky130_fd_sc_hd__nor2_1 _17165_ (.A(net1875),
    .B(_03490_),
    .Y(_01648_));
 sky130_fd_sc_hd__nand2_1 _17166_ (.A(net553),
    .B(_03327_),
    .Y(_03491_));
 sky130_fd_sc_hd__o2bb2a_1 _17167_ (.A1_N(\core.csr.traps.mcause.csrReadData[15] ),
    .A2_N(net534),
    .B1(_03491_),
    .B2(net620),
    .X(_03492_));
 sky130_fd_sc_hd__nor2_1 _17168_ (.A(net1875),
    .B(_03492_),
    .Y(_01649_));
 sky130_fd_sc_hd__nand2_1 _17169_ (.A(net551),
    .B(_03330_),
    .Y(_03493_));
 sky130_fd_sc_hd__o2bb2a_1 _17170_ (.A1_N(\core.csr.traps.mcause.csrReadData[16] ),
    .A2_N(net536),
    .B1(_03493_),
    .B2(net619),
    .X(_03494_));
 sky130_fd_sc_hd__nor2_1 _17171_ (.A(net1873),
    .B(_03494_),
    .Y(_01650_));
 sky130_fd_sc_hd__nand2_1 _17172_ (.A(net554),
    .B(_03333_),
    .Y(_03495_));
 sky130_fd_sc_hd__o2bb2a_1 _17173_ (.A1_N(\core.csr.traps.mcause.csrReadData[17] ),
    .A2_N(net534),
    .B1(_03495_),
    .B2(net620),
    .X(_03496_));
 sky130_fd_sc_hd__nor2_1 _17174_ (.A(net1875),
    .B(_03496_),
    .Y(_01651_));
 sky130_fd_sc_hd__nand2_1 _17175_ (.A(net551),
    .B(_03336_),
    .Y(_03497_));
 sky130_fd_sc_hd__o2bb2a_1 _17176_ (.A1_N(\core.csr.traps.mcause.csrReadData[18] ),
    .A2_N(net536),
    .B1(_03497_),
    .B2(net619),
    .X(_03498_));
 sky130_fd_sc_hd__nor2_1 _17177_ (.A(net1873),
    .B(_03498_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _17178_ (.A(net549),
    .B(_03339_),
    .Y(_03499_));
 sky130_fd_sc_hd__o2bb2a_1 _17179_ (.A1_N(\core.csr.traps.mcause.csrReadData[19] ),
    .A2_N(net533),
    .B1(_03499_),
    .B2(net619),
    .X(_03500_));
 sky130_fd_sc_hd__nor2_1 _17180_ (.A(net1871),
    .B(_03500_),
    .Y(_01653_));
 sky130_fd_sc_hd__nand2_1 _17181_ (.A(net549),
    .B(_03342_),
    .Y(_03501_));
 sky130_fd_sc_hd__o2bb2a_1 _17182_ (.A1_N(\core.csr.traps.mcause.csrReadData[20] ),
    .A2_N(net533),
    .B1(_03501_),
    .B2(net618),
    .X(_03502_));
 sky130_fd_sc_hd__nor2_1 _17183_ (.A(net1871),
    .B(_03502_),
    .Y(_01654_));
 sky130_fd_sc_hd__nand2_1 _17184_ (.A(net552),
    .B(_03345_),
    .Y(_03503_));
 sky130_fd_sc_hd__o2bb2a_1 _17185_ (.A1_N(\core.csr.traps.mcause.csrReadData[21] ),
    .A2_N(net536),
    .B1(_03503_),
    .B2(net619),
    .X(_03504_));
 sky130_fd_sc_hd__nor2_1 _17186_ (.A(net1873),
    .B(_03504_),
    .Y(_01655_));
 sky130_fd_sc_hd__nand2_2 _17187_ (.A(net552),
    .B(_03348_),
    .Y(_03505_));
 sky130_fd_sc_hd__o2bb2a_1 _17188_ (.A1_N(\core.csr.traps.mcause.csrReadData[22] ),
    .A2_N(net533),
    .B1(_03505_),
    .B2(net618),
    .X(_03506_));
 sky130_fd_sc_hd__nor2_1 _17189_ (.A(net1873),
    .B(_03506_),
    .Y(_01656_));
 sky130_fd_sc_hd__nand2_2 _17190_ (.A(net552),
    .B(_03351_),
    .Y(_03507_));
 sky130_fd_sc_hd__o2bb2a_1 _17191_ (.A1_N(\core.csr.traps.mcause.csrReadData[23] ),
    .A2_N(net533),
    .B1(_03507_),
    .B2(net618),
    .X(_03508_));
 sky130_fd_sc_hd__nor2_1 _17192_ (.A(net1872),
    .B(_03508_),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_2 _17193_ (.A(net551),
    .B(_03354_),
    .Y(_03509_));
 sky130_fd_sc_hd__o2bb2a_1 _17194_ (.A1_N(\core.csr.traps.mcause.csrReadData[24] ),
    .A2_N(net533),
    .B1(_03509_),
    .B2(net618),
    .X(_03510_));
 sky130_fd_sc_hd__nor2_1 _17195_ (.A(net1872),
    .B(_03510_),
    .Y(_01658_));
 sky130_fd_sc_hd__nand2_1 _17196_ (.A(net550),
    .B(_03357_),
    .Y(_03511_));
 sky130_fd_sc_hd__o2bb2a_1 _17197_ (.A1_N(\core.csr.traps.mcause.csrReadData[25] ),
    .A2_N(net533),
    .B1(_03511_),
    .B2(net618),
    .X(_03512_));
 sky130_fd_sc_hd__nor2_1 _17198_ (.A(net1872),
    .B(_03512_),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_1 _17199_ (.A(net550),
    .B(_03360_),
    .Y(_03513_));
 sky130_fd_sc_hd__o2bb2a_1 _17200_ (.A1_N(\core.csr.traps.mcause.csrReadData[26] ),
    .A2_N(net533),
    .B1(_03513_),
    .B2(net618),
    .X(_03514_));
 sky130_fd_sc_hd__nor2_1 _17201_ (.A(net1871),
    .B(_03514_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_2 _17202_ (.A(net552),
    .B(_03363_),
    .Y(_03515_));
 sky130_fd_sc_hd__o2bb2a_1 _17203_ (.A1_N(\core.csr.traps.mcause.csrReadData[27] ),
    .A2_N(net533),
    .B1(_03515_),
    .B2(net618),
    .X(_03516_));
 sky130_fd_sc_hd__nor2_1 _17204_ (.A(net1871),
    .B(_03516_),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_1 _17205_ (.A(net549),
    .B(_03366_),
    .Y(_03517_));
 sky130_fd_sc_hd__o2bb2a_1 _17206_ (.A1_N(\core.csr.traps.mcause.csrReadData[28] ),
    .A2_N(net533),
    .B1(_03517_),
    .B2(net618),
    .X(_03518_));
 sky130_fd_sc_hd__nor2_1 _17207_ (.A(net1871),
    .B(_03518_),
    .Y(_01662_));
 sky130_fd_sc_hd__nand2_2 _17208_ (.A(net549),
    .B(_03369_),
    .Y(_03519_));
 sky130_fd_sc_hd__o2bb2a_1 _17209_ (.A1_N(\core.csr.traps.mcause.csrReadData[29] ),
    .A2_N(net533),
    .B1(_03519_),
    .B2(net618),
    .X(_03520_));
 sky130_fd_sc_hd__nor2_1 _17210_ (.A(net1871),
    .B(_03520_),
    .Y(_01663_));
 sky130_fd_sc_hd__nand2_1 _17211_ (.A(net554),
    .B(_03372_),
    .Y(_03521_));
 sky130_fd_sc_hd__o2bb2a_1 _17212_ (.A1_N(\core.csr.traps.mcause.csrReadData[30] ),
    .A2_N(net534),
    .B1(_03521_),
    .B2(net620),
    .X(_03522_));
 sky130_fd_sc_hd__nor2_1 _17213_ (.A(net1875),
    .B(_03522_),
    .Y(_01664_));
 sky130_fd_sc_hd__nand2_1 _17214_ (.A(net551),
    .B(_03375_),
    .Y(_03523_));
 sky130_fd_sc_hd__a31o_1 _17215_ (.A1(net1102),
    .A2(_03460_),
    .A3(_03523_),
    .B1(net1873),
    .X(_03524_));
 sky130_fd_sc_hd__o21ba_1 _17216_ (.A1(\core.csr.traps.mcause.csrReadData[31] ),
    .A2(_03460_),
    .B1_N(_03524_),
    .X(_01665_));
 sky130_fd_sc_hd__or2_4 _17217_ (.A(_03264_),
    .B(_03382_),
    .X(_03525_));
 sky130_fd_sc_hd__inv_2 _17218_ (.A(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__nor2_2 _17219_ (.A(net544),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _17220_ (.A(\core.csr.trapReturnVector[0] ),
    .B(net518),
    .Y(_03528_));
 sky130_fd_sc_hd__o2bb2a_1 _17221_ (.A1_N(net450),
    .A2_N(net547),
    .B1(_03457_),
    .B2(net518),
    .X(_03529_));
 sky130_fd_sc_hd__a21oi_1 _17222_ (.A1(_03528_),
    .A2(_03529_),
    .B1(net1879),
    .Y(_01666_));
 sky130_fd_sc_hd__nand2_1 _17223_ (.A(\core.csr.trapReturnVector[1] ),
    .B(net519),
    .Y(_03530_));
 sky130_fd_sc_hd__o2bb2a_1 _17224_ (.A1_N(net461),
    .A2_N(net546),
    .B1(_03462_),
    .B2(net519),
    .X(_03531_));
 sky130_fd_sc_hd__a21oi_1 _17225_ (.A1(_03530_),
    .A2(_03531_),
    .B1(net1877),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _17226_ (.A(\core.csr.trapReturnVector[2] ),
    .B(net518),
    .Y(_03532_));
 sky130_fd_sc_hd__o22a_1 _17227_ (.A1(_03827_),
    .A2(net555),
    .B1(_03464_),
    .B2(net518),
    .X(_03533_));
 sky130_fd_sc_hd__a21oi_1 _17228_ (.A1(_03532_),
    .A2(_03533_),
    .B1(net1877),
    .Y(_01668_));
 sky130_fd_sc_hd__a22o_1 _17229_ (.A1(net475),
    .A2(net544),
    .B1(_03466_),
    .B2(_03526_),
    .X(_03534_));
 sky130_fd_sc_hd__a21oi_1 _17230_ (.A1(\core.csr.trapReturnVector[3] ),
    .A2(net520),
    .B1(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__nor2_1 _17231_ (.A(net1875),
    .B(_03535_),
    .Y(_01669_));
 sky130_fd_sc_hd__nand2_1 _17232_ (.A(\core.csr.trapReturnVector[4] ),
    .B(net519),
    .Y(_03536_));
 sky130_fd_sc_hd__o2bb2a_1 _17233_ (.A1_N(net476),
    .A2_N(net546),
    .B1(_03469_),
    .B2(net519),
    .X(_03537_));
 sky130_fd_sc_hd__a21oi_1 _17234_ (.A1(_03536_),
    .A2(_03537_),
    .B1(net1879),
    .Y(_01670_));
 sky130_fd_sc_hd__nand2_1 _17235_ (.A(\core.csr.trapReturnVector[5] ),
    .B(net518),
    .Y(_03538_));
 sky130_fd_sc_hd__o2bb2a_1 _17236_ (.A1_N(net477),
    .A2_N(net546),
    .B1(_03471_),
    .B2(net518),
    .X(_03539_));
 sky130_fd_sc_hd__a21oi_1 _17237_ (.A1(_03538_),
    .A2(_03539_),
    .B1(net1877),
    .Y(_01671_));
 sky130_fd_sc_hd__nand2_1 _17238_ (.A(\core.csr.trapReturnVector[6] ),
    .B(net518),
    .Y(_03540_));
 sky130_fd_sc_hd__o2bb2a_1 _17239_ (.A1_N(net478),
    .A2_N(net546),
    .B1(_03473_),
    .B2(net519),
    .X(_03541_));
 sky130_fd_sc_hd__a21oi_1 _17240_ (.A1(_03540_),
    .A2(_03541_),
    .B1(net1881),
    .Y(_01672_));
 sky130_fd_sc_hd__nand2_1 _17241_ (.A(\core.csr.trapReturnVector[7] ),
    .B(net519),
    .Y(_03542_));
 sky130_fd_sc_hd__o22a_1 _17242_ (.A1(_03826_),
    .A2(net556),
    .B1(_03475_),
    .B2(net519),
    .X(_03543_));
 sky130_fd_sc_hd__a21oi_1 _17243_ (.A1(_03542_),
    .A2(_03543_),
    .B1(net1878),
    .Y(_01673_));
 sky130_fd_sc_hd__nand2_1 _17244_ (.A(\core.csr.trapReturnVector[8] ),
    .B(net520),
    .Y(_03544_));
 sky130_fd_sc_hd__o2bb2a_1 _17245_ (.A1_N(net480),
    .A2_N(net545),
    .B1(_03477_),
    .B2(net520),
    .X(_03545_));
 sky130_fd_sc_hd__a21oi_1 _17246_ (.A1(_03544_),
    .A2(_03545_),
    .B1(net1878),
    .Y(_01674_));
 sky130_fd_sc_hd__nand2_1 _17247_ (.A(\core.csr.trapReturnVector[9] ),
    .B(net517),
    .Y(_03546_));
 sky130_fd_sc_hd__o22a_1 _17248_ (.A1(_03825_),
    .A2(net553),
    .B1(_03479_),
    .B2(net517),
    .X(_03547_));
 sky130_fd_sc_hd__a21oi_1 _17249_ (.A1(_03546_),
    .A2(_03547_),
    .B1(net1876),
    .Y(_01675_));
 sky130_fd_sc_hd__nor2_1 _17250_ (.A(_03481_),
    .B(_03525_),
    .Y(_03548_));
 sky130_fd_sc_hd__a22o_1 _17251_ (.A1(net451),
    .A2(net547),
    .B1(net519),
    .B2(\core.csr.trapReturnVector[10] ),
    .X(_03549_));
 sky130_fd_sc_hd__o21a_1 _17252_ (.A1(_03548_),
    .A2(_03549_),
    .B1(net1831),
    .X(_01676_));
 sky130_fd_sc_hd__a2bb2o_1 _17253_ (.A1_N(_03483_),
    .A2_N(_03525_),
    .B1(net452),
    .B2(net547),
    .X(_03550_));
 sky130_fd_sc_hd__a21oi_1 _17254_ (.A1(\core.csr.trapReturnVector[11] ),
    .A2(net518),
    .B1(_03550_),
    .Y(_03551_));
 sky130_fd_sc_hd__nor2_1 _17255_ (.A(net1878),
    .B(_03551_),
    .Y(_01677_));
 sky130_fd_sc_hd__nand2_1 _17256_ (.A(\core.csr.trapReturnVector[12] ),
    .B(net518),
    .Y(_03552_));
 sky130_fd_sc_hd__o2bb2a_1 _17257_ (.A1_N(net453),
    .A2_N(net547),
    .B1(_03485_),
    .B2(net518),
    .X(_03553_));
 sky130_fd_sc_hd__a21oi_1 _17258_ (.A1(_03552_),
    .A2(_03553_),
    .B1(net1880),
    .Y(_01678_));
 sky130_fd_sc_hd__a2bb2o_1 _17259_ (.A1_N(_03487_),
    .A2_N(_03525_),
    .B1(net454),
    .B2(net545),
    .X(_03554_));
 sky130_fd_sc_hd__a21oi_1 _17260_ (.A1(\core.csr.trapReturnVector[13] ),
    .A2(net517),
    .B1(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__nor2_1 _17261_ (.A(net1876),
    .B(_03555_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand2_1 _17262_ (.A(\core.csr.trapReturnVector[14] ),
    .B(net517),
    .Y(_03556_));
 sky130_fd_sc_hd__o2bb2a_1 _17263_ (.A1_N(net455),
    .A2_N(net545),
    .B1(_03489_),
    .B2(net520),
    .X(_03557_));
 sky130_fd_sc_hd__a21oi_1 _17264_ (.A1(_03556_),
    .A2(_03557_),
    .B1(net1876),
    .Y(_01680_));
 sky130_fd_sc_hd__nand2_1 _17265_ (.A(\core.csr.trapReturnVector[15] ),
    .B(net517),
    .Y(_03558_));
 sky130_fd_sc_hd__o2bb2a_1 _17266_ (.A1_N(net456),
    .A2_N(net545),
    .B1(_03491_),
    .B2(net517),
    .X(_03559_));
 sky130_fd_sc_hd__a21oi_1 _17267_ (.A1(_03558_),
    .A2(_03559_),
    .B1(net1875),
    .Y(_01681_));
 sky130_fd_sc_hd__nand2_1 _17268_ (.A(\core.csr.trapReturnVector[16] ),
    .B(net516),
    .Y(_03560_));
 sky130_fd_sc_hd__o2bb2a_1 _17269_ (.A1_N(net1747),
    .A2_N(net543),
    .B1(_03493_),
    .B2(net516),
    .X(_03561_));
 sky130_fd_sc_hd__a21oi_1 _17270_ (.A1(_03560_),
    .A2(_03561_),
    .B1(net1873),
    .Y(_01682_));
 sky130_fd_sc_hd__nand2_1 _17271_ (.A(\core.csr.trapReturnVector[17] ),
    .B(net517),
    .Y(_03562_));
 sky130_fd_sc_hd__o2bb2a_1 _17272_ (.A1_N(net458),
    .A2_N(net544),
    .B1(_03495_),
    .B2(net517),
    .X(_03563_));
 sky130_fd_sc_hd__a21oi_1 _17273_ (.A1(_03562_),
    .A2(_03563_),
    .B1(net1879),
    .Y(_01683_));
 sky130_fd_sc_hd__nand2_1 _17274_ (.A(\core.csr.trapReturnVector[18] ),
    .B(net516),
    .Y(_03564_));
 sky130_fd_sc_hd__o2bb2a_1 _17275_ (.A1_N(net459),
    .A2_N(net543),
    .B1(_03497_),
    .B2(net516),
    .X(_03565_));
 sky130_fd_sc_hd__a21oi_1 _17276_ (.A1(_03564_),
    .A2(_03565_),
    .B1(net1874),
    .Y(_01684_));
 sky130_fd_sc_hd__nand2_1 _17277_ (.A(\core.csr.trapReturnVector[19] ),
    .B(net515),
    .Y(_03566_));
 sky130_fd_sc_hd__o2bb2a_1 _17278_ (.A1_N(net460),
    .A2_N(net541),
    .B1(_03499_),
    .B2(net515),
    .X(_03567_));
 sky130_fd_sc_hd__a21oi_1 _17279_ (.A1(_03566_),
    .A2(_03567_),
    .B1(net1874),
    .Y(_01685_));
 sky130_fd_sc_hd__nand2_1 _17280_ (.A(\core.csr.trapReturnVector[20] ),
    .B(net515),
    .Y(_03568_));
 sky130_fd_sc_hd__o2bb2a_1 _17281_ (.A1_N(net462),
    .A2_N(net543),
    .B1(_03501_),
    .B2(net515),
    .X(_03569_));
 sky130_fd_sc_hd__a21oi_1 _17282_ (.A1(_03568_),
    .A2(_03569_),
    .B1(net1874),
    .Y(_01686_));
 sky130_fd_sc_hd__a2bb2o_1 _17283_ (.A1_N(_03503_),
    .A2_N(_03525_),
    .B1(net463),
    .B2(net543),
    .X(_03570_));
 sky130_fd_sc_hd__a21oi_1 _17284_ (.A1(\core.csr.trapReturnVector[21] ),
    .A2(net516),
    .B1(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__nor2_1 _17285_ (.A(net1873),
    .B(_03571_),
    .Y(_01687_));
 sky130_fd_sc_hd__nand2_1 _17286_ (.A(\core.csr.trapReturnVector[22] ),
    .B(net515),
    .Y(_03572_));
 sky130_fd_sc_hd__o2bb2a_1 _17287_ (.A1_N(net464),
    .A2_N(net542),
    .B1(_03505_),
    .B2(net516),
    .X(_03573_));
 sky130_fd_sc_hd__a21oi_1 _17288_ (.A1(_03572_),
    .A2(_03573_),
    .B1(net1872),
    .Y(_01688_));
 sky130_fd_sc_hd__nand2_1 _17289_ (.A(\core.csr.trapReturnVector[23] ),
    .B(net515),
    .Y(_03574_));
 sky130_fd_sc_hd__o22a_1 _17290_ (.A1(_03824_),
    .A2(net550),
    .B1(_03507_),
    .B2(net515),
    .X(_03575_));
 sky130_fd_sc_hd__a21oi_1 _17291_ (.A1(_03574_),
    .A2(_03575_),
    .B1(net1872),
    .Y(_01689_));
 sky130_fd_sc_hd__nand2_1 _17292_ (.A(\core.csr.trapReturnVector[24] ),
    .B(net514),
    .Y(_03576_));
 sky130_fd_sc_hd__o2bb2a_1 _17293_ (.A1_N(net466),
    .A2_N(net542),
    .B1(_03509_),
    .B2(net514),
    .X(_03577_));
 sky130_fd_sc_hd__a21oi_1 _17294_ (.A1(_03576_),
    .A2(_03577_),
    .B1(net1872),
    .Y(_01690_));
 sky130_fd_sc_hd__nand2_1 _17295_ (.A(\core.csr.trapReturnVector[25] ),
    .B(net514),
    .Y(_03578_));
 sky130_fd_sc_hd__o2bb2a_1 _17296_ (.A1_N(net467),
    .A2_N(net542),
    .B1(_03511_),
    .B2(net515),
    .X(_03579_));
 sky130_fd_sc_hd__a21oi_1 _17297_ (.A1(_03578_),
    .A2(_03579_),
    .B1(net1872),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_1 _17298_ (.A(\core.csr.trapReturnVector[26] ),
    .B(net514),
    .Y(_03580_));
 sky130_fd_sc_hd__o2bb2a_1 _17299_ (.A1_N(net468),
    .A2_N(net541),
    .B1(_03513_),
    .B2(net514),
    .X(_03581_));
 sky130_fd_sc_hd__a21oi_1 _17300_ (.A1(_03580_),
    .A2(_03581_),
    .B1(net1871),
    .Y(_01692_));
 sky130_fd_sc_hd__nand2_1 _17301_ (.A(\core.csr.trapReturnVector[27] ),
    .B(net514),
    .Y(_03582_));
 sky130_fd_sc_hd__o2bb2a_1 _17302_ (.A1_N(net469),
    .A2_N(net542),
    .B1(_03515_),
    .B2(net515),
    .X(_03583_));
 sky130_fd_sc_hd__a21oi_1 _17303_ (.A1(_03582_),
    .A2(_03583_),
    .B1(net1872),
    .Y(_01693_));
 sky130_fd_sc_hd__nand2_1 _17304_ (.A(\core.csr.trapReturnVector[28] ),
    .B(net514),
    .Y(_03584_));
 sky130_fd_sc_hd__o2bb2a_1 _17305_ (.A1_N(net470),
    .A2_N(net541),
    .B1(_03517_),
    .B2(net514),
    .X(_03585_));
 sky130_fd_sc_hd__a21oi_1 _17306_ (.A1(_03584_),
    .A2(_03585_),
    .B1(net1871),
    .Y(_01694_));
 sky130_fd_sc_hd__nand2_1 _17307_ (.A(\core.csr.trapReturnVector[29] ),
    .B(net514),
    .Y(_03586_));
 sky130_fd_sc_hd__o2bb2a_1 _17308_ (.A1_N(net471),
    .A2_N(net541),
    .B1(_03519_),
    .B2(net514),
    .X(_03587_));
 sky130_fd_sc_hd__a21oi_1 _17309_ (.A1(_03586_),
    .A2(_03587_),
    .B1(net1871),
    .Y(_01695_));
 sky130_fd_sc_hd__nand2_1 _17310_ (.A(\core.csr.trapReturnVector[30] ),
    .B(net517),
    .Y(_03588_));
 sky130_fd_sc_hd__o2bb2a_1 _17311_ (.A1_N(net473),
    .A2_N(net544),
    .B1(_03521_),
    .B2(net517),
    .X(_03589_));
 sky130_fd_sc_hd__a21oi_1 _17312_ (.A1(_03588_),
    .A2(_03589_),
    .B1(net1875),
    .Y(_01696_));
 sky130_fd_sc_hd__nand2_1 _17313_ (.A(\core.csr.trapReturnVector[31] ),
    .B(net516),
    .Y(_03590_));
 sky130_fd_sc_hd__o22a_1 _17314_ (.A1(_03823_),
    .A2(net551),
    .B1(_03523_),
    .B2(net516),
    .X(_03591_));
 sky130_fd_sc_hd__a21oi_1 _17315_ (.A1(_03590_),
    .A2(_03591_),
    .B1(net1874),
    .Y(_01697_));
 sky130_fd_sc_hd__nor2_8 _17316_ (.A(_03277_),
    .B(_03424_),
    .Y(_03592_));
 sky130_fd_sc_hd__mux2_1 _17317_ (.A0(\core.csr.traps.mtvec.csrReadData[0] ),
    .A1(_03281_),
    .S(net640),
    .X(_03593_));
 sky130_fd_sc_hd__and2_1 _17318_ (.A(net1845),
    .B(_03593_),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _17319_ (.A0(\core.csr.traps.mtvec.csrReadData[1] ),
    .A1(_03284_),
    .S(net641),
    .X(_03594_));
 sky130_fd_sc_hd__and2_1 _17320_ (.A(net1844),
    .B(_03594_),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _17321_ (.A0(\core.csr.traps.mtvec.csrReadData[2] ),
    .A1(_03287_),
    .S(net640),
    .X(_03595_));
 sky130_fd_sc_hd__and2_1 _17322_ (.A(net1846),
    .B(_03595_),
    .X(_01700_));
 sky130_fd_sc_hd__nor2_1 _17323_ (.A(\core.csr.traps.mtvec.csrReadData[3] ),
    .B(net640),
    .Y(_03596_));
 sky130_fd_sc_hd__a211oi_1 _17324_ (.A1(_03290_),
    .A2(net640),
    .B1(_03596_),
    .C1(net1881),
    .Y(_01701_));
 sky130_fd_sc_hd__mux2_1 _17325_ (.A0(\core.csr.traps.mtvec.csrReadData[4] ),
    .A1(_03293_),
    .S(net641),
    .X(_03597_));
 sky130_fd_sc_hd__and2_1 _17326_ (.A(net1832),
    .B(_03597_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _17327_ (.A0(\core.csr.traps.mtvec.csrReadData[5] ),
    .A1(_03296_),
    .S(net641),
    .X(_03598_));
 sky130_fd_sc_hd__and2_1 _17328_ (.A(net1844),
    .B(_03598_),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _17329_ (.A0(_03810_),
    .A1(_03300_),
    .S(net640),
    .X(_03599_));
 sky130_fd_sc_hd__nor2_1 _17330_ (.A(net1881),
    .B(_03599_),
    .Y(_01704_));
 sky130_fd_sc_hd__mux2_1 _17331_ (.A0(\core.csr.traps.mtvec.csrReadData[7] ),
    .A1(_03303_),
    .S(net640),
    .X(_03600_));
 sky130_fd_sc_hd__and2_1 _17332_ (.A(net1849),
    .B(_03600_),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_1 _17333_ (.A0(\core.csr.traps.mtvec.csrReadData[8] ),
    .A1(_03306_),
    .S(net641),
    .X(_03601_));
 sky130_fd_sc_hd__and2_1 _17334_ (.A(net1849),
    .B(_03601_),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_1 _17335_ (.A0(\core.csr.traps.mtvec.csrReadData[9] ),
    .A1(_03309_),
    .S(net639),
    .X(_03602_));
 sky130_fd_sc_hd__and2_1 _17336_ (.A(net1833),
    .B(_03602_),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_1 _17337_ (.A0(\core.csr.traps.mtvec.csrReadData[10] ),
    .A1(_03312_),
    .S(_03592_),
    .X(_03603_));
 sky130_fd_sc_hd__and2_1 _17338_ (.A(net1831),
    .B(_03603_),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _17339_ (.A0(\core.csr.traps.mtvec.csrReadData[11] ),
    .A1(_03315_),
    .S(net640),
    .X(_03604_));
 sky130_fd_sc_hd__and2_1 _17340_ (.A(net1847),
    .B(_03604_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _17341_ (.A0(\core.csr.traps.mtvec.csrReadData[12] ),
    .A1(_03318_),
    .S(net640),
    .X(_03605_));
 sky130_fd_sc_hd__and2_1 _17342_ (.A(net1849),
    .B(_03605_),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _17343_ (.A0(\core.csr.traps.mtvec.csrReadData[13] ),
    .A1(_03321_),
    .S(net640),
    .X(_03606_));
 sky130_fd_sc_hd__and2_1 _17344_ (.A(net1847),
    .B(_03606_),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_1 _17345_ (.A0(\core.csr.traps.mtvec.csrReadData[14] ),
    .A1(_03324_),
    .S(net641),
    .X(_03607_));
 sky130_fd_sc_hd__and2_1 _17346_ (.A(net1848),
    .B(_03607_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _17347_ (.A0(\core.csr.traps.mtvec.csrReadData[15] ),
    .A1(_03327_),
    .S(net639),
    .X(_03608_));
 sky130_fd_sc_hd__and2_1 _17348_ (.A(net1828),
    .B(_03608_),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _17349_ (.A0(\core.csr.traps.mtvec.csrReadData[16] ),
    .A1(_03330_),
    .S(net639),
    .X(_03609_));
 sky130_fd_sc_hd__and2_1 _17350_ (.A(net1826),
    .B(_03609_),
    .X(_01714_));
 sky130_fd_sc_hd__mux2_1 _17351_ (.A0(\core.csr.traps.mtvec.csrReadData[17] ),
    .A1(_03333_),
    .S(net639),
    .X(_03610_));
 sky130_fd_sc_hd__and2_1 _17352_ (.A(net1825),
    .B(_03610_),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _17353_ (.A0(\core.csr.traps.mtvec.csrReadData[18] ),
    .A1(_03336_),
    .S(net639),
    .X(_03611_));
 sky130_fd_sc_hd__and2_1 _17354_ (.A(net1815),
    .B(_03611_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _17355_ (.A0(\core.csr.traps.mtvec.csrReadData[19] ),
    .A1(_03339_),
    .S(net638),
    .X(_03612_));
 sky130_fd_sc_hd__and2_1 _17356_ (.A(net1814),
    .B(_03612_),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_1 _17357_ (.A0(\core.csr.traps.mtvec.csrReadData[20] ),
    .A1(_03342_),
    .S(net638),
    .X(_03613_));
 sky130_fd_sc_hd__and2_1 _17358_ (.A(net1810),
    .B(_03613_),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_1 _17359_ (.A0(\core.csr.traps.mtvec.csrReadData[21] ),
    .A1(_03345_),
    .S(net639),
    .X(_03614_));
 sky130_fd_sc_hd__and2_1 _17360_ (.A(net1828),
    .B(_03614_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _17361_ (.A0(\core.csr.traps.mtvec.csrReadData[22] ),
    .A1(_03348_),
    .S(net639),
    .X(_03615_));
 sky130_fd_sc_hd__and2_1 _17362_ (.A(net1818),
    .B(_03615_),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _17363_ (.A0(\core.csr.traps.mtvec.csrReadData[23] ),
    .A1(_03351_),
    .S(net638),
    .X(_03616_));
 sky130_fd_sc_hd__and2_1 _17364_ (.A(net1816),
    .B(_03616_),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _17365_ (.A0(\core.csr.traps.mtvec.csrReadData[24] ),
    .A1(_03354_),
    .S(net638),
    .X(_03617_));
 sky130_fd_sc_hd__and2_1 _17366_ (.A(net1819),
    .B(_03617_),
    .X(_01722_));
 sky130_fd_sc_hd__mux2_1 _17367_ (.A0(\core.csr.traps.mtvec.csrReadData[25] ),
    .A1(_03357_),
    .S(net638),
    .X(_03618_));
 sky130_fd_sc_hd__and2_1 _17368_ (.A(net1816),
    .B(_03618_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _17369_ (.A0(\core.csr.traps.mtvec.csrReadData[26] ),
    .A1(_03360_),
    .S(net638),
    .X(_03619_));
 sky130_fd_sc_hd__and2_1 _17370_ (.A(net1813),
    .B(_03619_),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _17371_ (.A0(\core.csr.traps.mtvec.csrReadData[27] ),
    .A1(_03363_),
    .S(net638),
    .X(_03620_));
 sky130_fd_sc_hd__and2_1 _17372_ (.A(net1818),
    .B(_03620_),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _17373_ (.A0(\core.csr.traps.mtvec.csrReadData[28] ),
    .A1(_03366_),
    .S(net638),
    .X(_03621_));
 sky130_fd_sc_hd__and2_1 _17374_ (.A(net1813),
    .B(_03621_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _17375_ (.A0(\core.csr.traps.mtvec.csrReadData[29] ),
    .A1(_03369_),
    .S(net638),
    .X(_03622_));
 sky130_fd_sc_hd__and2_1 _17376_ (.A(net1810),
    .B(_03622_),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _17377_ (.A0(\core.csr.traps.mtvec.csrReadData[30] ),
    .A1(_03372_),
    .S(net640),
    .X(_03623_));
 sky130_fd_sc_hd__and2_1 _17378_ (.A(net1845),
    .B(_03623_),
    .X(_01728_));
 sky130_fd_sc_hd__mux2_1 _17379_ (.A0(\core.csr.traps.mtvec.csrReadData[31] ),
    .A1(_03375_),
    .S(net638),
    .X(_03624_));
 sky130_fd_sc_hd__and2_1 _17380_ (.A(net1820),
    .B(_03624_),
    .X(_01729_));
 sky130_fd_sc_hd__nor3_4 _17381_ (.A(_03377_),
    .B(_03385_),
    .C(_03419_),
    .Y(_03625_));
 sky130_fd_sc_hd__nor2_1 _17382_ (.A(net546),
    .B(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__a22o_1 _17383_ (.A1(net482),
    .A2(_07057_),
    .B1(_03466_),
    .B2(_03625_),
    .X(_03627_));
 sky130_fd_sc_hd__a21o_1 _17384_ (.A1(\core.csr.traps.machineInterruptEnable ),
    .A2(_03626_),
    .B1(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__o311a_1 _17385_ (.A1(\core.csr.traps.machinePreviousInterruptEnable ),
    .A2(_03828_),
    .A3(net1127),
    .B1(_03628_),
    .C1(net1830),
    .X(_01730_));
 sky130_fd_sc_hd__and2_1 _17386_ (.A(\core.csr.traps.machinePreviousInterruptEnable ),
    .B(_03626_),
    .X(_03629_));
 sky130_fd_sc_hd__a2bb2o_1 _17387_ (.A1_N(_03626_),
    .A2_N(_03475_),
    .B1(net546),
    .B2(\core.csr.traps.machineInterruptEnable ),
    .X(_03630_));
 sky130_fd_sc_hd__o221a_1 _17388_ (.A1(_03828_),
    .A2(net1128),
    .B1(_03629_),
    .B2(_03630_),
    .C1(net1830),
    .X(_01731_));
 sky130_fd_sc_hd__a31o_1 _17389_ (.A1(_03262_),
    .A2(_03263_),
    .A3(_03383_),
    .B1(net547),
    .X(_03631_));
 sky130_fd_sc_hd__clkinv_2 _17390_ (.A(net507),
    .Y(_03632_));
 sky130_fd_sc_hd__a22o_1 _17391_ (.A1(net671),
    .A2(net604),
    .B1(net931),
    .B2(\core.csr.currentInstruction[0] ),
    .X(_03633_));
 sky130_fd_sc_hd__a211o_1 _17392_ (.A1(_03814_),
    .A2(_03633_),
    .B1(net1049),
    .C1(\core.fetchProgramCounter[0] ),
    .X(_03634_));
 sky130_fd_sc_hd__o21a_2 _17393_ (.A1(net450),
    .A2(net1100),
    .B1(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__nand2_1 _17394_ (.A(_03457_),
    .B(net511),
    .Y(_03636_));
 sky130_fd_sc_hd__o221a_1 _17395_ (.A1(\core.csr.traps.mtval.csrReadData[0] ),
    .A2(net511),
    .B1(_03635_),
    .B2(_03636_),
    .C1(net1844),
    .X(_01732_));
 sky130_fd_sc_hd__a22o_2 _17396_ (.A1(net635),
    .A2(net605),
    .B1(net932),
    .B2(\core.csr.currentInstruction[1] ),
    .X(_03637_));
 sky130_fd_sc_hd__a211o_1 _17397_ (.A1(_03815_),
    .A2(_03637_),
    .B1(net1049),
    .C1(\core.fetchProgramCounter[1] ),
    .X(_03638_));
 sky130_fd_sc_hd__o21ai_1 _17398_ (.A1(net461),
    .A2(net1101),
    .B1(_03638_),
    .Y(_03639_));
 sky130_fd_sc_hd__a31o_1 _17399_ (.A1(_03462_),
    .A2(net512),
    .A3(_03639_),
    .B1(net1877),
    .X(_03640_));
 sky130_fd_sc_hd__o21ba_1 _17400_ (.A1(\core.csr.traps.mtval.csrReadData[1] ),
    .A2(net512),
    .B1_N(_03640_),
    .X(_01733_));
 sky130_fd_sc_hd__a221o_1 _17401_ (.A1(_06713_),
    .A2(net604),
    .B1(net931),
    .B2(\core.csr.currentInstruction[2] ),
    .C1(net1605),
    .X(_03641_));
 sky130_fd_sc_hd__o21a_1 _17402_ (.A1(\core.fetchProgramCounter[2] ),
    .A2(net1609),
    .B1(net1101),
    .X(_03642_));
 sky130_fd_sc_hd__a22o_1 _17403_ (.A1(net472),
    .A2(net1049),
    .B1(_03641_),
    .B2(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__nand2_1 _17404_ (.A(_03464_),
    .B(net511),
    .Y(_03644_));
 sky130_fd_sc_hd__o221a_1 _17405_ (.A1(\core.csr.traps.mtval.csrReadData[2] ),
    .A2(net511),
    .B1(_03643_),
    .B2(_03644_),
    .C1(net1829),
    .X(_01734_));
 sky130_fd_sc_hd__a221o_1 _17406_ (.A1(_06715_),
    .A2(net604),
    .B1(net931),
    .B2(\core.csr.currentInstruction[3] ),
    .C1(net1605),
    .X(_03645_));
 sky130_fd_sc_hd__o211a_1 _17407_ (.A1(\core.fetchProgramCounter[3] ),
    .A2(net1609),
    .B1(_03645_),
    .C1(net1101),
    .X(_03646_));
 sky130_fd_sc_hd__a2111o_1 _17408_ (.A1(net475),
    .A2(net1049),
    .B1(_03466_),
    .C1(_03632_),
    .D1(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__o211a_1 _17409_ (.A1(\core.csr.traps.mtval.csrReadData[3] ),
    .A2(net512),
    .B1(_03647_),
    .C1(net1825),
    .X(_01735_));
 sky130_fd_sc_hd__a221o_1 _17410_ (.A1(_06716_),
    .A2(net604),
    .B1(net931),
    .B2(\core.csr.currentInstruction[4] ),
    .C1(net1605),
    .X(_03648_));
 sky130_fd_sc_hd__o21a_1 _17411_ (.A1(\core.fetchProgramCounter[4] ),
    .A2(net1609),
    .B1(net1101),
    .X(_03649_));
 sky130_fd_sc_hd__a22o_1 _17412_ (.A1(net476),
    .A2(net1049),
    .B1(_03648_),
    .B2(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__nand2_1 _17413_ (.A(_03469_),
    .B(net511),
    .Y(_03651_));
 sky130_fd_sc_hd__o221a_1 _17414_ (.A1(\core.csr.traps.mtval.csrReadData[4] ),
    .A2(net511),
    .B1(_03650_),
    .B2(_03651_),
    .C1(net1829),
    .X(_01736_));
 sky130_fd_sc_hd__a221o_1 _17415_ (.A1(_06718_),
    .A2(net604),
    .B1(net931),
    .B2(\core.csr.currentInstruction[5] ),
    .C1(net1605),
    .X(_03652_));
 sky130_fd_sc_hd__o21a_1 _17416_ (.A1(\core.fetchProgramCounter[5] ),
    .A2(net1609),
    .B1(net1100),
    .X(_03653_));
 sky130_fd_sc_hd__a22o_1 _17417_ (.A1(net477),
    .A2(net1049),
    .B1(_03652_),
    .B2(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__nand2_1 _17418_ (.A(_03471_),
    .B(net510),
    .Y(_03655_));
 sky130_fd_sc_hd__o221a_1 _17419_ (.A1(\core.csr.traps.mtval.csrReadData[5] ),
    .A2(net510),
    .B1(_03654_),
    .B2(_03655_),
    .C1(net1829),
    .X(_01737_));
 sky130_fd_sc_hd__a221o_1 _17420_ (.A1(_06720_),
    .A2(net605),
    .B1(net932),
    .B2(\core.csr.currentInstruction[6] ),
    .C1(net1605),
    .X(_03656_));
 sky130_fd_sc_hd__o21a_1 _17421_ (.A1(\core.fetchProgramCounter[6] ),
    .A2(net1609),
    .B1(net1101),
    .X(_03657_));
 sky130_fd_sc_hd__a22o_1 _17422_ (.A1(net478),
    .A2(net1049),
    .B1(_03656_),
    .B2(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__nand2_1 _17423_ (.A(_03473_),
    .B(net511),
    .Y(_03659_));
 sky130_fd_sc_hd__o221a_1 _17424_ (.A1(\core.csr.traps.mtval.csrReadData[6] ),
    .A2(net510),
    .B1(_03658_),
    .B2(_03659_),
    .C1(net1844),
    .X(_01738_));
 sky130_fd_sc_hd__a221o_1 _17425_ (.A1(_06722_),
    .A2(net605),
    .B1(net931),
    .B2(\core.csr.currentInstruction[7] ),
    .C1(net1606),
    .X(_03660_));
 sky130_fd_sc_hd__o21a_1 _17426_ (.A1(\core.fetchProgramCounter[7] ),
    .A2(net1609),
    .B1(net1101),
    .X(_03661_));
 sky130_fd_sc_hd__a22o_1 _17427_ (.A1(net479),
    .A2(net1049),
    .B1(_03660_),
    .B2(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__nand2_1 _17428_ (.A(_03475_),
    .B(net512),
    .Y(_03663_));
 sky130_fd_sc_hd__o221a_1 _17429_ (.A1(\core.csr.traps.mtval.csrReadData[7] ),
    .A2(net510),
    .B1(_03662_),
    .B2(_03663_),
    .C1(net1831),
    .X(_01739_));
 sky130_fd_sc_hd__a221o_1 _17430_ (.A1(_06723_),
    .A2(net605),
    .B1(net932),
    .B2(\core.csr.currentInstruction[8] ),
    .C1(net1606),
    .X(_03664_));
 sky130_fd_sc_hd__o21a_1 _17431_ (.A1(\core.fetchProgramCounter[8] ),
    .A2(net1609),
    .B1(net1100),
    .X(_03665_));
 sky130_fd_sc_hd__a22o_1 _17432_ (.A1(net480),
    .A2(net1049),
    .B1(_03664_),
    .B2(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__nand2_1 _17433_ (.A(_03477_),
    .B(net512),
    .Y(_03667_));
 sky130_fd_sc_hd__o221a_1 _17434_ (.A1(\core.csr.traps.mtval.csrReadData[8] ),
    .A2(net512),
    .B1(_03666_),
    .B2(_03667_),
    .C1(net1831),
    .X(_01740_));
 sky130_fd_sc_hd__a221o_1 _17435_ (.A1(_06725_),
    .A2(net606),
    .B1(net930),
    .B2(\core.csr.currentInstruction[9] ),
    .C1(net1605),
    .X(_03668_));
 sky130_fd_sc_hd__o21a_1 _17436_ (.A1(\core.fetchProgramCounter[9] ),
    .A2(net1608),
    .B1(net1100),
    .X(_03669_));
 sky130_fd_sc_hd__a22o_1 _17437_ (.A1(net481),
    .A2(net1049),
    .B1(_03668_),
    .B2(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__nand2_1 _17438_ (.A(_03479_),
    .B(net509),
    .Y(_03671_));
 sky130_fd_sc_hd__o221a_1 _17439_ (.A1(\core.csr.traps.mtval.csrReadData[9] ),
    .A2(net509),
    .B1(_03670_),
    .B2(_03671_),
    .C1(net1827),
    .X(_01741_));
 sky130_fd_sc_hd__a221o_1 _17440_ (.A1(_06726_),
    .A2(net604),
    .B1(net932),
    .B2(\core.csr.currentInstruction[10] ),
    .C1(net1606),
    .X(_03672_));
 sky130_fd_sc_hd__o21a_1 _17441_ (.A1(\core.fetchProgramCounter[10] ),
    .A2(_02239_),
    .B1(net1100),
    .X(_03673_));
 sky130_fd_sc_hd__a22o_1 _17442_ (.A1(net451),
    .A2(net1050),
    .B1(_03672_),
    .B2(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__nand2_1 _17443_ (.A(_03481_),
    .B(net510),
    .Y(_03675_));
 sky130_fd_sc_hd__o221a_1 _17444_ (.A1(\core.csr.traps.mtval.csrReadData[10] ),
    .A2(net510),
    .B1(_03674_),
    .B2(_03675_),
    .C1(net1831),
    .X(_01742_));
 sky130_fd_sc_hd__a221o_1 _17445_ (.A1(_05068_),
    .A2(net605),
    .B1(net932),
    .B2(\core.csr.currentInstruction[11] ),
    .C1(net1606),
    .X(_03676_));
 sky130_fd_sc_hd__o21a_1 _17446_ (.A1(\core.fetchProgramCounter[11] ),
    .A2(_02239_),
    .B1(net1100),
    .X(_03677_));
 sky130_fd_sc_hd__a22o_1 _17447_ (.A1(net452),
    .A2(net1050),
    .B1(_03676_),
    .B2(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__nand2_1 _17448_ (.A(_03483_),
    .B(net510),
    .Y(_03679_));
 sky130_fd_sc_hd__o221a_1 _17449_ (.A1(\core.csr.traps.mtval.csrReadData[11] ),
    .A2(net510),
    .B1(_03678_),
    .B2(_03679_),
    .C1(net1832),
    .X(_01743_));
 sky130_fd_sc_hd__a221o_1 _17450_ (.A1(_06670_),
    .A2(net606),
    .B1(net930),
    .B2(\core.csr.currentInstruction[12] ),
    .C1(net1605),
    .X(_03680_));
 sky130_fd_sc_hd__o21a_1 _17451_ (.A1(\core.fetchProgramCounter[12] ),
    .A2(net1608),
    .B1(net1100),
    .X(_03681_));
 sky130_fd_sc_hd__a22o_2 _17452_ (.A1(net453),
    .A2(net1050),
    .B1(_03680_),
    .B2(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__nand2_1 _17453_ (.A(_03485_),
    .B(net510),
    .Y(_03683_));
 sky130_fd_sc_hd__o221a_1 _17454_ (.A1(\core.csr.traps.mtval.csrReadData[12] ),
    .A2(net510),
    .B1(_03682_),
    .B2(_03683_),
    .C1(net1847),
    .X(_01744_));
 sky130_fd_sc_hd__a221o_1 _17455_ (.A1(_06668_),
    .A2(net604),
    .B1(net931),
    .B2(\core.csr.currentInstruction[13] ),
    .C1(net1605),
    .X(_03684_));
 sky130_fd_sc_hd__o211a_1 _17456_ (.A1(\core.fetchProgramCounter[13] ),
    .A2(net1609),
    .B1(_03684_),
    .C1(net1100),
    .X(_03685_));
 sky130_fd_sc_hd__nand2_1 _17457_ (.A(_03487_),
    .B(net512),
    .Y(_03686_));
 sky130_fd_sc_hd__a211o_1 _17458_ (.A1(net454),
    .A2(net1050),
    .B1(_03685_),
    .C1(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__o211a_1 _17459_ (.A1(\core.csr.traps.mtval.csrReadData[13] ),
    .A2(net512),
    .B1(_03687_),
    .C1(net1831),
    .X(_01745_));
 sky130_fd_sc_hd__a221o_1 _17460_ (.A1(_06667_),
    .A2(net604),
    .B1(net931),
    .B2(net1799),
    .C1(net1605),
    .X(_03688_));
 sky130_fd_sc_hd__o211a_1 _17461_ (.A1(\core.fetchProgramCounter[14] ),
    .A2(net1609),
    .B1(_03688_),
    .C1(net1100),
    .X(_03689_));
 sky130_fd_sc_hd__nand2_1 _17462_ (.A(_03489_),
    .B(net512),
    .Y(_03690_));
 sky130_fd_sc_hd__a211o_1 _17463_ (.A1(net455),
    .A2(net1050),
    .B1(_03689_),
    .C1(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__o211a_1 _17464_ (.A1(\core.csr.traps.mtval.csrReadData[14] ),
    .A2(net512),
    .B1(_03691_),
    .C1(net1825),
    .X(_01746_));
 sky130_fd_sc_hd__a221o_1 _17465_ (.A1(_06666_),
    .A2(net606),
    .B1(net930),
    .B2(\core.csr.currentInstruction[15] ),
    .C1(net1604),
    .X(_03692_));
 sky130_fd_sc_hd__o21a_1 _17466_ (.A1(\core.fetchProgramCounter[15] ),
    .A2(net1608),
    .B1(net1099),
    .X(_03693_));
 sky130_fd_sc_hd__a22o_1 _17467_ (.A1(net456),
    .A2(net1048),
    .B1(_03692_),
    .B2(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__nand2_1 _17468_ (.A(_03491_),
    .B(net509),
    .Y(_03695_));
 sky130_fd_sc_hd__o221a_1 _17469_ (.A1(\core.csr.traps.mtval.csrReadData[15] ),
    .A2(net509),
    .B1(_03694_),
    .B2(_03695_),
    .C1(net1827),
    .X(_01747_));
 sky130_fd_sc_hd__a221o_1 _17470_ (.A1(_06665_),
    .A2(net603),
    .B1(net928),
    .B2(\core.csr.currentInstruction[16] ),
    .C1(net1604),
    .X(_03696_));
 sky130_fd_sc_hd__o21a_1 _17471_ (.A1(\core.fetchProgramCounter[16] ),
    .A2(net1607),
    .B1(net1098),
    .X(_03697_));
 sky130_fd_sc_hd__a22o_1 _17472_ (.A1(net457),
    .A2(net1047),
    .B1(_03696_),
    .B2(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__nand2_1 _17473_ (.A(_03493_),
    .B(net506),
    .Y(_03699_));
 sky130_fd_sc_hd__o221a_1 _17474_ (.A1(\core.csr.traps.mtval.csrReadData[16] ),
    .A2(net509),
    .B1(_03698_),
    .B2(_03699_),
    .C1(net1826),
    .X(_01748_));
 sky130_fd_sc_hd__a221o_1 _17475_ (.A1(_06664_),
    .A2(net606),
    .B1(net930),
    .B2(\core.csr.currentInstruction[17] ),
    .C1(net1604),
    .X(_03700_));
 sky130_fd_sc_hd__o21a_1 _17476_ (.A1(\core.fetchProgramCounter[17] ),
    .A2(net1608),
    .B1(net1099),
    .X(_03701_));
 sky130_fd_sc_hd__a22o_1 _17477_ (.A1(net458),
    .A2(net1047),
    .B1(_03700_),
    .B2(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__nand2_1 _17478_ (.A(_03495_),
    .B(net509),
    .Y(_03703_));
 sky130_fd_sc_hd__o221a_1 _17479_ (.A1(\core.csr.traps.mtval.csrReadData[17] ),
    .A2(net509),
    .B1(_03702_),
    .B2(_03703_),
    .C1(net1826),
    .X(_01749_));
 sky130_fd_sc_hd__a221o_1 _17480_ (.A1(_06663_),
    .A2(net603),
    .B1(net928),
    .B2(\core.csr.currentInstruction[18] ),
    .C1(net1603),
    .X(_03704_));
 sky130_fd_sc_hd__o21a_1 _17481_ (.A1(\core.fetchProgramCounter[18] ),
    .A2(net1607),
    .B1(net1098),
    .X(_03705_));
 sky130_fd_sc_hd__a22o_1 _17482_ (.A1(net459),
    .A2(net1047),
    .B1(_03704_),
    .B2(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__nand2_1 _17483_ (.A(_03497_),
    .B(net507),
    .Y(_03707_));
 sky130_fd_sc_hd__o221a_1 _17484_ (.A1(\core.csr.traps.mtval.csrReadData[18] ),
    .A2(net507),
    .B1(_03706_),
    .B2(_03707_),
    .C1(net1815),
    .X(_01750_));
 sky130_fd_sc_hd__a221o_1 _17485_ (.A1(_06662_),
    .A2(net603),
    .B1(net928),
    .B2(\core.csr.currentInstruction[19] ),
    .C1(net1604),
    .X(_03708_));
 sky130_fd_sc_hd__o21a_1 _17486_ (.A1(\core.fetchProgramCounter[19] ),
    .A2(net1607),
    .B1(net1098),
    .X(_03709_));
 sky130_fd_sc_hd__a22o_1 _17487_ (.A1(net460),
    .A2(net1047),
    .B1(_03708_),
    .B2(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__nand2_1 _17488_ (.A(_03499_),
    .B(net506),
    .Y(_03711_));
 sky130_fd_sc_hd__o221a_1 _17489_ (.A1(\core.csr.traps.mtval.csrReadData[19] ),
    .A2(net506),
    .B1(_03710_),
    .B2(_03711_),
    .C1(net1814),
    .X(_01751_));
 sky130_fd_sc_hd__a221o_1 _17490_ (.A1(_06660_),
    .A2(net603),
    .B1(net928),
    .B2(\core.csr.currentInstruction[20] ),
    .C1(net1603),
    .X(_03712_));
 sky130_fd_sc_hd__o21a_1 _17491_ (.A1(\core.fetchProgramCounter[20] ),
    .A2(net1607),
    .B1(net1098),
    .X(_03713_));
 sky130_fd_sc_hd__a22o_1 _17492_ (.A1(net462),
    .A2(net1047),
    .B1(_03712_),
    .B2(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__nand2_1 _17493_ (.A(_03501_),
    .B(net506),
    .Y(_03715_));
 sky130_fd_sc_hd__o221a_1 _17494_ (.A1(\core.csr.traps.mtval.csrReadData[20] ),
    .A2(net506),
    .B1(_03714_),
    .B2(_03715_),
    .C1(net1814),
    .X(_01752_));
 sky130_fd_sc_hd__a221o_1 _17495_ (.A1(_06659_),
    .A2(net603),
    .B1(net929),
    .B2(\core.csr.currentInstruction[21] ),
    .C1(net1604),
    .X(_03716_));
 sky130_fd_sc_hd__o21a_1 _17496_ (.A1(\core.fetchProgramCounter[21] ),
    .A2(net1607),
    .B1(net1098),
    .X(_03717_));
 sky130_fd_sc_hd__a22o_1 _17497_ (.A1(net463),
    .A2(net1047),
    .B1(_03716_),
    .B2(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__nand2_1 _17498_ (.A(_03503_),
    .B(net509),
    .Y(_03719_));
 sky130_fd_sc_hd__o221a_1 _17499_ (.A1(\core.csr.traps.mtval.csrReadData[21] ),
    .A2(net513),
    .B1(_03718_),
    .B2(_03719_),
    .C1(net1828),
    .X(_01753_));
 sky130_fd_sc_hd__a221o_1 _17500_ (.A1(_06658_),
    .A2(net603),
    .B1(net928),
    .B2(\core.csr.currentInstruction[22] ),
    .C1(net1604),
    .X(_03720_));
 sky130_fd_sc_hd__o21a_1 _17501_ (.A1(\core.fetchProgramCounter[22] ),
    .A2(net1607),
    .B1(net1099),
    .X(_03721_));
 sky130_fd_sc_hd__a22o_1 _17502_ (.A1(net464),
    .A2(net1048),
    .B1(_03720_),
    .B2(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__nand2_1 _17503_ (.A(_03505_),
    .B(net507),
    .Y(_03723_));
 sky130_fd_sc_hd__o221a_1 _17504_ (.A1(\core.csr.traps.mtval.csrReadData[22] ),
    .A2(net507),
    .B1(_03722_),
    .B2(_03723_),
    .C1(net1818),
    .X(_01754_));
 sky130_fd_sc_hd__a221o_1 _17505_ (.A1(_06656_),
    .A2(net603),
    .B1(net928),
    .B2(\core.csr.currentInstruction[23] ),
    .C1(net1603),
    .X(_03724_));
 sky130_fd_sc_hd__o21a_1 _17506_ (.A1(\core.fetchProgramCounter[23] ),
    .A2(net1607),
    .B1(net1098),
    .X(_03725_));
 sky130_fd_sc_hd__a22o_2 _17507_ (.A1(net465),
    .A2(net1047),
    .B1(_03724_),
    .B2(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__nand2_1 _17508_ (.A(_03507_),
    .B(net508),
    .Y(_03727_));
 sky130_fd_sc_hd__o221a_1 _17509_ (.A1(\core.csr.traps.mtval.csrReadData[23] ),
    .A2(net507),
    .B1(_03726_),
    .B2(_03727_),
    .C1(net1816),
    .X(_01755_));
 sky130_fd_sc_hd__a221o_1 _17510_ (.A1(_06631_),
    .A2(net603),
    .B1(net928),
    .B2(\core.csr.currentInstruction[24] ),
    .C1(net1603),
    .X(_03728_));
 sky130_fd_sc_hd__o21a_1 _17511_ (.A1(\core.fetchProgramCounter[24] ),
    .A2(net1608),
    .B1(net1099),
    .X(_03729_));
 sky130_fd_sc_hd__a22o_1 _17512_ (.A1(net466),
    .A2(net1048),
    .B1(_03728_),
    .B2(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__nand2_1 _17513_ (.A(_03509_),
    .B(net507),
    .Y(_03731_));
 sky130_fd_sc_hd__o221a_1 _17514_ (.A1(\core.csr.traps.mtval.csrReadData[24] ),
    .A2(net507),
    .B1(_03730_),
    .B2(_03731_),
    .C1(net1818),
    .X(_01756_));
 sky130_fd_sc_hd__a221o_1 _17515_ (.A1(_06629_),
    .A2(net603),
    .B1(net928),
    .B2(\core.csr.currentInstruction[25] ),
    .C1(net1603),
    .X(_03732_));
 sky130_fd_sc_hd__o211a_1 _17516_ (.A1(\core.fetchProgramCounter[25] ),
    .A2(net1608),
    .B1(_03732_),
    .C1(net1099),
    .X(_03733_));
 sky130_fd_sc_hd__nand2_1 _17517_ (.A(_03511_),
    .B(net508),
    .Y(_03734_));
 sky130_fd_sc_hd__a211o_1 _17518_ (.A1(net467),
    .A2(net1051),
    .B1(_03733_),
    .C1(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__o211a_1 _17519_ (.A1(\core.csr.traps.mtval.csrReadData[25] ),
    .A2(net508),
    .B1(_03735_),
    .C1(net1816),
    .X(_01757_));
 sky130_fd_sc_hd__a221o_1 _17520_ (.A1(_06627_),
    .A2(net603),
    .B1(net929),
    .B2(\core.csr.currentInstruction[26] ),
    .C1(net1604),
    .X(_03736_));
 sky130_fd_sc_hd__o211a_1 _17521_ (.A1(\core.fetchProgramCounter[26] ),
    .A2(net1607),
    .B1(_03736_),
    .C1(net1098),
    .X(_03737_));
 sky130_fd_sc_hd__a22o_1 _17522_ (.A1(net468),
    .A2(net1047),
    .B1(net551),
    .B2(_03360_),
    .X(_03738_));
 sky130_fd_sc_hd__or2_1 _17523_ (.A(\core.csr.traps.mtval.csrReadData[26] ),
    .B(net507),
    .X(_03739_));
 sky130_fd_sc_hd__o311a_1 _17524_ (.A1(_03632_),
    .A2(_03737_),
    .A3(_03738_),
    .B1(_03739_),
    .C1(net1820),
    .X(_01758_));
 sky130_fd_sc_hd__o2bb2a_1 _17525_ (.A1_N(\core.csr.currentInstruction[27] ),
    .A2_N(net928),
    .B1(_02217_),
    .B2(_06626_),
    .X(_03740_));
 sky130_fd_sc_hd__nor2_1 _17526_ (.A(\core.fetchProgramCounter[27] ),
    .B(net1607),
    .Y(_03741_));
 sky130_fd_sc_hd__a211o_1 _17527_ (.A1(net1608),
    .A2(_03740_),
    .B1(_03741_),
    .C1(net1048),
    .X(_03742_));
 sky130_fd_sc_hd__nand2_1 _17528_ (.A(net469),
    .B(net1051),
    .Y(_03743_));
 sky130_fd_sc_hd__a41o_1 _17529_ (.A1(_03515_),
    .A2(net508),
    .A3(_03742_),
    .A4(_03743_),
    .B1(net1873),
    .X(_03744_));
 sky130_fd_sc_hd__o21ba_1 _17530_ (.A1(\core.csr.traps.mtval.csrReadData[27] ),
    .A2(net508),
    .B1_N(_03744_),
    .X(_01759_));
 sky130_fd_sc_hd__nor2_1 _17531_ (.A(_06625_),
    .B(_02217_),
    .Y(_03745_));
 sky130_fd_sc_hd__a211o_1 _17532_ (.A1(\core.csr.currentInstruction[28] ),
    .A2(net928),
    .B1(net1603),
    .C1(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__nand2_1 _17533_ (.A(_03821_),
    .B(net1603),
    .Y(_03747_));
 sky130_fd_sc_hd__a221o_1 _17534_ (.A1(net470),
    .A2(net1047),
    .B1(net551),
    .B2(_03366_),
    .C1(_03632_),
    .X(_03748_));
 sky130_fd_sc_hd__a31o_1 _17535_ (.A1(net1098),
    .A2(_03746_),
    .A3(_03747_),
    .B1(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__o211a_1 _17536_ (.A1(\core.csr.traps.mtval.csrReadData[28] ),
    .A2(net506),
    .B1(_03749_),
    .C1(net1814),
    .X(_01760_));
 sky130_fd_sc_hd__o2bb2a_1 _17537_ (.A1_N(\core.csr.currentInstruction[29] ),
    .A2_N(net929),
    .B1(_02217_),
    .B2(_06623_),
    .X(_03750_));
 sky130_fd_sc_hd__nor2_1 _17538_ (.A(net1603),
    .B(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__a211o_1 _17539_ (.A1(\core.fetchProgramCounter[29] ),
    .A2(net1603),
    .B1(_03751_),
    .C1(net1047),
    .X(_03752_));
 sky130_fd_sc_hd__o211ai_2 _17540_ (.A1(net471),
    .A2(net1098),
    .B1(net543),
    .C1(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__a31o_1 _17541_ (.A1(_03519_),
    .A2(net506),
    .A3(_03753_),
    .B1(net1874),
    .X(_03754_));
 sky130_fd_sc_hd__o21ba_1 _17542_ (.A1(\core.csr.traps.mtval.csrReadData[29] ),
    .A2(net506),
    .B1_N(_03754_),
    .X(_01761_));
 sky130_fd_sc_hd__a2bb2o_1 _17543_ (.A1_N(_06543_),
    .A2_N(_02217_),
    .B1(net929),
    .B2(\core.csr.currentInstruction[30] ),
    .X(_03755_));
 sky130_fd_sc_hd__and2_1 _17544_ (.A(net1607),
    .B(_03755_),
    .X(_03756_));
 sky130_fd_sc_hd__a211o_1 _17545_ (.A1(\core.fetchProgramCounter[30] ),
    .A2(net1604),
    .B1(_03756_),
    .C1(net1048),
    .X(_03757_));
 sky130_fd_sc_hd__o211a_1 _17546_ (.A1(net473),
    .A2(net1100),
    .B1(net544),
    .C1(_03757_),
    .X(_03758_));
 sky130_fd_sc_hd__nand2_1 _17547_ (.A(_03521_),
    .B(net509),
    .Y(_03759_));
 sky130_fd_sc_hd__o221a_1 _17548_ (.A1(\core.csr.traps.mtval.csrReadData[30] ),
    .A2(net509),
    .B1(_03758_),
    .B2(_03759_),
    .C1(net1825),
    .X(_01762_));
 sky130_fd_sc_hd__o2bb2a_1 _17549_ (.A1_N(\core.csr.currentInstruction[31] ),
    .A2_N(net929),
    .B1(_02217_),
    .B2(_06619_),
    .X(_03760_));
 sky130_fd_sc_hd__nor2_1 _17550_ (.A(net1604),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__a211oi_1 _17551_ (.A1(\core.fetchProgramCounter[31] ),
    .A2(net1603),
    .B1(_03761_),
    .C1(net1051),
    .Y(_03762_));
 sky130_fd_sc_hd__a211o_1 _17552_ (.A1(_03823_),
    .A2(net1051),
    .B1(net551),
    .C1(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__a31o_1 _17553_ (.A1(_03523_),
    .A2(net506),
    .A3(_03763_),
    .B1(net1874),
    .X(_03764_));
 sky130_fd_sc_hd__o21ba_1 _17554_ (.A1(\core.csr.traps.mtval.csrReadData[31] ),
    .A2(net506),
    .B1_N(_03764_),
    .X(_01763_));
 sky130_fd_sc_hd__or3_1 _17555_ (.A(_03276_),
    .B(_03377_),
    .C(_03381_),
    .X(_03765_));
 sky130_fd_sc_hd__and2_4 _17556_ (.A(net1102),
    .B(net637),
    .X(_03766_));
 sky130_fd_sc_hd__nand2_1 _17557_ (.A(net1103),
    .B(net636),
    .Y(_03767_));
 sky130_fd_sc_hd__or2_1 _17558_ (.A(\core.csr.traps.mip.csrReadData[0] ),
    .B(net617),
    .X(_03768_));
 sky130_fd_sc_hd__and2_1 _17559_ (.A(net1847),
    .B(net1103),
    .X(_03769_));
 sky130_fd_sc_hd__o211a_1 _17560_ (.A1(_03281_),
    .A2(net637),
    .B1(_03768_),
    .C1(net1054),
    .X(_01764_));
 sky130_fd_sc_hd__or2_1 _17561_ (.A(\core.csr.traps.mip.csrReadData[1] ),
    .B(net616),
    .X(_03770_));
 sky130_fd_sc_hd__o211a_1 _17562_ (.A1(_03284_),
    .A2(net636),
    .B1(net1053),
    .C1(_03770_),
    .X(_01765_));
 sky130_fd_sc_hd__or2_1 _17563_ (.A(_03287_),
    .B(net636),
    .X(_03771_));
 sky130_fd_sc_hd__o211a_1 _17564_ (.A1(\core.csr.traps.mip.csrReadData[2] ),
    .A2(net616),
    .B1(net1053),
    .C1(_03771_),
    .X(_01766_));
 sky130_fd_sc_hd__nand2b_1 _17565_ (.A_N(net637),
    .B(_03290_),
    .Y(_03772_));
 sky130_fd_sc_hd__o211a_1 _17566_ (.A1(\core.csr.traps.mip.csrReadData[3] ),
    .A2(net616),
    .B1(net1053),
    .C1(_03772_),
    .X(_01767_));
 sky130_fd_sc_hd__or2_1 _17567_ (.A(_03293_),
    .B(net636),
    .X(_03773_));
 sky130_fd_sc_hd__o211a_1 _17568_ (.A1(\core.csr.traps.mip.csrReadData[4] ),
    .A2(net616),
    .B1(net1053),
    .C1(_03773_),
    .X(_01768_));
 sky130_fd_sc_hd__or2_1 _17569_ (.A(_03296_),
    .B(net636),
    .X(_03774_));
 sky130_fd_sc_hd__o211a_1 _17570_ (.A1(\core.csr.traps.mip.csrReadData[5] ),
    .A2(net616),
    .B1(net1053),
    .C1(_03774_),
    .X(_01769_));
 sky130_fd_sc_hd__or2_1 _17571_ (.A(_03299_),
    .B(net636),
    .X(_03775_));
 sky130_fd_sc_hd__o211a_1 _17572_ (.A1(\core.csr.traps.mip.csrReadData[6] ),
    .A2(net616),
    .B1(net1053),
    .C1(_03775_),
    .X(_01770_));
 sky130_fd_sc_hd__or2_1 _17573_ (.A(_03303_),
    .B(net636),
    .X(_03776_));
 sky130_fd_sc_hd__o211a_1 _17574_ (.A1(\core.csr.traps.mip.csrReadData[7] ),
    .A2(net617),
    .B1(net1054),
    .C1(_03776_),
    .X(_01771_));
 sky130_fd_sc_hd__or2_1 _17575_ (.A(_03306_),
    .B(net637),
    .X(_03777_));
 sky130_fd_sc_hd__o211a_1 _17576_ (.A1(\core.csr.traps.mip.csrReadData[8] ),
    .A2(net616),
    .B1(net1053),
    .C1(_03777_),
    .X(_01772_));
 sky130_fd_sc_hd__or2_1 _17577_ (.A(_03309_),
    .B(net637),
    .X(_03778_));
 sky130_fd_sc_hd__o211a_1 _17578_ (.A1(\core.csr.traps.mip.csrReadData[9] ),
    .A2(net615),
    .B1(net1054),
    .C1(_03778_),
    .X(_01773_));
 sky130_fd_sc_hd__or2_1 _17579_ (.A(_03312_),
    .B(net636),
    .X(_03779_));
 sky130_fd_sc_hd__o211a_1 _17580_ (.A1(\core.csr.traps.mip.csrReadData[10] ),
    .A2(net616),
    .B1(net1053),
    .C1(_03779_),
    .X(_01774_));
 sky130_fd_sc_hd__or2_1 _17581_ (.A(_03315_),
    .B(net636),
    .X(_03780_));
 sky130_fd_sc_hd__o211a_1 _17582_ (.A1(\core.csr.traps.mip.csrReadData[11] ),
    .A2(net617),
    .B1(net1054),
    .C1(_03780_),
    .X(_01775_));
 sky130_fd_sc_hd__or2_1 _17583_ (.A(_03318_),
    .B(net636),
    .X(_03781_));
 sky130_fd_sc_hd__o211a_1 _17584_ (.A1(\core.csr.traps.mip.csrReadData[12] ),
    .A2(net617),
    .B1(net1054),
    .C1(_03781_),
    .X(_01776_));
 sky130_fd_sc_hd__or2_1 _17585_ (.A(_03321_),
    .B(net637),
    .X(_03782_));
 sky130_fd_sc_hd__o211a_1 _17586_ (.A1(\core.csr.traps.mip.csrReadData[13] ),
    .A2(net616),
    .B1(net1053),
    .C1(_03782_),
    .X(_01777_));
 sky130_fd_sc_hd__or2_1 _17587_ (.A(_03324_),
    .B(net637),
    .X(_03783_));
 sky130_fd_sc_hd__o211a_1 _17588_ (.A1(\core.csr.traps.mip.csrReadData[14] ),
    .A2(net616),
    .B1(net1053),
    .C1(_03783_),
    .X(_01778_));
 sky130_fd_sc_hd__or2_1 _17589_ (.A(_03327_),
    .B(net637),
    .X(_03784_));
 sky130_fd_sc_hd__o211a_1 _17590_ (.A1(\core.csr.traps.mip.csrReadData[15] ),
    .A2(net615),
    .B1(net1052),
    .C1(_03784_),
    .X(_01779_));
 sky130_fd_sc_hd__or4_4 _17591_ (.A(_02229_),
    .B(_02237_),
    .C(_03381_),
    .D(_03420_),
    .X(_03785_));
 sky130_fd_sc_hd__and2_4 _17592_ (.A(\core.csr.traps.machineInterruptEnable ),
    .B(net1818),
    .X(_03786_));
 sky130_fd_sc_hd__a41o_1 _17593_ (.A1(\core.csr.traps.mie.currentValue[16] ),
    .A2(net1731),
    .A3(net171),
    .A4(_03786_),
    .B1(net1052),
    .X(_03787_));
 sky130_fd_sc_hd__o221a_1 _17594_ (.A1(\core.csr.traps.mip.csrReadData[16] ),
    .A2(net615),
    .B1(_03785_),
    .B2(_03330_),
    .C1(_03787_),
    .X(_01780_));
 sky130_fd_sc_hd__a41o_1 _17595_ (.A1(\core.csr.traps.mie.currentValue[17] ),
    .A2(net1731),
    .A3(net178),
    .A4(_03786_),
    .B1(net1052),
    .X(_03788_));
 sky130_fd_sc_hd__o221a_1 _17596_ (.A1(\core.csr.traps.mip.csrReadData[17] ),
    .A2(net615),
    .B1(_03785_),
    .B2(_03333_),
    .C1(_03788_),
    .X(_01781_));
 sky130_fd_sc_hd__a41o_1 _17597_ (.A1(\core.csr.traps.mie.currentValue[18] ),
    .A2(net1731),
    .A3(net179),
    .A4(_03786_),
    .B1(net1052),
    .X(_03789_));
 sky130_fd_sc_hd__o221a_1 _17598_ (.A1(\core.csr.traps.mip.csrReadData[18] ),
    .A2(net615),
    .B1(_03785_),
    .B2(_03336_),
    .C1(_03789_),
    .X(_01782_));
 sky130_fd_sc_hd__a221o_1 _17599_ (.A1(\core.csr.traps.machineInterruptEnable ),
    .A2(_02228_),
    .B1(net1102),
    .B2(_03339_),
    .C1(_03766_),
    .X(_03790_));
 sky130_fd_sc_hd__o211a_1 _17600_ (.A1(\core.csr.traps.mip.csrReadData[19] ),
    .A2(net614),
    .B1(_03790_),
    .C1(net1814),
    .X(_01783_));
 sky130_fd_sc_hd__a21o_1 _17601_ (.A1(_02220_),
    .A2(_03786_),
    .B1(net1052),
    .X(_03791_));
 sky130_fd_sc_hd__o221a_1 _17602_ (.A1(\core.csr.traps.mip.csrReadData[20] ),
    .A2(net614),
    .B1(_03785_),
    .B2(_03342_),
    .C1(_03791_),
    .X(_01784_));
 sky130_fd_sc_hd__a21o_1 _17603_ (.A1(_02222_),
    .A2(_03786_),
    .B1(net1054),
    .X(_03792_));
 sky130_fd_sc_hd__o221a_1 _17604_ (.A1(\core.csr.traps.mip.csrReadData[21] ),
    .A2(net615),
    .B1(_03785_),
    .B2(_03345_),
    .C1(_03792_),
    .X(_01785_));
 sky130_fd_sc_hd__a41o_1 _17605_ (.A1(\core.csr.traps.mie.currentValue[22] ),
    .A2(net1731),
    .A3(net183),
    .A4(_03786_),
    .B1(net1052),
    .X(_03793_));
 sky130_fd_sc_hd__o221a_1 _17606_ (.A1(\core.csr.traps.mip.csrReadData[22] ),
    .A2(net614),
    .B1(_03785_),
    .B2(_03348_),
    .C1(_03793_),
    .X(_01786_));
 sky130_fd_sc_hd__a221o_1 _17607_ (.A1(\core.csr.traps.machineInterruptEnable ),
    .A2(_02221_),
    .B1(net1102),
    .B2(_03351_),
    .C1(_03766_),
    .X(_03794_));
 sky130_fd_sc_hd__o211a_1 _17608_ (.A1(\core.csr.traps.mip.csrReadData[23] ),
    .A2(net614),
    .B1(_03794_),
    .C1(net1816),
    .X(_01787_));
 sky130_fd_sc_hd__a41o_1 _17609_ (.A1(\core.csr.traps.mie.currentValue[24] ),
    .A2(net1733),
    .A3(net185),
    .A4(_03786_),
    .B1(net1052),
    .X(_03795_));
 sky130_fd_sc_hd__o221a_1 _17610_ (.A1(\core.csr.traps.mip.csrReadData[24] ),
    .A2(net615),
    .B1(_03785_),
    .B2(_03354_),
    .C1(_03795_),
    .X(_01788_));
 sky130_fd_sc_hd__a21o_1 _17611_ (.A1(_02226_),
    .A2(_03786_),
    .B1(net1052),
    .X(_03796_));
 sky130_fd_sc_hd__o221a_1 _17612_ (.A1(\core.csr.traps.mip.csrReadData[25] ),
    .A2(net614),
    .B1(_03785_),
    .B2(_03357_),
    .C1(_03796_),
    .X(_01789_));
 sky130_fd_sc_hd__a221o_1 _17613_ (.A1(\core.csr.traps.machineInterruptEnable ),
    .A2(_02227_),
    .B1(net1102),
    .B2(_03360_),
    .C1(_03766_),
    .X(_03797_));
 sky130_fd_sc_hd__o211a_1 _17614_ (.A1(\core.csr.traps.mip.csrReadData[26] ),
    .A2(net614),
    .B1(_03797_),
    .C1(net1818),
    .X(_01790_));
 sky130_fd_sc_hd__a221o_1 _17615_ (.A1(\core.csr.traps.machineInterruptEnable ),
    .A2(_02224_),
    .B1(net1102),
    .B2(_03363_),
    .C1(_03766_),
    .X(_03798_));
 sky130_fd_sc_hd__o211a_1 _17616_ (.A1(\core.csr.traps.mip.csrReadData[27] ),
    .A2(net614),
    .B1(_03798_),
    .C1(net1818),
    .X(_01791_));
 sky130_fd_sc_hd__a221o_1 _17617_ (.A1(\core.csr.traps.machineInterruptEnable ),
    .A2(_02225_),
    .B1(net1102),
    .B2(_03366_),
    .C1(_03766_),
    .X(_03799_));
 sky130_fd_sc_hd__o211a_1 _17618_ (.A1(\core.csr.traps.mip.csrReadData[28] ),
    .A2(net614),
    .B1(_03799_),
    .C1(net1816),
    .X(_01792_));
 sky130_fd_sc_hd__a41o_1 _17619_ (.A1(\core.csr.traps.mie.currentValue[29] ),
    .A2(net1732),
    .A3(net175),
    .A4(_03786_),
    .B1(net1052),
    .X(_03800_));
 sky130_fd_sc_hd__o221a_1 _17620_ (.A1(\core.csr.traps.mip.csrReadData[29] ),
    .A2(net614),
    .B1(_03785_),
    .B2(_03369_),
    .C1(_03800_),
    .X(_01793_));
 sky130_fd_sc_hd__a221o_1 _17621_ (.A1(\core.csr.traps.machineInterruptEnable ),
    .A2(_02223_),
    .B1(net1102),
    .B2(_03372_),
    .C1(_03766_),
    .X(_03801_));
 sky130_fd_sc_hd__o211a_1 _17622_ (.A1(\core.csr.traps.mip.csrReadData[30] ),
    .A2(net615),
    .B1(_03801_),
    .C1(net1825),
    .X(_01794_));
 sky130_fd_sc_hd__a41o_1 _17623_ (.A1(\core.csr.traps.mie.currentValue[31] ),
    .A2(net1732),
    .A3(net177),
    .A4(_03786_),
    .B1(net1052),
    .X(_03802_));
 sky130_fd_sc_hd__o221a_1 _17624_ (.A1(\core.csr.traps.mip.csrReadData[31] ),
    .A2(net614),
    .B1(_03785_),
    .B2(_03375_),
    .C1(_03802_),
    .X(_01795_));
 sky130_fd_sc_hd__nand2_8 _17625_ (.A(_06851_),
    .B(_08676_),
    .Y(_03803_));
 sky130_fd_sc_hd__mux2_1 _17626_ (.A0(net1079),
    .A1(\core.registers[23][0] ),
    .S(net774),
    .X(_01796_));
 sky130_fd_sc_hd__mux2_1 _17627_ (.A0(net1083),
    .A1(\core.registers[23][1] ),
    .S(net776),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _17628_ (.A0(net1085),
    .A1(\core.registers[23][2] ),
    .S(net774),
    .X(_01798_));
 sky130_fd_sc_hd__mux2_1 _17629_ (.A0(net1091),
    .A1(\core.registers[23][3] ),
    .S(net774),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _17630_ (.A0(net1028),
    .A1(\core.registers[23][4] ),
    .S(net776),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_1 _17631_ (.A0(net1033),
    .A1(\core.registers[23][5] ),
    .S(net776),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _17632_ (.A0(net1037),
    .A1(\core.registers[23][6] ),
    .S(net776),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _17633_ (.A0(net1138),
    .A1(\core.registers[23][7] ),
    .S(net776),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _17634_ (.A0(net899),
    .A1(\core.registers[23][8] ),
    .S(net775),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _17635_ (.A0(net901),
    .A1(\core.registers[23][9] ),
    .S(net776),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _17636_ (.A0(net759),
    .A1(\core.registers[23][10] ),
    .S(net775),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _17637_ (.A0(net761),
    .A1(\core.registers[23][11] ),
    .S(net775),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_1 _17638_ (.A0(net729),
    .A1(\core.registers[23][12] ),
    .S(net775),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _17639_ (.A0(net733),
    .A1(\core.registers[23][13] ),
    .S(net775),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _17640_ (.A0(net737),
    .A1(\core.registers[23][14] ),
    .S(net773),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _17641_ (.A0(net743),
    .A1(\core.registers[23][15] ),
    .S(net773),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _17642_ (.A0(net830),
    .A1(\core.registers[23][16] ),
    .S(net774),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _17643_ (.A0(net835),
    .A1(\core.registers[23][17] ),
    .S(net773),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _17644_ (.A0(net839),
    .A1(\core.registers[23][18] ),
    .S(net775),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _17645_ (.A0(net843),
    .A1(\core.registers[23][19] ),
    .S(net773),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _17646_ (.A0(net848),
    .A1(\core.registers[23][20] ),
    .S(net773),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _17647_ (.A0(net852),
    .A1(\core.registers[23][21] ),
    .S(net773),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _17648_ (.A0(net858),
    .A1(\core.registers[23][22] ),
    .S(net774),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _17649_ (.A0(net862),
    .A1(\core.registers[23][23] ),
    .S(net773),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _17650_ (.A0(net994),
    .A1(\core.registers[23][24] ),
    .S(net773),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _17651_ (.A0(net999),
    .A1(\core.registers[23][25] ),
    .S(net773),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _17652_ (.A0(net1002),
    .A1(\core.registers[23][26] ),
    .S(net775),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _17653_ (.A0(net867),
    .A1(\core.registers[23][27] ),
    .S(net775),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_1 _17654_ (.A0(net869),
    .A1(\core.registers[23][28] ),
    .S(net776),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _17655_ (.A0(net874),
    .A1(\core.registers[23][29] ),
    .S(net775),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _17656_ (.A0(net878),
    .A1(\core.registers[23][30] ),
    .S(net775),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _17657_ (.A0(net1023),
    .A1(\core.registers[23][31] ),
    .S(net773),
    .X(_01827_));
 sky130_fd_sc_hd__nand2_8 _17658_ (.A(_08676_),
    .B(_08761_),
    .Y(_03804_));
 sky130_fd_sc_hd__mux2_1 _17659_ (.A0(net1079),
    .A1(\core.registers[22][0] ),
    .S(net770),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _17660_ (.A0(net1083),
    .A1(\core.registers[22][1] ),
    .S(net772),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _17661_ (.A0(net1086),
    .A1(\core.registers[22][2] ),
    .S(net770),
    .X(_01830_));
 sky130_fd_sc_hd__mux2_1 _17662_ (.A0(net1091),
    .A1(\core.registers[22][3] ),
    .S(net770),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _17663_ (.A0(net1028),
    .A1(\core.registers[22][4] ),
    .S(net772),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _17664_ (.A0(net1033),
    .A1(\core.registers[22][5] ),
    .S(net772),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _17665_ (.A0(net1037),
    .A1(\core.registers[22][6] ),
    .S(net772),
    .X(_01834_));
 sky130_fd_sc_hd__mux2_1 _17666_ (.A0(net1138),
    .A1(\core.registers[22][7] ),
    .S(net772),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _17667_ (.A0(net899),
    .A1(\core.registers[22][8] ),
    .S(net771),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_1 _17668_ (.A0(net901),
    .A1(\core.registers[22][9] ),
    .S(net772),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _17669_ (.A0(net759),
    .A1(\core.registers[22][10] ),
    .S(net771),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_1 _17670_ (.A0(net762),
    .A1(\core.registers[22][11] ),
    .S(net771),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _17671_ (.A0(net729),
    .A1(\core.registers[22][12] ),
    .S(net771),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _17672_ (.A0(net733),
    .A1(\core.registers[22][13] ),
    .S(net771),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _17673_ (.A0(net737),
    .A1(\core.registers[22][14] ),
    .S(net769),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _17674_ (.A0(net742),
    .A1(\core.registers[22][15] ),
    .S(net769),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _17675_ (.A0(net830),
    .A1(\core.registers[22][16] ),
    .S(net770),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _17676_ (.A0(net835),
    .A1(\core.registers[22][17] ),
    .S(net769),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _17677_ (.A0(net838),
    .A1(\core.registers[22][18] ),
    .S(net771),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _17678_ (.A0(net843),
    .A1(\core.registers[22][19] ),
    .S(net769),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _17679_ (.A0(net848),
    .A1(\core.registers[22][20] ),
    .S(net769),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _17680_ (.A0(net852),
    .A1(\core.registers[22][21] ),
    .S(net769),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _17681_ (.A0(net858),
    .A1(\core.registers[22][22] ),
    .S(net770),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _17682_ (.A0(net862),
    .A1(\core.registers[22][23] ),
    .S(net769),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _17683_ (.A0(net994),
    .A1(\core.registers[22][24] ),
    .S(net769),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_1 _17684_ (.A0(net999),
    .A1(\core.registers[22][25] ),
    .S(net769),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _17685_ (.A0(net1002),
    .A1(\core.registers[22][26] ),
    .S(net771),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _17686_ (.A0(net867),
    .A1(\core.registers[22][27] ),
    .S(net771),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _17687_ (.A0(net869),
    .A1(\core.registers[22][28] ),
    .S(net772),
    .X(_01856_));
 sky130_fd_sc_hd__mux2_1 _17688_ (.A0(net874),
    .A1(\core.registers[22][29] ),
    .S(net771),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _17689_ (.A0(net878),
    .A1(\core.registers[22][30] ),
    .S(net771),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _17690_ (.A0(net1023),
    .A1(\core.registers[22][31] ),
    .S(net769),
    .X(_01859_));
 sky130_fd_sc_hd__nand2_2 _17691_ (.A(_08761_),
    .B(_08770_),
    .Y(_03805_));
 sky130_fd_sc_hd__mux2_1 _17692_ (.A0(net1076),
    .A1(\core.registers[14][0] ),
    .S(net768),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _17693_ (.A0(net1080),
    .A1(\core.registers[14][1] ),
    .S(net766),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _17694_ (.A0(net1085),
    .A1(\core.registers[14][2] ),
    .S(net768),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _17695_ (.A0(net1089),
    .A1(\core.registers[14][3] ),
    .S(net765),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _17696_ (.A0(net1027),
    .A1(\core.registers[14][4] ),
    .S(net766),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _17697_ (.A0(net1031),
    .A1(\core.registers[14][5] ),
    .S(net766),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _17698_ (.A0(net1038),
    .A1(\core.registers[14][6] ),
    .S(net766),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _17699_ (.A0(net1137),
    .A1(\core.registers[14][7] ),
    .S(net766),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _17700_ (.A0(net896),
    .A1(\core.registers[14][8] ),
    .S(net767),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _17701_ (.A0(net900),
    .A1(\core.registers[14][9] ),
    .S(net766),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _17702_ (.A0(net758),
    .A1(\core.registers[14][10] ),
    .S(net767),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _17703_ (.A0(net761),
    .A1(\core.registers[14][11] ),
    .S(net767),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _17704_ (.A0(net728),
    .A1(\core.registers[14][12] ),
    .S(net767),
    .X(_01872_));
 sky130_fd_sc_hd__mux2_1 _17705_ (.A0(net732),
    .A1(\core.registers[14][13] ),
    .S(net767),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _17706_ (.A0(net737),
    .A1(\core.registers[14][14] ),
    .S(net765),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _17707_ (.A0(net740),
    .A1(\core.registers[14][15] ),
    .S(net765),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _17708_ (.A0(net830),
    .A1(\core.registers[14][16] ),
    .S(net766),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _17709_ (.A0(net834),
    .A1(\core.registers[14][17] ),
    .S(net768),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _17710_ (.A0(net840),
    .A1(\core.registers[14][18] ),
    .S(net766),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _17711_ (.A0(net844),
    .A1(\core.registers[14][19] ),
    .S(net765),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _17712_ (.A0(net846),
    .A1(\core.registers[14][20] ),
    .S(net765),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _17713_ (.A0(net850),
    .A1(\core.registers[14][21] ),
    .S(net765),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _17714_ (.A0(net855),
    .A1(\core.registers[14][22] ),
    .S(net766),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _17715_ (.A0(net860),
    .A1(\core.registers[14][23] ),
    .S(net765),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _17716_ (.A0(net992),
    .A1(\core.registers[14][24] ),
    .S(net765),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _17717_ (.A0(net996),
    .A1(\core.registers[14][25] ),
    .S(net765),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _17718_ (.A0(net1000),
    .A1(\core.registers[14][26] ),
    .S(net765),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _17719_ (.A0(net865),
    .A1(\core.registers[14][27] ),
    .S(net766),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _17720_ (.A0(net869),
    .A1(\core.registers[14][28] ),
    .S(net767),
    .X(_01888_));
 sky130_fd_sc_hd__mux2_1 _17721_ (.A0(net876),
    .A1(\core.registers[14][29] ),
    .S(net767),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _17722_ (.A0(net878),
    .A1(\core.registers[14][30] ),
    .S(net767),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_1 _17723_ (.A0(net1025),
    .A1(\core.registers[14][31] ),
    .S(net768),
    .X(_01891_));
 sky130_fd_sc_hd__nor2_1 _17724_ (.A(_03807_),
    .B(net602),
    .Y(_03806_));
 sky130_fd_sc_hd__a211o_1 _17725_ (.A1(net1797),
    .A2(net602),
    .B1(_03806_),
    .C1(net1886),
    .X(_01892_));
 sky130_fd_sc_hd__clkbuf_2 _17726_ (.A(\core.registers[0][0] ),
    .X(_00868_));
 sky130_fd_sc_hd__clkbuf_2 _17727_ (.A(\core.registers[0][1] ),
    .X(_00869_));
 sky130_fd_sc_hd__clkbuf_2 _17728_ (.A(\core.registers[0][2] ),
    .X(_00870_));
 sky130_fd_sc_hd__clkbuf_2 _17729_ (.A(\core.registers[0][3] ),
    .X(_00871_));
 sky130_fd_sc_hd__clkbuf_2 _17730_ (.A(\core.registers[0][4] ),
    .X(_00872_));
 sky130_fd_sc_hd__clkbuf_2 _17731_ (.A(\core.registers[0][5] ),
    .X(_00873_));
 sky130_fd_sc_hd__clkbuf_2 _17732_ (.A(\core.registers[0][6] ),
    .X(_00874_));
 sky130_fd_sc_hd__clkbuf_2 _17733_ (.A(\core.registers[0][7] ),
    .X(_00875_));
 sky130_fd_sc_hd__clkbuf_2 _17734_ (.A(\core.registers[0][8] ),
    .X(_00876_));
 sky130_fd_sc_hd__clkbuf_2 _17735_ (.A(\core.registers[0][9] ),
    .X(_00877_));
 sky130_fd_sc_hd__clkbuf_2 _17736_ (.A(\core.registers[0][10] ),
    .X(_00878_));
 sky130_fd_sc_hd__clkbuf_2 _17737_ (.A(\core.registers[0][11] ),
    .X(_00879_));
 sky130_fd_sc_hd__clkbuf_2 _17738_ (.A(\core.registers[0][12] ),
    .X(_00880_));
 sky130_fd_sc_hd__clkbuf_2 _17739_ (.A(\core.registers[0][13] ),
    .X(_00881_));
 sky130_fd_sc_hd__clkbuf_2 _17740_ (.A(\core.registers[0][14] ),
    .X(_00882_));
 sky130_fd_sc_hd__clkbuf_2 _17741_ (.A(\core.registers[0][15] ),
    .X(_00883_));
 sky130_fd_sc_hd__clkbuf_2 _17742_ (.A(\core.registers[0][16] ),
    .X(_00884_));
 sky130_fd_sc_hd__clkbuf_2 _17743_ (.A(\core.registers[0][17] ),
    .X(_00885_));
 sky130_fd_sc_hd__clkbuf_2 _17744_ (.A(\core.registers[0][18] ),
    .X(_00886_));
 sky130_fd_sc_hd__clkbuf_2 _17745_ (.A(\core.registers[0][19] ),
    .X(_00887_));
 sky130_fd_sc_hd__clkbuf_2 _17746_ (.A(\core.registers[0][20] ),
    .X(_00888_));
 sky130_fd_sc_hd__clkbuf_2 _17747_ (.A(\core.registers[0][21] ),
    .X(_00889_));
 sky130_fd_sc_hd__clkbuf_2 _17748_ (.A(\core.registers[0][22] ),
    .X(_00890_));
 sky130_fd_sc_hd__clkbuf_2 _17749_ (.A(\core.registers[0][23] ),
    .X(_00891_));
 sky130_fd_sc_hd__clkbuf_2 _17750_ (.A(\core.registers[0][24] ),
    .X(_00892_));
 sky130_fd_sc_hd__clkbuf_2 _17751_ (.A(\core.registers[0][25] ),
    .X(_00893_));
 sky130_fd_sc_hd__clkbuf_2 _17752_ (.A(\core.registers[0][26] ),
    .X(_00894_));
 sky130_fd_sc_hd__clkbuf_2 _17753_ (.A(\core.registers[0][27] ),
    .X(_00895_));
 sky130_fd_sc_hd__clkbuf_2 _17754_ (.A(\core.registers[0][28] ),
    .X(_00896_));
 sky130_fd_sc_hd__clkbuf_2 _17755_ (.A(\core.registers[0][29] ),
    .X(_00897_));
 sky130_fd_sc_hd__clkbuf_2 _17756_ (.A(\core.registers[0][30] ),
    .X(_00898_));
 sky130_fd_sc_hd__clkbuf_2 _17757_ (.A(\core.registers[0][31] ),
    .X(_00899_));
 sky130_fd_sc_hd__dfxtp_1 _17758_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00000_),
    .Q(\core.registers[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17759_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00001_),
    .Q(\core.registers[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17760_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00002_),
    .Q(\core.registers[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17761_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00003_),
    .Q(\core.registers[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17762_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00004_),
    .Q(\core.registers[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17763_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00005_),
    .Q(\core.registers[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17764_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00006_),
    .Q(\core.registers[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17765_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_00007_),
    .Q(\core.registers[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17766_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00008_),
    .Q(\core.registers[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17767_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00009_),
    .Q(\core.registers[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17768_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00010_),
    .Q(\core.registers[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17769_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00011_),
    .Q(\core.registers[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17770_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00012_),
    .Q(\core.registers[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17771_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00013_),
    .Q(\core.registers[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17772_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00014_),
    .Q(\core.registers[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17773_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00015_),
    .Q(\core.registers[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17774_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00016_),
    .Q(\core.registers[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17775_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00017_),
    .Q(\core.registers[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17776_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_00018_),
    .Q(\core.registers[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17777_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00019_),
    .Q(\core.registers[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17778_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_00020_),
    .Q(\core.registers[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17779_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00021_),
    .Q(\core.registers[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17780_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00022_),
    .Q(\core.registers[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17781_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00023_),
    .Q(\core.registers[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17782_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00024_),
    .Q(\core.registers[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17783_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_00025_),
    .Q(\core.registers[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17784_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00026_),
    .Q(\core.registers[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17785_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00027_),
    .Q(\core.registers[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17786_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00028_),
    .Q(\core.registers[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17787_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00029_),
    .Q(\core.registers[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17788_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00030_),
    .Q(\core.registers[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17789_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00031_),
    .Q(\core.registers[19][31] ));
 sky130_fd_sc_hd__dfxtp_4 _17790_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00032_),
    .Q(\core.csr.currentInstruction[0] ));
 sky130_fd_sc_hd__dfxtp_4 _17791_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00033_),
    .Q(\core.csr.currentInstruction[1] ));
 sky130_fd_sc_hd__dfxtp_4 _17792_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00034_),
    .Q(\core.csr.currentInstruction[2] ));
 sky130_fd_sc_hd__dfxtp_4 _17793_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00035_),
    .Q(\core.csr.currentInstruction[3] ));
 sky130_fd_sc_hd__dfxtp_4 _17794_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00036_),
    .Q(\core.csr.currentInstruction[4] ));
 sky130_fd_sc_hd__dfxtp_4 _17795_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00037_),
    .Q(\core.csr.currentInstruction[5] ));
 sky130_fd_sc_hd__dfxtp_4 _17796_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00038_),
    .Q(\core.csr.currentInstruction[6] ));
 sky130_fd_sc_hd__dfxtp_4 _17797_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00039_),
    .Q(\core.csr.currentInstruction[7] ));
 sky130_fd_sc_hd__dfxtp_4 _17798_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00040_),
    .Q(\core.csr.currentInstruction[8] ));
 sky130_fd_sc_hd__dfxtp_4 _17799_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00041_),
    .Q(\core.csr.currentInstruction[9] ));
 sky130_fd_sc_hd__dfxtp_4 _17800_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00042_),
    .Q(\core.csr.currentInstruction[10] ));
 sky130_fd_sc_hd__dfxtp_4 _17801_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00043_),
    .Q(\core.csr.currentInstruction[11] ));
 sky130_fd_sc_hd__dfxtp_4 _17802_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00044_),
    .Q(\core.csr.currentInstruction[12] ));
 sky130_fd_sc_hd__dfxtp_2 _17803_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00045_),
    .Q(\core.csr.currentInstruction[13] ));
 sky130_fd_sc_hd__dfxtp_2 _17804_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00046_),
    .Q(\core.csr.currentInstruction[14] ));
 sky130_fd_sc_hd__dfxtp_2 _17805_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00047_),
    .Q(\core.csr.currentInstruction[15] ));
 sky130_fd_sc_hd__dfxtp_2 _17806_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00048_),
    .Q(\core.csr.currentInstruction[16] ));
 sky130_fd_sc_hd__dfxtp_2 _17807_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00049_),
    .Q(\core.csr.currentInstruction[17] ));
 sky130_fd_sc_hd__dfxtp_4 _17808_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00050_),
    .Q(\core.csr.currentInstruction[18] ));
 sky130_fd_sc_hd__dfxtp_4 _17809_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00051_),
    .Q(\core.csr.currentInstruction[19] ));
 sky130_fd_sc_hd__dfxtp_4 _17810_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00052_),
    .Q(\core.csr.currentInstruction[20] ));
 sky130_fd_sc_hd__dfxtp_4 _17811_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00053_),
    .Q(\core.csr.currentInstruction[21] ));
 sky130_fd_sc_hd__dfxtp_4 _17812_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00054_),
    .Q(\core.csr.currentInstruction[22] ));
 sky130_fd_sc_hd__dfxtp_4 _17813_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00055_),
    .Q(\core.csr.currentInstruction[23] ));
 sky130_fd_sc_hd__dfxtp_4 _17814_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00056_),
    .Q(\core.csr.currentInstruction[24] ));
 sky130_fd_sc_hd__dfxtp_4 _17815_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00057_),
    .Q(\core.csr.currentInstruction[25] ));
 sky130_fd_sc_hd__dfxtp_4 _17816_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00058_),
    .Q(\core.csr.currentInstruction[26] ));
 sky130_fd_sc_hd__dfxtp_4 _17817_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00059_),
    .Q(\core.csr.currentInstruction[27] ));
 sky130_fd_sc_hd__dfxtp_4 _17818_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00060_),
    .Q(\core.csr.currentInstruction[28] ));
 sky130_fd_sc_hd__dfxtp_4 _17819_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00061_),
    .Q(\core.csr.currentInstruction[29] ));
 sky130_fd_sc_hd__dfxtp_4 _17820_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00062_),
    .Q(\core.csr.currentInstruction[30] ));
 sky130_fd_sc_hd__dfxtp_4 _17821_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00063_),
    .Q(\core.csr.currentInstruction[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17822_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00064_),
    .Q(\core.pipe1_operation.currentPipeStall ));
 sky130_fd_sc_hd__dfxtp_2 _17823_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00065_),
    .Q(\core.csr.cycleTimer.currentValue[0] ));
 sky130_fd_sc_hd__dfxtp_2 _17824_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00066_),
    .Q(\core.csr.cycleTimer.currentValue[1] ));
 sky130_fd_sc_hd__dfxtp_1 _17825_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00067_),
    .Q(\core.csr.cycleTimer.currentValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _17826_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00068_),
    .Q(\core.csr.cycleTimer.currentValue[3] ));
 sky130_fd_sc_hd__dfxtp_1 _17827_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00069_),
    .Q(\core.csr.cycleTimer.currentValue[4] ));
 sky130_fd_sc_hd__dfxtp_1 _17828_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00070_),
    .Q(\core.csr.cycleTimer.currentValue[5] ));
 sky130_fd_sc_hd__dfxtp_1 _17829_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00071_),
    .Q(\core.csr.cycleTimer.currentValue[6] ));
 sky130_fd_sc_hd__dfxtp_2 _17830_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00072_),
    .Q(\core.csr.cycleTimer.currentValue[7] ));
 sky130_fd_sc_hd__dfxtp_1 _17831_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00073_),
    .Q(\core.csr.cycleTimer.currentValue[8] ));
 sky130_fd_sc_hd__dfxtp_1 _17832_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00074_),
    .Q(\core.csr.cycleTimer.currentValue[9] ));
 sky130_fd_sc_hd__dfxtp_2 _17833_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00075_),
    .Q(\core.csr.cycleTimer.currentValue[10] ));
 sky130_fd_sc_hd__dfxtp_1 _17834_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00076_),
    .Q(\core.csr.cycleTimer.currentValue[11] ));
 sky130_fd_sc_hd__dfxtp_1 _17835_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00077_),
    .Q(\core.csr.cycleTimer.currentValue[12] ));
 sky130_fd_sc_hd__dfxtp_2 _17836_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00078_),
    .Q(\core.csr.cycleTimer.currentValue[13] ));
 sky130_fd_sc_hd__dfxtp_1 _17837_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00079_),
    .Q(\core.csr.cycleTimer.currentValue[14] ));
 sky130_fd_sc_hd__dfxtp_1 _17838_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00080_),
    .Q(\core.csr.cycleTimer.currentValue[15] ));
 sky130_fd_sc_hd__dfxtp_2 _17839_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00081_),
    .Q(\core.csr.cycleTimer.currentValue[16] ));
 sky130_fd_sc_hd__dfxtp_1 _17840_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00082_),
    .Q(\core.csr.cycleTimer.currentValue[17] ));
 sky130_fd_sc_hd__dfxtp_1 _17841_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_00083_),
    .Q(\core.csr.cycleTimer.currentValue[18] ));
 sky130_fd_sc_hd__dfxtp_2 _17842_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_00084_),
    .Q(\core.csr.cycleTimer.currentValue[19] ));
 sky130_fd_sc_hd__dfxtp_1 _17843_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00085_),
    .Q(\core.csr.cycleTimer.currentValue[20] ));
 sky130_fd_sc_hd__dfxtp_1 _17844_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00086_),
    .Q(\core.csr.cycleTimer.currentValue[21] ));
 sky130_fd_sc_hd__dfxtp_2 _17845_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00087_),
    .Q(\core.csr.cycleTimer.currentValue[22] ));
 sky130_fd_sc_hd__dfxtp_1 _17846_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00088_),
    .Q(\core.csr.cycleTimer.currentValue[23] ));
 sky130_fd_sc_hd__dfxtp_1 _17847_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00089_),
    .Q(\core.csr.cycleTimer.currentValue[24] ));
 sky130_fd_sc_hd__dfxtp_2 _17848_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00090_),
    .Q(\core.csr.cycleTimer.currentValue[25] ));
 sky130_fd_sc_hd__dfxtp_1 _17849_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00091_),
    .Q(\core.csr.cycleTimer.currentValue[26] ));
 sky130_fd_sc_hd__dfxtp_1 _17850_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00092_),
    .Q(\core.csr.cycleTimer.currentValue[27] ));
 sky130_fd_sc_hd__dfxtp_2 _17851_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00093_),
    .Q(\core.csr.cycleTimer.currentValue[28] ));
 sky130_fd_sc_hd__dfxtp_1 _17852_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00094_),
    .Q(\core.csr.cycleTimer.currentValue[29] ));
 sky130_fd_sc_hd__dfxtp_1 _17853_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00095_),
    .Q(\core.csr.cycleTimer.currentValue[30] ));
 sky130_fd_sc_hd__dfxtp_2 _17854_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_00096_),
    .Q(\core.csr.cycleTimer.currentValue[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17855_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_00097_),
    .Q(\core.csr.cycleTimer.currentValue[32] ));
 sky130_fd_sc_hd__dfxtp_1 _17856_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00098_),
    .Q(\core.csr.cycleTimer.currentValue[33] ));
 sky130_fd_sc_hd__dfxtp_2 _17857_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00099_),
    .Q(\core.csr.cycleTimer.currentValue[34] ));
 sky130_fd_sc_hd__dfxtp_1 _17858_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00100_),
    .Q(\core.csr.cycleTimer.currentValue[35] ));
 sky130_fd_sc_hd__dfxtp_1 _17859_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00101_),
    .Q(\core.csr.cycleTimer.currentValue[36] ));
 sky130_fd_sc_hd__dfxtp_2 _17860_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00102_),
    .Q(\core.csr.cycleTimer.currentValue[37] ));
 sky130_fd_sc_hd__dfxtp_1 _17861_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00103_),
    .Q(\core.csr.cycleTimer.currentValue[38] ));
 sky130_fd_sc_hd__dfxtp_1 _17862_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00104_),
    .Q(\core.csr.cycleTimer.currentValue[39] ));
 sky130_fd_sc_hd__dfxtp_2 _17863_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00105_),
    .Q(\core.csr.cycleTimer.currentValue[40] ));
 sky130_fd_sc_hd__dfxtp_1 _17864_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00106_),
    .Q(\core.csr.cycleTimer.currentValue[41] ));
 sky130_fd_sc_hd__dfxtp_1 _17865_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00107_),
    .Q(\core.csr.cycleTimer.currentValue[42] ));
 sky130_fd_sc_hd__dfxtp_2 _17866_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00108_),
    .Q(\core.csr.cycleTimer.currentValue[43] ));
 sky130_fd_sc_hd__dfxtp_1 _17867_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00109_),
    .Q(\core.csr.cycleTimer.currentValue[44] ));
 sky130_fd_sc_hd__dfxtp_1 _17868_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00110_),
    .Q(\core.csr.cycleTimer.currentValue[45] ));
 sky130_fd_sc_hd__dfxtp_2 _17869_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00111_),
    .Q(\core.csr.cycleTimer.currentValue[46] ));
 sky130_fd_sc_hd__dfxtp_1 _17870_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00112_),
    .Q(\core.csr.cycleTimer.currentValue[47] ));
 sky130_fd_sc_hd__dfxtp_1 _17871_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00113_),
    .Q(\core.csr.cycleTimer.currentValue[48] ));
 sky130_fd_sc_hd__dfxtp_2 _17872_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00114_),
    .Q(\core.csr.cycleTimer.currentValue[49] ));
 sky130_fd_sc_hd__dfxtp_1 _17873_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00115_),
    .Q(\core.csr.cycleTimer.currentValue[50] ));
 sky130_fd_sc_hd__dfxtp_1 _17874_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00116_),
    .Q(\core.csr.cycleTimer.currentValue[51] ));
 sky130_fd_sc_hd__dfxtp_2 _17875_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00117_),
    .Q(\core.csr.cycleTimer.currentValue[52] ));
 sky130_fd_sc_hd__dfxtp_1 _17876_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00118_),
    .Q(\core.csr.cycleTimer.currentValue[53] ));
 sky130_fd_sc_hd__dfxtp_1 _17877_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00119_),
    .Q(\core.csr.cycleTimer.currentValue[54] ));
 sky130_fd_sc_hd__dfxtp_2 _17878_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00120_),
    .Q(\core.csr.cycleTimer.currentValue[55] ));
 sky130_fd_sc_hd__dfxtp_1 _17879_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00121_),
    .Q(\core.csr.cycleTimer.currentValue[56] ));
 sky130_fd_sc_hd__dfxtp_1 _17880_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00122_),
    .Q(\core.csr.cycleTimer.currentValue[57] ));
 sky130_fd_sc_hd__dfxtp_2 _17881_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00123_),
    .Q(\core.csr.cycleTimer.currentValue[58] ));
 sky130_fd_sc_hd__dfxtp_1 _17882_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00124_),
    .Q(\core.csr.cycleTimer.currentValue[59] ));
 sky130_fd_sc_hd__dfxtp_1 _17883_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00125_),
    .Q(\core.csr.cycleTimer.currentValue[60] ));
 sky130_fd_sc_hd__dfxtp_1 _17884_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00126_),
    .Q(\core.csr.cycleTimer.currentValue[61] ));
 sky130_fd_sc_hd__dfxtp_1 _17885_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00127_),
    .Q(\core.csr.cycleTimer.currentValue[62] ));
 sky130_fd_sc_hd__dfxtp_1 _17886_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00128_),
    .Q(\core.csr.cycleTimer.currentValue[63] ));
 sky130_fd_sc_hd__dfxtp_4 _17887_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00129_),
    .Q(\core.pipe0_fetch.currentPipeStall ));
 sky130_fd_sc_hd__dfxtp_2 _17888_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00130_),
    .Q(\core.pipe0_currentInstruction[0] ));
 sky130_fd_sc_hd__dfxtp_2 _17889_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00131_),
    .Q(\core.pipe0_currentInstruction[1] ));
 sky130_fd_sc_hd__dfxtp_2 _17890_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00132_),
    .Q(\core.pipe0_currentInstruction[2] ));
 sky130_fd_sc_hd__dfxtp_2 _17891_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00133_),
    .Q(\core.pipe0_currentInstruction[3] ));
 sky130_fd_sc_hd__dfxtp_4 _17892_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00134_),
    .Q(\core.pipe0_currentInstruction[4] ));
 sky130_fd_sc_hd__dfxtp_4 _17893_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00135_),
    .Q(\core.pipe0_currentInstruction[5] ));
 sky130_fd_sc_hd__dfxtp_4 _17894_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00136_),
    .Q(\core.pipe0_currentInstruction[6] ));
 sky130_fd_sc_hd__dfxtp_4 _17895_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00137_),
    .Q(\core.pipe0_currentInstruction[7] ));
 sky130_fd_sc_hd__dfxtp_4 _17896_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00138_),
    .Q(\core.pipe0_currentInstruction[8] ));
 sky130_fd_sc_hd__dfxtp_4 _17897_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00139_),
    .Q(\core.pipe0_currentInstruction[9] ));
 sky130_fd_sc_hd__dfxtp_4 _17898_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00140_),
    .Q(\core.pipe0_currentInstruction[10] ));
 sky130_fd_sc_hd__dfxtp_4 _17899_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00141_),
    .Q(\core.pipe0_currentInstruction[11] ));
 sky130_fd_sc_hd__dfxtp_4 _17900_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00142_),
    .Q(\core.pipe0_currentInstruction[12] ));
 sky130_fd_sc_hd__dfxtp_4 _17901_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00143_),
    .Q(\core.pipe0_currentInstruction[13] ));
 sky130_fd_sc_hd__dfxtp_4 _17902_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00144_),
    .Q(\core.pipe0_currentInstruction[14] ));
 sky130_fd_sc_hd__dfxtp_2 _17903_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00145_),
    .Q(\core.pipe0_currentInstruction[15] ));
 sky130_fd_sc_hd__dfxtp_4 _17904_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00146_),
    .Q(\core.pipe0_currentInstruction[16] ));
 sky130_fd_sc_hd__dfxtp_4 _17905_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00147_),
    .Q(\core.pipe0_currentInstruction[17] ));
 sky130_fd_sc_hd__dfxtp_4 _17906_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00148_),
    .Q(\core.pipe0_currentInstruction[18] ));
 sky130_fd_sc_hd__dfxtp_4 _17907_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00149_),
    .Q(\core.pipe0_currentInstruction[19] ));
 sky130_fd_sc_hd__dfxtp_4 _17908_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00150_),
    .Q(\core.pipe0_currentInstruction[20] ));
 sky130_fd_sc_hd__dfxtp_4 _17909_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00151_),
    .Q(\core.pipe0_currentInstruction[21] ));
 sky130_fd_sc_hd__dfxtp_1 _17910_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00152_),
    .Q(\core.pipe0_currentInstruction[22] ));
 sky130_fd_sc_hd__dfxtp_1 _17911_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00153_),
    .Q(\core.pipe0_currentInstruction[23] ));
 sky130_fd_sc_hd__dfxtp_4 _17912_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00154_),
    .Q(\core.pipe0_currentInstruction[24] ));
 sky130_fd_sc_hd__dfxtp_4 _17913_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00155_),
    .Q(\core.pipe0_currentInstruction[25] ));
 sky130_fd_sc_hd__dfxtp_4 _17914_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00156_),
    .Q(\core.pipe0_currentInstruction[26] ));
 sky130_fd_sc_hd__dfxtp_4 _17915_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00157_),
    .Q(\core.pipe0_currentInstruction[27] ));
 sky130_fd_sc_hd__dfxtp_4 _17916_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00158_),
    .Q(\core.pipe0_currentInstruction[28] ));
 sky130_fd_sc_hd__dfxtp_4 _17917_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00159_),
    .Q(\core.pipe0_currentInstruction[29] ));
 sky130_fd_sc_hd__dfxtp_4 _17918_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00160_),
    .Q(\core.pipe0_currentInstruction[30] ));
 sky130_fd_sc_hd__dfxtp_4 _17919_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00161_),
    .Q(\core.pipe0_currentInstruction[31] ));
 sky130_fd_sc_hd__dfxtp_4 _17920_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00162_),
    .Q(\core.pipe1_resultRegister[0] ));
 sky130_fd_sc_hd__dfxtp_4 _17921_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00163_),
    .Q(\core.pipe1_resultRegister[1] ));
 sky130_fd_sc_hd__dfxtp_4 _17922_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00164_),
    .Q(\core.pipe1_resultRegister[2] ));
 sky130_fd_sc_hd__dfxtp_4 _17923_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00165_),
    .Q(\core.pipe1_resultRegister[3] ));
 sky130_fd_sc_hd__dfxtp_4 _17924_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00166_),
    .Q(\core.pipe1_resultRegister[4] ));
 sky130_fd_sc_hd__dfxtp_4 _17925_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00167_),
    .Q(\core.pipe1_resultRegister[5] ));
 sky130_fd_sc_hd__dfxtp_4 _17926_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00168_),
    .Q(\core.pipe1_resultRegister[6] ));
 sky130_fd_sc_hd__dfxtp_4 _17927_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00169_),
    .Q(\core.pipe1_resultRegister[7] ));
 sky130_fd_sc_hd__dfxtp_4 _17928_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00170_),
    .Q(\core.pipe1_resultRegister[8] ));
 sky130_fd_sc_hd__dfxtp_4 _17929_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_00171_),
    .Q(\core.pipe1_resultRegister[9] ));
 sky130_fd_sc_hd__dfxtp_4 _17930_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00172_),
    .Q(\core.pipe1_resultRegister[10] ));
 sky130_fd_sc_hd__dfxtp_4 _17931_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_00173_),
    .Q(\core.pipe1_resultRegister[11] ));
 sky130_fd_sc_hd__dfxtp_2 _17932_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00174_),
    .Q(\core.pipe1_resultRegister[12] ));
 sky130_fd_sc_hd__dfxtp_2 _17933_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00175_),
    .Q(\core.pipe1_resultRegister[13] ));
 sky130_fd_sc_hd__dfxtp_2 _17934_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00176_),
    .Q(\core.pipe1_resultRegister[14] ));
 sky130_fd_sc_hd__dfxtp_2 _17935_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00177_),
    .Q(\core.pipe1_resultRegister[15] ));
 sky130_fd_sc_hd__dfxtp_2 _17936_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00178_),
    .Q(\core.pipe1_resultRegister[16] ));
 sky130_fd_sc_hd__dfxtp_2 _17937_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00179_),
    .Q(\core.pipe1_resultRegister[17] ));
 sky130_fd_sc_hd__dfxtp_2 _17938_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00180_),
    .Q(\core.pipe1_resultRegister[18] ));
 sky130_fd_sc_hd__dfxtp_2 _17939_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00181_),
    .Q(\core.pipe1_resultRegister[19] ));
 sky130_fd_sc_hd__dfxtp_2 _17940_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00182_),
    .Q(\core.pipe1_resultRegister[20] ));
 sky130_fd_sc_hd__dfxtp_4 _17941_ (.CLK(clknet_leaf_182_wb_clk_i),
    .D(_00183_),
    .Q(\core.pipe1_resultRegister[21] ));
 sky130_fd_sc_hd__dfxtp_1 _17942_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00184_),
    .Q(\core.pipe1_resultRegister[22] ));
 sky130_fd_sc_hd__dfxtp_2 _17943_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00185_),
    .Q(\core.pipe1_resultRegister[23] ));
 sky130_fd_sc_hd__dfxtp_2 _17944_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00186_),
    .Q(\core.pipe1_resultRegister[24] ));
 sky130_fd_sc_hd__dfxtp_2 _17945_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00187_),
    .Q(\core.pipe1_resultRegister[25] ));
 sky130_fd_sc_hd__dfxtp_2 _17946_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00188_),
    .Q(\core.pipe1_resultRegister[26] ));
 sky130_fd_sc_hd__dfxtp_2 _17947_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00189_),
    .Q(\core.pipe1_resultRegister[27] ));
 sky130_fd_sc_hd__dfxtp_1 _17948_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00190_),
    .Q(\core.pipe1_resultRegister[28] ));
 sky130_fd_sc_hd__dfxtp_4 _17949_ (.CLK(clknet_leaf_182_wb_clk_i),
    .D(_00191_),
    .Q(\core.pipe1_resultRegister[29] ));
 sky130_fd_sc_hd__dfxtp_2 _17950_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00192_),
    .Q(\core.pipe1_resultRegister[30] ));
 sky130_fd_sc_hd__dfxtp_4 _17951_ (.CLK(clknet_leaf_182_wb_clk_i),
    .D(_00193_),
    .Q(\core.pipe1_resultRegister[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17952_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00194_),
    .Q(\core.pipe1_csrData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _17953_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00195_),
    .Q(\core.pipe1_csrData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _17954_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00196_),
    .Q(\core.pipe1_csrData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _17955_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00197_),
    .Q(\core.pipe1_csrData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _17956_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00198_),
    .Q(\core.pipe1_csrData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _17957_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00199_),
    .Q(\core.pipe1_csrData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _17958_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00200_),
    .Q(\core.pipe1_csrData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _17959_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00201_),
    .Q(\core.pipe1_csrData[7] ));
 sky130_fd_sc_hd__dfxtp_2 _17960_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00202_),
    .Q(\core.pipe1_csrData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _17961_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00203_),
    .Q(\core.pipe1_csrData[9] ));
 sky130_fd_sc_hd__dfxtp_1 _17962_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00204_),
    .Q(\core.pipe1_csrData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _17963_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00205_),
    .Q(\core.pipe1_csrData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _17964_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00206_),
    .Q(\core.pipe1_csrData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _17965_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00207_),
    .Q(\core.pipe1_csrData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _17966_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00208_),
    .Q(\core.pipe1_csrData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _17967_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00209_),
    .Q(\core.pipe1_csrData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _17968_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00210_),
    .Q(\core.pipe1_csrData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _17969_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00211_),
    .Q(\core.pipe1_csrData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _17970_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00212_),
    .Q(\core.pipe1_csrData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _17971_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00213_),
    .Q(\core.pipe1_csrData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _17972_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00214_),
    .Q(\core.pipe1_csrData[20] ));
 sky130_fd_sc_hd__dfxtp_1 _17973_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00215_),
    .Q(\core.pipe1_csrData[21] ));
 sky130_fd_sc_hd__dfxtp_1 _17974_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00216_),
    .Q(\core.pipe1_csrData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _17975_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00217_),
    .Q(\core.pipe1_csrData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _17976_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00218_),
    .Q(\core.pipe1_csrData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _17977_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00219_),
    .Q(\core.pipe1_csrData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _17978_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00220_),
    .Q(\core.pipe1_csrData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _17979_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00221_),
    .Q(\core.pipe1_csrData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _17980_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00222_),
    .Q(\core.pipe1_csrData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _17981_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00223_),
    .Q(\core.pipe1_csrData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _17982_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00224_),
    .Q(\core.pipe1_csrData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _17983_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00225_),
    .Q(\core.pipe1_csrData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17984_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00226_),
    .Q(\core.registers[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17985_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00227_),
    .Q(\core.registers[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17986_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_00228_),
    .Q(\core.registers[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17987_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00229_),
    .Q(\core.registers[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17988_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00230_),
    .Q(\core.registers[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17989_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00231_),
    .Q(\core.registers[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17990_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00232_),
    .Q(\core.registers[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17991_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00233_),
    .Q(\core.registers[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17992_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_00234_),
    .Q(\core.registers[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17993_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00235_),
    .Q(\core.registers[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17994_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00236_),
    .Q(\core.registers[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17995_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_00237_),
    .Q(\core.registers[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17996_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00238_),
    .Q(\core.registers[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17997_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00239_),
    .Q(\core.registers[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17998_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00240_),
    .Q(\core.registers[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17999_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00241_),
    .Q(\core.registers[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18000_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00242_),
    .Q(\core.registers[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18001_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00243_),
    .Q(\core.registers[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18002_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00244_),
    .Q(\core.registers[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18003_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00245_),
    .Q(\core.registers[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18004_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_00246_),
    .Q(\core.registers[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18005_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00247_),
    .Q(\core.registers[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18006_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00248_),
    .Q(\core.registers[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18007_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00249_),
    .Q(\core.registers[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18008_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00250_),
    .Q(\core.registers[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18009_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00251_),
    .Q(\core.registers[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18010_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00252_),
    .Q(\core.registers[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18011_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00253_),
    .Q(\core.registers[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18012_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_00254_),
    .Q(\core.registers[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18013_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00255_),
    .Q(\core.registers[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18014_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00256_),
    .Q(\core.registers[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18015_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00257_),
    .Q(\core.registers[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18016_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00258_),
    .Q(\core.registers[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18017_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00259_),
    .Q(\core.registers[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18018_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_00260_),
    .Q(\core.registers[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18019_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00261_),
    .Q(\core.registers[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18020_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00262_),
    .Q(\core.registers[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18021_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00263_),
    .Q(\core.registers[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18022_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00264_),
    .Q(\core.registers[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18023_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00265_),
    .Q(\core.registers[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18024_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_00266_),
    .Q(\core.registers[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18025_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00267_),
    .Q(\core.registers[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18026_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00268_),
    .Q(\core.registers[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18027_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_00269_),
    .Q(\core.registers[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18028_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00270_),
    .Q(\core.registers[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18029_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00271_),
    .Q(\core.registers[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18030_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00272_),
    .Q(\core.registers[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18031_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00273_),
    .Q(\core.registers[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18032_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00274_),
    .Q(\core.registers[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18033_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_00275_),
    .Q(\core.registers[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18034_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00276_),
    .Q(\core.registers[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18035_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00277_),
    .Q(\core.registers[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18036_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00278_),
    .Q(\core.registers[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18037_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00279_),
    .Q(\core.registers[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18038_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00280_),
    .Q(\core.registers[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18039_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_00281_),
    .Q(\core.registers[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18040_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00282_),
    .Q(\core.registers[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18041_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_00283_),
    .Q(\core.registers[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18042_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00284_),
    .Q(\core.registers[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18043_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00285_),
    .Q(\core.registers[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18044_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_00286_),
    .Q(\core.registers[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18045_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00287_),
    .Q(\core.registers[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18046_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00288_),
    .Q(\core.registers[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18047_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00289_),
    .Q(\core.registers[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18048_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00290_),
    .Q(\core.registers[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18049_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00291_),
    .Q(\core.registers[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18050_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00292_),
    .Q(\core.registers[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18051_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00293_),
    .Q(\core.registers[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18052_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00294_),
    .Q(\core.registers[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18053_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00295_),
    .Q(\core.registers[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18054_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00296_),
    .Q(\core.registers[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18055_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_00297_),
    .Q(\core.registers[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18056_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00298_),
    .Q(\core.registers[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18057_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00299_),
    .Q(\core.registers[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18058_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00300_),
    .Q(\core.registers[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18059_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00301_),
    .Q(\core.registers[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18060_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00302_),
    .Q(\core.registers[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18061_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00303_),
    .Q(\core.registers[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18062_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00304_),
    .Q(\core.registers[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18063_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00305_),
    .Q(\core.registers[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18064_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00306_),
    .Q(\core.registers[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18065_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00307_),
    .Q(\core.registers[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18066_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00308_),
    .Q(\core.registers[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18067_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00309_),
    .Q(\core.registers[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18068_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_00310_),
    .Q(\core.registers[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18069_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00311_),
    .Q(\core.registers[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18070_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00312_),
    .Q(\core.registers[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18071_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_00313_),
    .Q(\core.registers[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18072_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_00314_),
    .Q(\core.registers[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18073_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00315_),
    .Q(\core.registers[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18074_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00316_),
    .Q(\core.registers[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18075_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00317_),
    .Q(\core.registers[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18076_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00318_),
    .Q(\core.registers[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18077_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00319_),
    .Q(\core.registers[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18078_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00320_),
    .Q(\core.registers[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18079_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00321_),
    .Q(\core.registers[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18080_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00322_),
    .Q(\core.cancelStall ));
 sky130_fd_sc_hd__dfxtp_1 _18081_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00323_),
    .Q(\jtag.managementAddress[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18082_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00324_),
    .Q(\jtag.managementAddress[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18083_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00325_),
    .Q(\jtag.managementAddress[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18084_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00326_),
    .Q(\jtag.managementAddress[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18085_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00327_),
    .Q(\jtag.managementAddress[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18086_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00328_),
    .Q(\jtag.managementAddress[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18087_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00329_),
    .Q(\jtag.managementAddress[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18088_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00330_),
    .Q(\jtag.managementAddress[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18089_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00331_),
    .Q(\jtag.managementAddress[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18090_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00332_),
    .Q(\jtag.managementAddress[9] ));
 sky130_fd_sc_hd__dfxtp_2 _18091_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00333_),
    .Q(\jtag.managementAddress[10] ));
 sky130_fd_sc_hd__dfxtp_2 _18092_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00334_),
    .Q(\jtag.managementAddress[11] ));
 sky130_fd_sc_hd__dfxtp_2 _18093_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00335_),
    .Q(\jtag.managementAddress[12] ));
 sky130_fd_sc_hd__dfxtp_1 _18094_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00336_),
    .Q(\jtag.managementAddress[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18095_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00337_),
    .Q(\jtag.managementAddress[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18096_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00338_),
    .Q(\jtag.managementAddress[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18097_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00339_),
    .Q(\jtag.managementAddress[16] ));
 sky130_fd_sc_hd__dfxtp_1 _18098_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00340_),
    .Q(\jtag.managementAddress[17] ));
 sky130_fd_sc_hd__dfxtp_1 _18099_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00341_),
    .Q(\jtag.managementAddress[18] ));
 sky130_fd_sc_hd__dfxtp_1 _18100_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00342_),
    .Q(\jtag.managementAddress[19] ));
 sky130_fd_sc_hd__dfxtp_4 _18101_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00343_),
    .Q(net450));
 sky130_fd_sc_hd__dfxtp_4 _18102_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00344_),
    .Q(net461));
 sky130_fd_sc_hd__dfxtp_4 _18103_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00345_),
    .Q(net472));
 sky130_fd_sc_hd__dfxtp_4 _18104_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00346_),
    .Q(net475));
 sky130_fd_sc_hd__dfxtp_4 _18105_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00347_),
    .Q(net476));
 sky130_fd_sc_hd__dfxtp_4 _18106_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00348_),
    .Q(net477));
 sky130_fd_sc_hd__dfxtp_4 _18107_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00349_),
    .Q(net478));
 sky130_fd_sc_hd__dfxtp_4 _18108_ (.CLK(clknet_leaf_145_wb_clk_i),
    .D(_00350_),
    .Q(net479));
 sky130_fd_sc_hd__dfxtp_4 _18109_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_00351_),
    .Q(net480));
 sky130_fd_sc_hd__dfxtp_4 _18110_ (.CLK(clknet_leaf_145_wb_clk_i),
    .D(_00352_),
    .Q(net481));
 sky130_fd_sc_hd__dfxtp_4 _18111_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00353_),
    .Q(net451));
 sky130_fd_sc_hd__dfxtp_4 _18112_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00354_),
    .Q(net452));
 sky130_fd_sc_hd__dfxtp_4 _18113_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_00355_),
    .Q(net453));
 sky130_fd_sc_hd__dfxtp_4 _18114_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00356_),
    .Q(net454));
 sky130_fd_sc_hd__dfxtp_4 _18115_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00357_),
    .Q(net455));
 sky130_fd_sc_hd__dfxtp_4 _18116_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00358_),
    .Q(net456));
 sky130_fd_sc_hd__dfxtp_4 _18117_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00359_),
    .Q(net457));
 sky130_fd_sc_hd__dfxtp_4 _18118_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00360_),
    .Q(net458));
 sky130_fd_sc_hd__dfxtp_4 _18119_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00361_),
    .Q(net459));
 sky130_fd_sc_hd__dfxtp_4 _18120_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00362_),
    .Q(net460));
 sky130_fd_sc_hd__dfxtp_4 _18121_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00363_),
    .Q(net462));
 sky130_fd_sc_hd__dfxtp_4 _18122_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00364_),
    .Q(net463));
 sky130_fd_sc_hd__dfxtp_4 _18123_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00365_),
    .Q(net464));
 sky130_fd_sc_hd__dfxtp_4 _18124_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_00366_),
    .Q(net465));
 sky130_fd_sc_hd__dfxtp_4 _18125_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_00367_),
    .Q(net466));
 sky130_fd_sc_hd__dfxtp_4 _18126_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00368_),
    .Q(net467));
 sky130_fd_sc_hd__dfxtp_4 _18127_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00369_),
    .Q(net468));
 sky130_fd_sc_hd__dfxtp_4 _18128_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00370_),
    .Q(net469));
 sky130_fd_sc_hd__dfxtp_4 _18129_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00371_),
    .Q(net470));
 sky130_fd_sc_hd__dfxtp_4 _18130_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00372_),
    .Q(net471));
 sky130_fd_sc_hd__dfxtp_4 _18131_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00373_),
    .Q(net473));
 sky130_fd_sc_hd__dfxtp_4 _18132_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_00374_),
    .Q(net474));
 sky130_fd_sc_hd__dfxtp_1 _18133_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00375_),
    .Q(\core.registers[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18134_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00376_),
    .Q(\core.registers[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18135_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_00377_),
    .Q(\core.registers[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18136_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00378_),
    .Q(\core.registers[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18137_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_00379_),
    .Q(\core.registers[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18138_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00380_),
    .Q(\core.registers[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18139_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00381_),
    .Q(\core.registers[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18140_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00382_),
    .Q(\core.registers[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18141_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00383_),
    .Q(\core.registers[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18142_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00384_),
    .Q(\core.registers[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18143_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00385_),
    .Q(\core.registers[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18144_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00386_),
    .Q(\core.registers[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18145_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00387_),
    .Q(\core.registers[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18146_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00388_),
    .Q(\core.registers[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18147_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00389_),
    .Q(\core.registers[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18148_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00390_),
    .Q(\core.registers[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18149_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00391_),
    .Q(\core.registers[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18150_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_00392_),
    .Q(\core.registers[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18151_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00393_),
    .Q(\core.registers[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18152_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00394_),
    .Q(\core.registers[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18153_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_00395_),
    .Q(\core.registers[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18154_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_00396_),
    .Q(\core.registers[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18155_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00397_),
    .Q(\core.registers[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18156_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_00398_),
    .Q(\core.registers[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18157_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_00399_),
    .Q(\core.registers[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18158_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_00400_),
    .Q(\core.registers[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18159_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_00401_),
    .Q(\core.registers[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18160_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00402_),
    .Q(\core.registers[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18161_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00403_),
    .Q(\core.registers[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18162_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00404_),
    .Q(\core.registers[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18163_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00405_),
    .Q(\core.registers[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18164_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_00406_),
    .Q(\core.registers[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18165_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00407_),
    .Q(\core.registers[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18166_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00408_),
    .Q(\core.registers[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18167_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00409_),
    .Q(\core.registers[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18168_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00410_),
    .Q(\core.registers[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18169_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_00411_),
    .Q(\core.registers[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18170_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00412_),
    .Q(\core.registers[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18171_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00413_),
    .Q(\core.registers[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18172_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00414_),
    .Q(\core.registers[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18173_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00415_),
    .Q(\core.registers[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18174_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00416_),
    .Q(\core.registers[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18175_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00417_),
    .Q(\core.registers[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18176_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_00418_),
    .Q(\core.registers[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18177_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00419_),
    .Q(\core.registers[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18178_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00420_),
    .Q(\core.registers[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18179_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00421_),
    .Q(\core.registers[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18180_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00422_),
    .Q(\core.registers[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18181_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00423_),
    .Q(\core.registers[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18182_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00424_),
    .Q(\core.registers[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18183_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_00425_),
    .Q(\core.registers[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18184_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00426_),
    .Q(\core.registers[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18185_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_00427_),
    .Q(\core.registers[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18186_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_00428_),
    .Q(\core.registers[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18187_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00429_),
    .Q(\core.registers[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18188_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00430_),
    .Q(\core.registers[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18189_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00431_),
    .Q(\core.registers[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18190_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_00432_),
    .Q(\core.registers[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18191_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_00433_),
    .Q(\core.registers[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18192_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00434_),
    .Q(\core.registers[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18193_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00435_),
    .Q(\core.registers[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18194_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00436_),
    .Q(\core.registers[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18195_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00437_),
    .Q(\core.registers[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18196_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_00438_),
    .Q(\core.registers[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18197_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00439_),
    .Q(\localMemoryInterface.lastCoreByteSelect[0] ));
 sky130_fd_sc_hd__dfxtp_2 _18198_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00440_),
    .Q(\localMemoryInterface.lastCoreByteSelect[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18199_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00441_),
    .Q(\localMemoryInterface.lastCoreByteSelect[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18200_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00442_),
    .Q(\localMemoryInterface.lastCoreByteSelect[3] ));
 sky130_fd_sc_hd__dfxtp_2 _18201_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00443_),
    .Q(\memoryController.last_instruction_enableLocalMemory ));
 sky130_fd_sc_hd__dfxtp_2 _18202_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00444_),
    .Q(\memoryController.last_data_enableLocalMemory ));
 sky130_fd_sc_hd__dfxtp_1 _18203_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00445_),
    .Q(\memoryController.last_instruction_enableWB ));
 sky130_fd_sc_hd__dfxtp_1 _18204_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00446_),
    .Q(\core.registers[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18205_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00447_),
    .Q(\core.registers[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18206_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_00448_),
    .Q(\core.registers[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18207_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00449_),
    .Q(\core.registers[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18208_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00450_),
    .Q(\core.registers[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18209_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00451_),
    .Q(\core.registers[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18210_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00452_),
    .Q(\core.registers[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18211_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00453_),
    .Q(\core.registers[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18212_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00454_),
    .Q(\core.registers[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18213_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00455_),
    .Q(\core.registers[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18214_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00456_),
    .Q(\core.registers[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18215_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_00457_),
    .Q(\core.registers[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18216_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00458_),
    .Q(\core.registers[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18217_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00459_),
    .Q(\core.registers[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18218_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00460_),
    .Q(\core.registers[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18219_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00461_),
    .Q(\core.registers[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18220_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00462_),
    .Q(\core.registers[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18221_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00463_),
    .Q(\core.registers[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18222_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_00464_),
    .Q(\core.registers[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18223_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00465_),
    .Q(\core.registers[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18224_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00466_),
    .Q(\core.registers[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18225_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00467_),
    .Q(\core.registers[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18226_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00468_),
    .Q(\core.registers[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18227_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_00469_),
    .Q(\core.registers[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18228_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_00470_),
    .Q(\core.registers[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18229_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00471_),
    .Q(\core.registers[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18230_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00472_),
    .Q(\core.registers[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18231_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00473_),
    .Q(\core.registers[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18232_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00474_),
    .Q(\core.registers[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18233_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00475_),
    .Q(\core.registers[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18234_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00476_),
    .Q(\core.registers[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18235_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00477_),
    .Q(\core.registers[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18236_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00478_),
    .Q(\core.registers[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18237_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00479_),
    .Q(\core.registers[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18238_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_00480_),
    .Q(\core.registers[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18239_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00481_),
    .Q(\core.registers[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18240_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00482_),
    .Q(\core.registers[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18241_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00483_),
    .Q(\core.registers[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18242_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00484_),
    .Q(\core.registers[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18243_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00485_),
    .Q(\core.registers[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18244_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00486_),
    .Q(\core.registers[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18245_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00487_),
    .Q(\core.registers[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18246_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00488_),
    .Q(\core.registers[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18247_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00489_),
    .Q(\core.registers[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18248_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_00490_),
    .Q(\core.registers[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18249_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00491_),
    .Q(\core.registers[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18250_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00492_),
    .Q(\core.registers[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18251_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00493_),
    .Q(\core.registers[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18252_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00494_),
    .Q(\core.registers[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18253_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00495_),
    .Q(\core.registers[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18254_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00496_),
    .Q(\core.registers[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18255_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00497_),
    .Q(\core.registers[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18256_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00498_),
    .Q(\core.registers[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18257_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_00499_),
    .Q(\core.registers[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18258_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00500_),
    .Q(\core.registers[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18259_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_00501_),
    .Q(\core.registers[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18260_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00502_),
    .Q(\core.registers[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18261_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_00503_),
    .Q(\core.registers[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18262_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_00504_),
    .Q(\core.registers[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18263_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00505_),
    .Q(\core.registers[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18264_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00506_),
    .Q(\core.registers[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18265_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00507_),
    .Q(\core.registers[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18266_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00508_),
    .Q(\core.registers[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18267_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_00509_),
    .Q(\core.registers[8][31] ));
 sky130_fd_sc_hd__dfxtp_4 _18268_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_00510_),
    .Q(\localMemoryInterface.coreReadReady ));
 sky130_fd_sc_hd__dfxtp_2 _18269_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00511_),
    .Q(\localMemoryInterface.lastWBByteSelect[0] ));
 sky130_fd_sc_hd__dfxtp_2 _18270_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00512_),
    .Q(\localMemoryInterface.lastWBByteSelect[1] ));
 sky130_fd_sc_hd__dfxtp_2 _18271_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00513_),
    .Q(\localMemoryInterface.lastWBByteSelect[2] ));
 sky130_fd_sc_hd__dfxtp_2 _18272_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00514_),
    .Q(\localMemoryInterface.lastWBByteSelect[3] ));
 sky130_fd_sc_hd__dfxtp_4 _18273_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00515_),
    .Q(\localMemoryInterface.lastRWBankSelect ));
 sky130_fd_sc_hd__dfxtp_1 _18274_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00516_),
    .Q(\localMemoryInterface.wbReadReady ));
 sky130_fd_sc_hd__dfxtp_1 _18275_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00517_),
    .Q(\core.pipe0_fetch.lastProgramCounter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18276_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00518_),
    .Q(\core.pipe0_fetch.lastProgramCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18277_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_00519_),
    .Q(\core.pipe0_fetch.lastProgramCounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18278_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00520_),
    .Q(\core.pipe0_fetch.lastProgramCounter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18279_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_00521_),
    .Q(\core.pipe0_fetch.lastProgramCounter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18280_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00522_),
    .Q(\core.pipe0_fetch.lastProgramCounter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18281_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00523_),
    .Q(\core.pipe0_fetch.lastProgramCounter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18282_ (.CLK(clknet_leaf_145_wb_clk_i),
    .D(_00524_),
    .Q(\core.pipe0_fetch.lastProgramCounter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18283_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_00525_),
    .Q(\core.pipe0_fetch.lastProgramCounter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18284_ (.CLK(clknet_leaf_145_wb_clk_i),
    .D(_00526_),
    .Q(\core.pipe0_fetch.lastProgramCounter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _18285_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00527_),
    .Q(\core.pipe0_fetch.lastProgramCounter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18286_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00528_),
    .Q(\core.pipe0_fetch.lastProgramCounter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _18287_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_00529_),
    .Q(\core.pipe0_fetch.lastProgramCounter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _18288_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00530_),
    .Q(\core.pipe0_fetch.lastProgramCounter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18289_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00531_),
    .Q(\core.pipe0_fetch.lastProgramCounter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18290_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00532_),
    .Q(\core.pipe0_fetch.lastProgramCounter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18291_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00533_),
    .Q(\core.pipe0_fetch.lastProgramCounter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _18292_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00534_),
    .Q(\core.pipe0_fetch.lastProgramCounter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _18293_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00535_),
    .Q(\core.pipe0_fetch.lastProgramCounter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _18294_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00536_),
    .Q(\core.pipe0_fetch.lastProgramCounter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _18295_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00537_),
    .Q(\core.pipe0_fetch.lastProgramCounter[20] ));
 sky130_fd_sc_hd__dfxtp_1 _18296_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00538_),
    .Q(\core.pipe0_fetch.lastProgramCounter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _18297_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00539_),
    .Q(\core.pipe0_fetch.lastProgramCounter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _18298_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_00540_),
    .Q(\core.pipe0_fetch.lastProgramCounter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _18299_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_00541_),
    .Q(\core.pipe0_fetch.lastProgramCounter[24] ));
 sky130_fd_sc_hd__dfxtp_1 _18300_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00542_),
    .Q(\core.pipe0_fetch.lastProgramCounter[25] ));
 sky130_fd_sc_hd__dfxtp_1 _18301_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00543_),
    .Q(\core.pipe0_fetch.lastProgramCounter[26] ));
 sky130_fd_sc_hd__dfxtp_1 _18302_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00544_),
    .Q(\core.pipe0_fetch.lastProgramCounter[27] ));
 sky130_fd_sc_hd__dfxtp_1 _18303_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00545_),
    .Q(\core.pipe0_fetch.lastProgramCounter[28] ));
 sky130_fd_sc_hd__dfxtp_1 _18304_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00546_),
    .Q(\core.pipe0_fetch.lastProgramCounter[29] ));
 sky130_fd_sc_hd__dfxtp_1 _18305_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00547_),
    .Q(\core.pipe0_fetch.lastProgramCounter[30] ));
 sky130_fd_sc_hd__dfxtp_1 _18306_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_00548_),
    .Q(\core.pipe0_fetch.lastProgramCounter[31] ));
 sky130_fd_sc_hd__dfxtp_1 _18307_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00549_),
    .Q(\core.registers[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18308_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00550_),
    .Q(\core.registers[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18309_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00551_),
    .Q(\core.registers[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18310_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00552_),
    .Q(\core.registers[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18311_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00553_),
    .Q(\core.registers[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18312_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00554_),
    .Q(\core.registers[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18313_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00555_),
    .Q(\core.registers[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18314_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_00556_),
    .Q(\core.registers[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18315_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00557_),
    .Q(\core.registers[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18316_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00558_),
    .Q(\core.registers[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18317_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00559_),
    .Q(\core.registers[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18318_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00560_),
    .Q(\core.registers[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18319_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00561_),
    .Q(\core.registers[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18320_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00562_),
    .Q(\core.registers[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18321_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00563_),
    .Q(\core.registers[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18322_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00564_),
    .Q(\core.registers[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18323_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00565_),
    .Q(\core.registers[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18324_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00566_),
    .Q(\core.registers[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18325_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_00567_),
    .Q(\core.registers[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18326_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00568_),
    .Q(\core.registers[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18327_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_00569_),
    .Q(\core.registers[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18328_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00570_),
    .Q(\core.registers[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18329_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00571_),
    .Q(\core.registers[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18330_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00572_),
    .Q(\core.registers[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18331_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00573_),
    .Q(\core.registers[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18332_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_00574_),
    .Q(\core.registers[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18333_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00575_),
    .Q(\core.registers[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18334_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00576_),
    .Q(\core.registers[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18335_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00577_),
    .Q(\core.registers[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18336_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00578_),
    .Q(\core.registers[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18337_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00579_),
    .Q(\core.registers[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18338_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00580_),
    .Q(\core.registers[18][31] ));
 sky130_fd_sc_hd__dfxtp_4 _18339_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_00581_),
    .Q(\localMemoryInterface.lastRBankSelect ));
 sky130_fd_sc_hd__dfxtp_1 _18340_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00582_),
    .Q(\core.registers[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18341_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00583_),
    .Q(\core.registers[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18342_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00584_),
    .Q(\core.registers[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18343_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00585_),
    .Q(\core.registers[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18344_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00586_),
    .Q(\core.registers[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18345_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00587_),
    .Q(\core.registers[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18346_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00588_),
    .Q(\core.registers[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18347_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_00589_),
    .Q(\core.registers[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18348_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_00590_),
    .Q(\core.registers[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18349_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00591_),
    .Q(\core.registers[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18350_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00592_),
    .Q(\core.registers[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18351_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_00593_),
    .Q(\core.registers[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18352_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00594_),
    .Q(\core.registers[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18353_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_00595_),
    .Q(\core.registers[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18354_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00596_),
    .Q(\core.registers[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18355_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00597_),
    .Q(\core.registers[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18356_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00598_),
    .Q(\core.registers[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18357_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00599_),
    .Q(\core.registers[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18358_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00600_),
    .Q(\core.registers[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18359_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00601_),
    .Q(\core.registers[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18360_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00602_),
    .Q(\core.registers[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18361_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00603_),
    .Q(\core.registers[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18362_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00604_),
    .Q(\core.registers[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18363_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00605_),
    .Q(\core.registers[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18364_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_00606_),
    .Q(\core.registers[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18365_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00607_),
    .Q(\core.registers[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18366_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_00608_),
    .Q(\core.registers[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18367_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00609_),
    .Q(\core.registers[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18368_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00610_),
    .Q(\core.registers[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18369_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00611_),
    .Q(\core.registers[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18370_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00612_),
    .Q(\core.registers[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18371_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_00613_),
    .Q(\core.registers[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _18372_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_00614_),
    .Q(net370));
 sky130_fd_sc_hd__dfxtp_4 _18373_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00615_),
    .Q(\coreWBInterface.readDataBuffered[0] ));
 sky130_fd_sc_hd__dfxtp_4 _18374_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00616_),
    .Q(\coreWBInterface.readDataBuffered[1] ));
 sky130_fd_sc_hd__dfxtp_4 _18375_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_00617_),
    .Q(\coreWBInterface.readDataBuffered[2] ));
 sky130_fd_sc_hd__dfxtp_4 _18376_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00618_),
    .Q(\coreWBInterface.readDataBuffered[3] ));
 sky130_fd_sc_hd__dfxtp_4 _18377_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_00619_),
    .Q(\coreWBInterface.readDataBuffered[4] ));
 sky130_fd_sc_hd__dfxtp_4 _18378_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_00620_),
    .Q(\coreWBInterface.readDataBuffered[5] ));
 sky130_fd_sc_hd__dfxtp_4 _18379_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00621_),
    .Q(\coreWBInterface.readDataBuffered[6] ));
 sky130_fd_sc_hd__dfxtp_4 _18380_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_00622_),
    .Q(\coreWBInterface.readDataBuffered[7] ));
 sky130_fd_sc_hd__dfxtp_4 _18381_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_00623_),
    .Q(\coreWBInterface.readDataBuffered[8] ));
 sky130_fd_sc_hd__dfxtp_4 _18382_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00624_),
    .Q(\coreWBInterface.readDataBuffered[9] ));
 sky130_fd_sc_hd__dfxtp_4 _18383_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00625_),
    .Q(\coreWBInterface.readDataBuffered[10] ));
 sky130_fd_sc_hd__dfxtp_4 _18384_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00626_),
    .Q(\coreWBInterface.readDataBuffered[11] ));
 sky130_fd_sc_hd__dfxtp_4 _18385_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_00627_),
    .Q(\coreWBInterface.readDataBuffered[12] ));
 sky130_fd_sc_hd__dfxtp_4 _18386_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_00628_),
    .Q(\coreWBInterface.readDataBuffered[13] ));
 sky130_fd_sc_hd__dfxtp_4 _18387_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_00629_),
    .Q(\coreWBInterface.readDataBuffered[14] ));
 sky130_fd_sc_hd__dfxtp_4 _18388_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00630_),
    .Q(\coreWBInterface.readDataBuffered[15] ));
 sky130_fd_sc_hd__dfxtp_4 _18389_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00631_),
    .Q(\coreWBInterface.readDataBuffered[16] ));
 sky130_fd_sc_hd__dfxtp_4 _18390_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00632_),
    .Q(\coreWBInterface.readDataBuffered[17] ));
 sky130_fd_sc_hd__dfxtp_4 _18391_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00633_),
    .Q(\coreWBInterface.readDataBuffered[18] ));
 sky130_fd_sc_hd__dfxtp_4 _18392_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00634_),
    .Q(\coreWBInterface.readDataBuffered[19] ));
 sky130_fd_sc_hd__dfxtp_4 _18393_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00635_),
    .Q(\coreWBInterface.readDataBuffered[20] ));
 sky130_fd_sc_hd__dfxtp_4 _18394_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00636_),
    .Q(\coreWBInterface.readDataBuffered[21] ));
 sky130_fd_sc_hd__dfxtp_4 _18395_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00637_),
    .Q(\coreWBInterface.readDataBuffered[22] ));
 sky130_fd_sc_hd__dfxtp_4 _18396_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00638_),
    .Q(\coreWBInterface.readDataBuffered[23] ));
 sky130_fd_sc_hd__dfxtp_4 _18397_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00639_),
    .Q(\coreWBInterface.readDataBuffered[24] ));
 sky130_fd_sc_hd__dfxtp_4 _18398_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00640_),
    .Q(\coreWBInterface.readDataBuffered[25] ));
 sky130_fd_sc_hd__dfxtp_4 _18399_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_00641_),
    .Q(\coreWBInterface.readDataBuffered[26] ));
 sky130_fd_sc_hd__dfxtp_4 _18400_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_00642_),
    .Q(\coreWBInterface.readDataBuffered[27] ));
 sky130_fd_sc_hd__dfxtp_4 _18401_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_00643_),
    .Q(\coreWBInterface.readDataBuffered[28] ));
 sky130_fd_sc_hd__dfxtp_4 _18402_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_00644_),
    .Q(\coreWBInterface.readDataBuffered[29] ));
 sky130_fd_sc_hd__dfxtp_4 _18403_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00645_),
    .Q(\coreWBInterface.readDataBuffered[30] ));
 sky130_fd_sc_hd__dfxtp_4 _18404_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00646_),
    .Q(\coreWBInterface.readDataBuffered[31] ));
 sky130_fd_sc_hd__dfxtp_2 _18405_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_00647_),
    .Q(\coreWBInterface.state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _18406_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_00648_),
    .Q(\coreWBInterface.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18407_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00649_),
    .Q(\core.registers[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18408_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00650_),
    .Q(\core.registers[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18409_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00651_),
    .Q(\core.registers[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18410_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00652_),
    .Q(\core.registers[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18411_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00653_),
    .Q(\core.registers[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18412_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00654_),
    .Q(\core.registers[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18413_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00655_),
    .Q(\core.registers[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18414_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00656_),
    .Q(\core.registers[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18415_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00657_),
    .Q(\core.registers[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18416_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00658_),
    .Q(\core.registers[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18417_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00659_),
    .Q(\core.registers[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18418_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_00660_),
    .Q(\core.registers[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18419_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00661_),
    .Q(\core.registers[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18420_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00662_),
    .Q(\core.registers[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18421_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00663_),
    .Q(\core.registers[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18422_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00664_),
    .Q(\core.registers[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18423_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00665_),
    .Q(\core.registers[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18424_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00666_),
    .Q(\core.registers[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18425_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00667_),
    .Q(\core.registers[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18426_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00668_),
    .Q(\core.registers[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18427_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00669_),
    .Q(\core.registers[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18428_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00670_),
    .Q(\core.registers[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18429_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00671_),
    .Q(\core.registers[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18430_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_00672_),
    .Q(\core.registers[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18431_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00673_),
    .Q(\core.registers[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18432_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00674_),
    .Q(\core.registers[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18433_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00675_),
    .Q(\core.registers[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18434_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00676_),
    .Q(\core.registers[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18435_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_00677_),
    .Q(\core.registers[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18436_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00678_),
    .Q(\core.registers[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18437_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00679_),
    .Q(\core.registers[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18438_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00680_),
    .Q(\core.registers[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18439_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00681_),
    .Q(\core.registers[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18440_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00682_),
    .Q(\core.registers[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18441_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00683_),
    .Q(\core.registers[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18442_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00684_),
    .Q(\core.registers[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18443_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00685_),
    .Q(\core.registers[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18444_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00686_),
    .Q(\core.registers[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18445_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00687_),
    .Q(\core.registers[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18446_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_00688_),
    .Q(\core.registers[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18447_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_00689_),
    .Q(\core.registers[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18448_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00690_),
    .Q(\core.registers[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18449_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00691_),
    .Q(\core.registers[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18450_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00692_),
    .Q(\core.registers[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18451_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_00693_),
    .Q(\core.registers[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18452_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_00694_),
    .Q(\core.registers[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18453_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00695_),
    .Q(\core.registers[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18454_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00696_),
    .Q(\core.registers[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18455_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00697_),
    .Q(\core.registers[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18456_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00698_),
    .Q(\core.registers[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18457_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00699_),
    .Q(\core.registers[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18458_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00700_),
    .Q(\core.registers[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18459_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00701_),
    .Q(\core.registers[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18460_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00702_),
    .Q(\core.registers[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18461_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00703_),
    .Q(\core.registers[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18462_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00704_),
    .Q(\core.registers[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18463_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_00705_),
    .Q(\core.registers[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18464_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_00706_),
    .Q(\core.registers[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18465_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_00707_),
    .Q(\core.registers[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18466_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00708_),
    .Q(\core.registers[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18467_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00709_),
    .Q(\core.registers[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18468_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00710_),
    .Q(\core.registers[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18469_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00711_),
    .Q(\core.registers[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18470_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_00712_),
    .Q(\core.registers[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18471_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00713_),
    .Q(net410));
 sky130_fd_sc_hd__dfxtp_1 _18472_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00714_),
    .Q(net421));
 sky130_fd_sc_hd__dfxtp_1 _18473_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00715_),
    .Q(net432));
 sky130_fd_sc_hd__dfxtp_1 _18474_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00716_),
    .Q(net435));
 sky130_fd_sc_hd__dfxtp_1 _18475_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00717_),
    .Q(net436));
 sky130_fd_sc_hd__dfxtp_1 _18476_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00718_),
    .Q(net437));
 sky130_fd_sc_hd__dfxtp_1 _18477_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00719_),
    .Q(net438));
 sky130_fd_sc_hd__dfxtp_1 _18478_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00720_),
    .Q(net439));
 sky130_fd_sc_hd__dfxtp_1 _18479_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00721_),
    .Q(net440));
 sky130_fd_sc_hd__dfxtp_1 _18480_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00722_),
    .Q(net441));
 sky130_fd_sc_hd__dfxtp_1 _18481_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00723_),
    .Q(net411));
 sky130_fd_sc_hd__dfxtp_1 _18482_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00724_),
    .Q(net412));
 sky130_fd_sc_hd__dfxtp_1 _18483_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00725_),
    .Q(net413));
 sky130_fd_sc_hd__dfxtp_1 _18484_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00726_),
    .Q(net414));
 sky130_fd_sc_hd__dfxtp_1 _18485_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00727_),
    .Q(net415));
 sky130_fd_sc_hd__dfxtp_1 _18486_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00728_),
    .Q(net416));
 sky130_fd_sc_hd__dfxtp_1 _18487_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00729_),
    .Q(net417));
 sky130_fd_sc_hd__dfxtp_1 _18488_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00730_),
    .Q(net418));
 sky130_fd_sc_hd__dfxtp_1 _18489_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00731_),
    .Q(net419));
 sky130_fd_sc_hd__dfxtp_1 _18490_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00732_),
    .Q(net420));
 sky130_fd_sc_hd__dfxtp_1 _18491_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00733_),
    .Q(net422));
 sky130_fd_sc_hd__dfxtp_1 _18492_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00734_),
    .Q(net423));
 sky130_fd_sc_hd__dfxtp_1 _18493_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00735_),
    .Q(net424));
 sky130_fd_sc_hd__dfxtp_1 _18494_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00736_),
    .Q(net425));
 sky130_fd_sc_hd__dfxtp_1 _18495_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00737_),
    .Q(net426));
 sky130_fd_sc_hd__dfxtp_1 _18496_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00738_),
    .Q(net427));
 sky130_fd_sc_hd__dfxtp_1 _18497_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00739_),
    .Q(net428));
 sky130_fd_sc_hd__dfxtp_1 _18498_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00740_),
    .Q(net429));
 sky130_fd_sc_hd__dfxtp_1 _18499_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00741_),
    .Q(net430));
 sky130_fd_sc_hd__dfxtp_1 _18500_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00742_),
    .Q(net431));
 sky130_fd_sc_hd__dfxtp_1 _18501_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00743_),
    .Q(net433));
 sky130_fd_sc_hd__dfxtp_1 _18502_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00744_),
    .Q(net434));
 sky130_fd_sc_hd__dfxtp_1 _18503_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00745_),
    .Q(net409));
 sky130_fd_sc_hd__dfxtp_1 _18504_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00746_),
    .Q(\wbSRAMInterface.currentAddress[0] ));
 sky130_fd_sc_hd__dfxtp_2 _18505_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00747_),
    .Q(\wbSRAMInterface.currentAddress[1] ));
 sky130_fd_sc_hd__dfxtp_4 _18506_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00748_),
    .Q(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__dfxtp_4 _18507_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00749_),
    .Q(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__dfxtp_4 _18508_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00750_),
    .Q(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__dfxtp_4 _18509_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00751_),
    .Q(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__dfxtp_4 _18510_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00752_),
    .Q(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__dfxtp_4 _18511_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00753_),
    .Q(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__dfxtp_4 _18512_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00754_),
    .Q(\wbSRAMInterface.currentAddress[8] ));
 sky130_fd_sc_hd__dfxtp_4 _18513_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00755_),
    .Q(\wbSRAMInterface.currentAddress[9] ));
 sky130_fd_sc_hd__dfxtp_4 _18514_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00756_),
    .Q(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__dfxtp_4 _18515_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00757_),
    .Q(\wbSRAMInterface.currentAddress[11] ));
 sky130_fd_sc_hd__dfxtp_4 _18516_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00758_),
    .Q(\wbSRAMInterface.currentAddress[12] ));
 sky130_fd_sc_hd__dfxtp_2 _18517_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00759_),
    .Q(\wbSRAMInterface.currentAddress[13] ));
 sky130_fd_sc_hd__dfxtp_2 _18518_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00760_),
    .Q(\wbSRAMInterface.currentAddress[14] ));
 sky130_fd_sc_hd__dfxtp_2 _18519_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00761_),
    .Q(\wbSRAMInterface.currentAddress[15] ));
 sky130_fd_sc_hd__dfxtp_2 _18520_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00762_),
    .Q(\wbSRAMInterface.currentAddress[16] ));
 sky130_fd_sc_hd__dfxtp_1 _18521_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00763_),
    .Q(\wbSRAMInterface.currentAddress[17] ));
 sky130_fd_sc_hd__dfxtp_1 _18522_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00764_),
    .Q(\wbSRAMInterface.currentAddress[18] ));
 sky130_fd_sc_hd__dfxtp_1 _18523_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00765_),
    .Q(\wbSRAMInterface.currentAddress[19] ));
 sky130_fd_sc_hd__dfxtp_1 _18524_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00766_),
    .Q(\wbSRAMInterface.currentAddress[20] ));
 sky130_fd_sc_hd__dfxtp_1 _18525_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00767_),
    .Q(\wbSRAMInterface.currentAddress[21] ));
 sky130_fd_sc_hd__dfxtp_1 _18526_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00768_),
    .Q(\wbSRAMInterface.currentAddress[22] ));
 sky130_fd_sc_hd__dfxtp_1 _18527_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00769_),
    .Q(\wbSRAMInterface.currentAddress[23] ));
 sky130_fd_sc_hd__dfxtp_1 _18528_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00770_),
    .Q(\memoryController.last_data_enableWB ));
 sky130_fd_sc_hd__dfxtp_1 _18529_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00771_),
    .Q(net442));
 sky130_fd_sc_hd__dfxtp_4 _18530_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00772_),
    .Q(\wbSRAMInterface.state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _18531_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00773_),
    .Q(\wbSRAMInterface.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18532_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00774_),
    .Q(\core.registers[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18533_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00775_),
    .Q(\core.registers[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18534_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00776_),
    .Q(\core.registers[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18535_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00777_),
    .Q(\core.registers[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18536_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00778_),
    .Q(\core.registers[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18537_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00779_),
    .Q(\core.registers[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18538_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00780_),
    .Q(\core.registers[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18539_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00781_),
    .Q(\core.registers[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18540_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00782_),
    .Q(\core.registers[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18541_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00783_),
    .Q(\core.registers[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18542_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00784_),
    .Q(\core.registers[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18543_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_00785_),
    .Q(\core.registers[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18544_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00786_),
    .Q(\core.registers[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18545_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00787_),
    .Q(\core.registers[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18546_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00788_),
    .Q(\core.registers[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18547_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00789_),
    .Q(\core.registers[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18548_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00790_),
    .Q(\core.registers[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18549_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00791_),
    .Q(\core.registers[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18550_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00792_),
    .Q(\core.registers[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18551_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00793_),
    .Q(\core.registers[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18552_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00794_),
    .Q(\core.registers[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18553_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00795_),
    .Q(\core.registers[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18554_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00796_),
    .Q(\core.registers[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18555_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00797_),
    .Q(\core.registers[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18556_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00798_),
    .Q(\core.registers[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18557_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00799_),
    .Q(\core.registers[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18558_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00800_),
    .Q(\core.registers[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18559_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00801_),
    .Q(\core.registers[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18560_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00802_),
    .Q(\core.registers[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18561_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00803_),
    .Q(\core.registers[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18562_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00804_),
    .Q(\core.registers[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18563_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00805_),
    .Q(\core.registers[16][31] ));
 sky130_fd_sc_hd__dfxtp_4 _18564_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00806_),
    .Q(\core.fetchProgramCounter[2] ));
 sky130_fd_sc_hd__dfxtp_4 _18565_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00807_),
    .Q(\core.fetchProgramCounter[3] ));
 sky130_fd_sc_hd__dfxtp_4 _18566_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_00808_),
    .Q(\core.fetchProgramCounter[4] ));
 sky130_fd_sc_hd__dfxtp_4 _18567_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_00809_),
    .Q(\core.fetchProgramCounter[5] ));
 sky130_fd_sc_hd__dfxtp_4 _18568_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_00810_),
    .Q(\core.fetchProgramCounter[6] ));
 sky130_fd_sc_hd__dfxtp_4 _18569_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00811_),
    .Q(\core.fetchProgramCounter[7] ));
 sky130_fd_sc_hd__dfxtp_4 _18570_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00812_),
    .Q(\core.fetchProgramCounter[8] ));
 sky130_fd_sc_hd__dfxtp_4 _18571_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00813_),
    .Q(\core.fetchProgramCounter[9] ));
 sky130_fd_sc_hd__dfxtp_4 _18572_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00814_),
    .Q(\core.fetchProgramCounter[10] ));
 sky130_fd_sc_hd__dfxtp_4 _18573_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00815_),
    .Q(\core.fetchProgramCounter[11] ));
 sky130_fd_sc_hd__dfxtp_4 _18574_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_00816_),
    .Q(\core.fetchProgramCounter[12] ));
 sky130_fd_sc_hd__dfxtp_4 _18575_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00817_),
    .Q(\core.fetchProgramCounter[13] ));
 sky130_fd_sc_hd__dfxtp_4 _18576_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_00818_),
    .Q(\core.fetchProgramCounter[14] ));
 sky130_fd_sc_hd__dfxtp_4 _18577_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_00819_),
    .Q(\core.fetchProgramCounter[15] ));
 sky130_fd_sc_hd__dfxtp_2 _18578_ (.CLK(clknet_leaf_161_wb_clk_i),
    .D(_00820_),
    .Q(\core.fetchProgramCounter[16] ));
 sky130_fd_sc_hd__dfxtp_4 _18579_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00821_),
    .Q(\core.fetchProgramCounter[17] ));
 sky130_fd_sc_hd__dfxtp_4 _18580_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_00822_),
    .Q(\core.fetchProgramCounter[18] ));
 sky130_fd_sc_hd__dfxtp_4 _18581_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_00823_),
    .Q(\core.fetchProgramCounter[19] ));
 sky130_fd_sc_hd__dfxtp_4 _18582_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_00824_),
    .Q(\core.fetchProgramCounter[20] ));
 sky130_fd_sc_hd__dfxtp_4 _18583_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_00825_),
    .Q(\core.fetchProgramCounter[21] ));
 sky130_fd_sc_hd__dfxtp_4 _18584_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_00826_),
    .Q(\core.fetchProgramCounter[22] ));
 sky130_fd_sc_hd__dfxtp_4 _18585_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_00827_),
    .Q(\core.fetchProgramCounter[23] ));
 sky130_fd_sc_hd__dfxtp_4 _18586_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_00828_),
    .Q(\core.fetchProgramCounter[24] ));
 sky130_fd_sc_hd__dfxtp_4 _18587_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_00829_),
    .Q(\core.fetchProgramCounter[25] ));
 sky130_fd_sc_hd__dfxtp_4 _18588_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_00830_),
    .Q(\core.fetchProgramCounter[26] ));
 sky130_fd_sc_hd__dfxtp_4 _18589_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_00831_),
    .Q(\core.fetchProgramCounter[27] ));
 sky130_fd_sc_hd__dfxtp_4 _18590_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00832_),
    .Q(\core.fetchProgramCounter[28] ));
 sky130_fd_sc_hd__dfxtp_4 _18591_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00833_),
    .Q(\core.fetchProgramCounter[29] ));
 sky130_fd_sc_hd__dfxtp_4 _18592_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_00834_),
    .Q(\core.fetchProgramCounter[30] ));
 sky130_fd_sc_hd__dfxtp_2 _18593_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00835_),
    .Q(\core.fetchProgramCounter[31] ));
 sky130_fd_sc_hd__dfxtp_1 _18594_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00836_),
    .Q(\core.registers[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18595_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00837_),
    .Q(\core.registers[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18596_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_00838_),
    .Q(\core.registers[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18597_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00839_),
    .Q(\core.registers[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18598_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00840_),
    .Q(\core.registers[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18599_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00841_),
    .Q(\core.registers[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18600_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00842_),
    .Q(\core.registers[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18601_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00843_),
    .Q(\core.registers[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18602_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00844_),
    .Q(\core.registers[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18603_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00845_),
    .Q(\core.registers[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18604_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00846_),
    .Q(\core.registers[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18605_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_00847_),
    .Q(\core.registers[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18606_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00848_),
    .Q(\core.registers[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18607_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00849_),
    .Q(\core.registers[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18608_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00850_),
    .Q(\core.registers[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18609_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00851_),
    .Q(\core.registers[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18610_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00852_),
    .Q(\core.registers[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18611_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00853_),
    .Q(\core.registers[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18612_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00854_),
    .Q(\core.registers[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18613_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00855_),
    .Q(\core.registers[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18614_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_00856_),
    .Q(\core.registers[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18615_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_00857_),
    .Q(\core.registers[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18616_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00858_),
    .Q(\core.registers[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18617_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00859_),
    .Q(\core.registers[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18618_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00860_),
    .Q(\core.registers[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18619_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_00861_),
    .Q(\core.registers[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18620_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_00862_),
    .Q(\core.registers[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18621_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00863_),
    .Q(\core.registers[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18622_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00864_),
    .Q(\core.registers[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18623_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00865_),
    .Q(\core.registers[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18624_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00866_),
    .Q(\core.registers[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18625_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_00867_),
    .Q(\core.registers[10][31] ));
 sky130_fd_sc_hd__dfxtp_4 _18626_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00868_),
    .Q(\core.registers[0][0] ));
 sky130_fd_sc_hd__dfxtp_4 _18627_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00869_),
    .Q(\core.registers[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _18628_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00870_),
    .Q(\core.registers[0][2] ));
 sky130_fd_sc_hd__dfxtp_4 _18629_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00871_),
    .Q(\core.registers[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _18630_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00872_),
    .Q(\core.registers[0][4] ));
 sky130_fd_sc_hd__dfxtp_4 _18631_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00873_),
    .Q(\core.registers[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _18632_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00874_),
    .Q(\core.registers[0][6] ));
 sky130_fd_sc_hd__dfxtp_4 _18633_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00875_),
    .Q(\core.registers[0][7] ));
 sky130_fd_sc_hd__dfxtp_4 _18634_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00876_),
    .Q(\core.registers[0][8] ));
 sky130_fd_sc_hd__dfxtp_4 _18635_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00877_),
    .Q(\core.registers[0][9] ));
 sky130_fd_sc_hd__dfxtp_4 _18636_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00878_),
    .Q(\core.registers[0][10] ));
 sky130_fd_sc_hd__dfxtp_4 _18637_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00879_),
    .Q(\core.registers[0][11] ));
 sky130_fd_sc_hd__dfxtp_4 _18638_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00880_),
    .Q(\core.registers[0][12] ));
 sky130_fd_sc_hd__dfxtp_4 _18639_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00881_),
    .Q(\core.registers[0][13] ));
 sky130_fd_sc_hd__dfxtp_4 _18640_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00882_),
    .Q(\core.registers[0][14] ));
 sky130_fd_sc_hd__dfxtp_4 _18641_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00883_),
    .Q(\core.registers[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _18642_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_00884_),
    .Q(\core.registers[0][16] ));
 sky130_fd_sc_hd__dfxtp_4 _18643_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00885_),
    .Q(\core.registers[0][17] ));
 sky130_fd_sc_hd__dfxtp_4 _18644_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00886_),
    .Q(\core.registers[0][18] ));
 sky130_fd_sc_hd__dfxtp_4 _18645_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00887_),
    .Q(\core.registers[0][19] ));
 sky130_fd_sc_hd__dfxtp_4 _18646_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_00888_),
    .Q(\core.registers[0][20] ));
 sky130_fd_sc_hd__dfxtp_4 _18647_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00889_),
    .Q(\core.registers[0][21] ));
 sky130_fd_sc_hd__dfxtp_4 _18648_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00890_),
    .Q(\core.registers[0][22] ));
 sky130_fd_sc_hd__dfxtp_4 _18649_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00891_),
    .Q(\core.registers[0][23] ));
 sky130_fd_sc_hd__dfxtp_4 _18650_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00892_),
    .Q(\core.registers[0][24] ));
 sky130_fd_sc_hd__dfxtp_4 _18651_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00893_),
    .Q(\core.registers[0][25] ));
 sky130_fd_sc_hd__dfxtp_4 _18652_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00894_),
    .Q(\core.registers[0][26] ));
 sky130_fd_sc_hd__dfxtp_4 _18653_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00895_),
    .Q(\core.registers[0][27] ));
 sky130_fd_sc_hd__dfxtp_4 _18654_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00896_),
    .Q(\core.registers[0][28] ));
 sky130_fd_sc_hd__dfxtp_4 _18655_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00897_),
    .Q(\core.registers[0][29] ));
 sky130_fd_sc_hd__dfxtp_4 _18656_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00898_),
    .Q(\core.registers[0][30] ));
 sky130_fd_sc_hd__dfxtp_4 _18657_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00899_),
    .Q(\core.registers[0][31] ));
 sky130_fd_sc_hd__dfxtp_4 _18658_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00900_),
    .Q(\core.management_interruptEnable ));
 sky130_fd_sc_hd__dfxtp_1 _18659_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00901_),
    .Q(\coreManagement.control[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18660_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00902_),
    .Q(\core.management_run ));
 sky130_fd_sc_hd__dfxtp_1 _18661_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00903_),
    .Q(\jtag.dataIDRegister.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18662_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00904_),
    .Q(\jtag.dataIDRegister.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18663_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00905_),
    .Q(\jtag.dataIDRegister.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18664_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00906_),
    .Q(\jtag.dataIDRegister.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18665_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00907_),
    .Q(\jtag.dataIDRegister.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18666_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00908_),
    .Q(\jtag.dataIDRegister.data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18667_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00909_),
    .Q(\jtag.dataIDRegister.data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18668_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00910_),
    .Q(\jtag.dataIDRegister.data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18669_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00911_),
    .Q(\jtag.dataIDRegister.data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18670_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00912_),
    .Q(\jtag.dataIDRegister.data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _18671_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00913_),
    .Q(\jtag.dataIDRegister.data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18672_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00914_),
    .Q(\jtag.dataIDRegister.data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _18673_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00915_),
    .Q(\jtag.dataIDRegister.data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _18674_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00916_),
    .Q(\jtag.dataIDRegister.data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18675_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00917_),
    .Q(\jtag.dataIDRegister.data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18676_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00918_),
    .Q(\jtag.dataIDRegister.data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18677_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00919_),
    .Q(\jtag.dataIDRegister.data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _18678_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00920_),
    .Q(\jtag.dataIDRegister.data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _18679_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00921_),
    .Q(\jtag.dataIDRegister.data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _18680_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00922_),
    .Q(\jtag.dataIDRegister.data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _18681_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00923_),
    .Q(\jtag.dataIDRegister.data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _18682_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00924_),
    .Q(\jtag.dataIDRegister.data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _18683_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00925_),
    .Q(\jtag.dataIDRegister.data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _18684_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00926_),
    .Q(\jtag.dataIDRegister.data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _18685_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00927_),
    .Q(\jtag.dataIDRegister.data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _18686_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00928_),
    .Q(\jtag.dataIDRegister.data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _18687_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00929_),
    .Q(\jtag.dataIDRegister.data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _18688_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00930_),
    .Q(\jtag.dataIDRegister.data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _18689_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00931_),
    .Q(\jtag.dataIDRegister.data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _18690_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00932_),
    .Q(\jtag.dataIDRegister.data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _18691_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00933_),
    .Q(\jtag.dataIDRegister.data[30] ));
 sky130_fd_sc_hd__dfxtp_4 _18692_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00934_),
    .Q(\jtag.dataIDRegister.data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _18693_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00935_),
    .Q(\jtag.dataBypassRegister.data ));
 sky130_fd_sc_hd__dfxtp_1 _18694_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00936_),
    .Q(\jtag.dataBSRRegister.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18695_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00937_),
    .Q(\jtag.dataBSRRegister.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18696_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00938_),
    .Q(\jtag.dataBSRRegister.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18697_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00939_),
    .Q(\jtag.dataBSRRegister.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18698_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00940_),
    .Q(\jtag.dataBSRRegister.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18699_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00941_),
    .Q(\jtag.dataBSRRegister.data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18700_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00942_),
    .Q(\jtag.dataBSRRegister.data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18701_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00943_),
    .Q(\jtag.dataBSRRegister.data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18702_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00944_),
    .Q(\jtag.dataBSRRegister.data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18703_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00945_),
    .Q(\jtag.dataBSRRegister.data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _18704_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00946_),
    .Q(\jtag.dataBSRRegister.data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18705_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00947_),
    .Q(\jtag.dataBSRRegister.data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _18706_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00948_),
    .Q(\jtag.dataBSRRegister.data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _18707_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00949_),
    .Q(\jtag.dataBSRRegister.data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18708_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00950_),
    .Q(\jtag.dataBSRRegister.data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18709_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00951_),
    .Q(\jtag.dataBSRRegister.data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18710_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00952_),
    .Q(\jtag.dataBSRRegister.data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _18711_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00953_),
    .Q(\jtag.dataBSRRegister.data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _18712_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00954_),
    .Q(\jtag.dataBSRRegister.data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _18713_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00955_),
    .Q(\jtag.dataBSRRegister.data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _18714_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00956_),
    .Q(\jtag.dataBSRRegister.data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _18715_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00957_),
    .Q(\jtag.dataBSRRegister.data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _18716_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00958_),
    .Q(\jtag.dataBSRRegister.data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _18717_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00959_),
    .Q(\jtag.dataBSRRegister.data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _18718_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_00960_),
    .Q(\jtag.dataBSRRegister.data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _18719_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_00961_),
    .Q(\jtag.dataBSRRegister.data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _18720_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_00962_),
    .Q(\jtag.dataBSRRegister.data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _18721_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_00963_),
    .Q(\jtag.dataBSRRegister.data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _18722_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_00964_),
    .Q(\jtag.dataBSRRegister.data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _18723_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00965_),
    .Q(\jtag.dataBSRRegister.data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _18724_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00966_),
    .Q(\jtag.dataBSRRegister.data[30] ));
 sky130_fd_sc_hd__dfxtp_4 _18725_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00967_),
    .Q(\jtag.dataBSRRegister.data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _18726_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00968_),
    .Q(\jtag.instructionRegister.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18727_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00969_),
    .Q(\jtag.instructionRegister.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18728_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00970_),
    .Q(\jtag.instructionRegister.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18729_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00971_),
    .Q(\jtag.instructionRegister.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18730_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00972_),
    .Q(\jtag.instructionRegister.data[4] ));
 sky130_fd_sc_hd__dfxtp_4 _18731_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00973_),
    .Q(\jtag.tckRisingEdge ));
 sky130_fd_sc_hd__dfxtp_1 _18732_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00974_),
    .Q(\jtag.tckState ));
 sky130_fd_sc_hd__dfxtp_4 _18733_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00975_),
    .Q(net445));
 sky130_fd_sc_hd__dfxtp_4 _18734_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00976_),
    .Q(net446));
 sky130_fd_sc_hd__dfxtp_4 _18735_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00977_),
    .Q(net447));
 sky130_fd_sc_hd__dfxtp_4 _18736_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00978_),
    .Q(net448));
 sky130_fd_sc_hd__dfxtp_4 _18737_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00979_),
    .Q(net449));
 sky130_fd_sc_hd__dfxtp_2 _18738_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00980_),
    .Q(\jtag.state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _18739_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00981_),
    .Q(\jtag.state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _18740_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00982_),
    .Q(\jtag.state[2] ));
 sky130_fd_sc_hd__dfxtp_2 _18741_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00983_),
    .Q(\jtag.state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _18742_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00984_),
    .Q(\jtag.managementReadData[0] ));
 sky130_fd_sc_hd__dfxtp_2 _18743_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00985_),
    .Q(\jtag.managementReadData[1] ));
 sky130_fd_sc_hd__dfxtp_2 _18744_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00986_),
    .Q(\jtag.managementReadData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18745_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00987_),
    .Q(\jtag.managementReadData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18746_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00988_),
    .Q(\jtag.managementReadData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18747_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00989_),
    .Q(\jtag.managementReadData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18748_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00990_),
    .Q(\jtag.managementReadData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18749_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00991_),
    .Q(\jtag.managementReadData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18750_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00992_),
    .Q(\jtag.managementReadData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18751_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00993_),
    .Q(\jtag.managementReadData[9] ));
 sky130_fd_sc_hd__dfxtp_1 _18752_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00994_),
    .Q(\jtag.managementReadData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18753_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00995_),
    .Q(\jtag.managementReadData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _18754_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00996_),
    .Q(\jtag.managementReadData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _18755_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00997_),
    .Q(\jtag.managementReadData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18756_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00998_),
    .Q(\jtag.managementReadData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18757_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00999_),
    .Q(\jtag.managementReadData[15] ));
 sky130_fd_sc_hd__dfxtp_2 _18758_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_01000_),
    .Q(\jtag.managementReadData[16] ));
 sky130_fd_sc_hd__dfxtp_2 _18759_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_01001_),
    .Q(\jtag.managementReadData[17] ));
 sky130_fd_sc_hd__dfxtp_2 _18760_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01002_),
    .Q(\jtag.managementReadData[18] ));
 sky130_fd_sc_hd__dfxtp_2 _18761_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_01003_),
    .Q(\jtag.managementReadData[19] ));
 sky130_fd_sc_hd__dfxtp_2 _18762_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01004_),
    .Q(\jtag.managementReadData[20] ));
 sky130_fd_sc_hd__dfxtp_2 _18763_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01005_),
    .Q(\jtag.managementReadData[21] ));
 sky130_fd_sc_hd__dfxtp_2 _18764_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01006_),
    .Q(\jtag.managementReadData[22] ));
 sky130_fd_sc_hd__dfxtp_2 _18765_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01007_),
    .Q(\jtag.managementReadData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _18766_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01008_),
    .Q(\jtag.managementReadData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _18767_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01009_),
    .Q(\jtag.managementReadData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _18768_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01010_),
    .Q(\jtag.managementReadData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _18769_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01011_),
    .Q(\jtag.managementReadData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _18770_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01012_),
    .Q(\jtag.managementReadData[28] ));
 sky130_fd_sc_hd__dfxtp_2 _18771_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01013_),
    .Q(\jtag.managementReadData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _18772_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01014_),
    .Q(\jtag.managementReadData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _18773_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01015_),
    .Q(\jtag.managementReadData[31] ));
 sky130_fd_sc_hd__dfxtp_2 _18774_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01016_),
    .Q(\jtag.managementState[0] ));
 sky130_fd_sc_hd__dfxtp_2 _18775_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01017_),
    .Q(\jtag.managementState[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18776_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_01018_),
    .Q(\jtag.managementState[2] ));
 sky130_fd_sc_hd__dfxtp_4 _18777_ (.CLK(clknet_leaf_145_wb_clk_i),
    .D(_01019_),
    .Q(\core.fetchProgramCounter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _18778_ (.CLK(clknet_leaf_145_wb_clk_i),
    .D(_01020_),
    .Q(\core.fetchProgramCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18779_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01021_),
    .Q(\core.registers[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18780_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01022_),
    .Q(\core.registers[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18781_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_01023_),
    .Q(\core.registers[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18782_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01024_),
    .Q(\core.registers[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18783_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01025_),
    .Q(\core.registers[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18784_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01026_),
    .Q(\core.registers[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18785_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_01027_),
    .Q(\core.registers[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18786_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01028_),
    .Q(\core.registers[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18787_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01029_),
    .Q(\core.registers[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18788_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01030_),
    .Q(\core.registers[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18789_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01031_),
    .Q(\core.registers[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18790_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01032_),
    .Q(\core.registers[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18791_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01033_),
    .Q(\core.registers[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18792_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01034_),
    .Q(\core.registers[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18793_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_01035_),
    .Q(\core.registers[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18794_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_01036_),
    .Q(\core.registers[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18795_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01037_),
    .Q(\core.registers[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18796_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01038_),
    .Q(\core.registers[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18797_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_01039_),
    .Q(\core.registers[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18798_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01040_),
    .Q(\core.registers[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18799_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01041_),
    .Q(\core.registers[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18800_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01042_),
    .Q(\core.registers[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18801_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_01043_),
    .Q(\core.registers[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18802_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_01044_),
    .Q(\core.registers[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18803_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_01045_),
    .Q(\core.registers[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18804_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_01046_),
    .Q(\core.registers[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18805_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01047_),
    .Q(\core.registers[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18806_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01048_),
    .Q(\core.registers[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18807_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01049_),
    .Q(\core.registers[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18808_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01050_),
    .Q(\core.registers[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18809_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01051_),
    .Q(\core.registers[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18810_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01052_),
    .Q(\core.registers[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18811_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01053_),
    .Q(\core.registers[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18812_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01054_),
    .Q(\core.registers[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18813_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01055_),
    .Q(\core.registers[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18814_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01056_),
    .Q(\core.registers[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18815_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01057_),
    .Q(\core.registers[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18816_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01058_),
    .Q(\core.registers[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18817_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_01059_),
    .Q(\core.registers[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18818_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01060_),
    .Q(\core.registers[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18819_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01061_),
    .Q(\core.registers[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18820_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01062_),
    .Q(\core.registers[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18821_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01063_),
    .Q(\core.registers[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18822_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01064_),
    .Q(\core.registers[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18823_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01065_),
    .Q(\core.registers[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18824_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01066_),
    .Q(\core.registers[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18825_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01067_),
    .Q(\core.registers[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18826_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01068_),
    .Q(\core.registers[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18827_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_01069_),
    .Q(\core.registers[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18828_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01070_),
    .Q(\core.registers[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18829_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01071_),
    .Q(\core.registers[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18830_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01072_),
    .Q(\core.registers[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18831_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_01073_),
    .Q(\core.registers[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18832_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01074_),
    .Q(\core.registers[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18833_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_01075_),
    .Q(\core.registers[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18834_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_01076_),
    .Q(\core.registers[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18835_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_01077_),
    .Q(\core.registers[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18836_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_01078_),
    .Q(\core.registers[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18837_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01079_),
    .Q(\core.registers[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18838_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01080_),
    .Q(\core.registers[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18839_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01081_),
    .Q(\core.registers[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18840_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_01082_),
    .Q(\core.registers[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18841_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01083_),
    .Q(\core.registers[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18842_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01084_),
    .Q(\core.registers[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18843_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01085_),
    .Q(\core.registers[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18844_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01086_),
    .Q(\core.registers[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18845_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01087_),
    .Q(\core.registers[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18846_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01088_),
    .Q(\core.registers[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18847_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01089_),
    .Q(\core.registers[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18848_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01090_),
    .Q(\core.registers[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18849_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_01091_),
    .Q(\core.registers[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18850_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01092_),
    .Q(\core.registers[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18851_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01093_),
    .Q(\core.registers[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18852_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01094_),
    .Q(\core.registers[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18853_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01095_),
    .Q(\core.registers[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18854_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01096_),
    .Q(\core.registers[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18855_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01097_),
    .Q(\core.registers[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18856_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01098_),
    .Q(\core.registers[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18857_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_01099_),
    .Q(\core.registers[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18858_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01100_),
    .Q(\core.registers[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18859_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_01101_),
    .Q(\core.registers[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18860_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_01102_),
    .Q(\core.registers[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18861_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01103_),
    .Q(\core.registers[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18862_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01104_),
    .Q(\core.registers[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18863_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01105_),
    .Q(\core.registers[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18864_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01106_),
    .Q(\core.registers[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18865_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01107_),
    .Q(\core.registers[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18866_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_01108_),
    .Q(\core.registers[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18867_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01109_),
    .Q(\core.registers[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18868_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_01110_),
    .Q(\core.registers[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18869_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01111_),
    .Q(\core.registers[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18870_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01112_),
    .Q(\core.registers[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18871_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01113_),
    .Q(\core.registers[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18872_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_01114_),
    .Q(\core.registers[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18873_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_01115_),
    .Q(\core.registers[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18874_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01116_),
    .Q(\core.registers[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18875_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01117_),
    .Q(\core.registers[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18876_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01118_),
    .Q(\core.registers[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18877_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01119_),
    .Q(\core.registers[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18878_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01120_),
    .Q(\core.registers[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18879_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01121_),
    .Q(\core.registers[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18880_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01122_),
    .Q(\core.registers[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18881_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_01123_),
    .Q(\core.registers[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18882_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01124_),
    .Q(\core.registers[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18883_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01125_),
    .Q(\core.registers[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18884_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01126_),
    .Q(\core.registers[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18885_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01127_),
    .Q(\core.registers[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18886_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01128_),
    .Q(\core.registers[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18887_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01129_),
    .Q(\core.registers[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18888_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01130_),
    .Q(\core.registers[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18889_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_01131_),
    .Q(\core.registers[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18890_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01132_),
    .Q(\core.registers[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18891_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01133_),
    .Q(\core.registers[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18892_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01134_),
    .Q(\core.registers[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18893_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01135_),
    .Q(\core.registers[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18894_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01136_),
    .Q(\core.registers[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18895_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01137_),
    .Q(\core.registers[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18896_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01138_),
    .Q(\core.registers[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18897_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01139_),
    .Q(\core.registers[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18898_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_01140_),
    .Q(\core.registers[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18899_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01141_),
    .Q(\core.registers[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18900_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_01142_),
    .Q(\core.registers[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18901_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01143_),
    .Q(\core.registers[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18902_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01144_),
    .Q(\core.registers[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18903_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01145_),
    .Q(\core.registers[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18904_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_01146_),
    .Q(\core.registers[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18905_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_01147_),
    .Q(\core.registers[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18906_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01148_),
    .Q(\core.registers[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18907_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01149_),
    .Q(\core.registers[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18908_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01150_),
    .Q(\core.registers[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18909_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01151_),
    .Q(\core.registers[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18910_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01152_),
    .Q(\core.registers[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18911_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01153_),
    .Q(\core.registers[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18912_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01154_),
    .Q(\core.registers[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18913_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_01155_),
    .Q(\core.registers[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18914_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01156_),
    .Q(\core.registers[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18915_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01157_),
    .Q(\core.registers[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18916_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01158_),
    .Q(\core.registers[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18917_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01159_),
    .Q(\core.registers[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18918_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01160_),
    .Q(\core.registers[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18919_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01161_),
    .Q(\core.registers[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18920_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01162_),
    .Q(\core.registers[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18921_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01163_),
    .Q(\core.registers[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18922_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01164_),
    .Q(\core.registers[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18923_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_01165_),
    .Q(\core.registers[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18924_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01166_),
    .Q(\core.registers[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18925_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01167_),
    .Q(\core.registers[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18926_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01168_),
    .Q(\core.registers[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18927_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_01169_),
    .Q(\core.registers[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18928_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01170_),
    .Q(\core.registers[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18929_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01171_),
    .Q(\core.registers[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18930_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_01172_),
    .Q(\core.registers[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18931_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_01173_),
    .Q(\core.registers[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18932_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_01174_),
    .Q(\core.registers[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18933_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_01175_),
    .Q(\core.registers[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18934_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_01176_),
    .Q(\core.registers[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18935_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01177_),
    .Q(\core.registers[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18936_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01178_),
    .Q(\core.registers[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18937_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_01179_),
    .Q(\core.registers[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18938_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_01180_),
    .Q(\core.registers[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18939_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_01181_),
    .Q(\core.registers[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18940_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01182_),
    .Q(\core.registers[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18941_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01183_),
    .Q(\core.registers[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18942_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_01184_),
    .Q(\core.registers[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18943_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01185_),
    .Q(\core.registers[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18944_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01186_),
    .Q(\core.registers[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18945_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01187_),
    .Q(\core.registers[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18946_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01188_),
    .Q(\core.registers[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18947_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01189_),
    .Q(\core.registers[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18948_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01190_),
    .Q(\core.registers[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18949_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01191_),
    .Q(\core.registers[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18950_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_01192_),
    .Q(\core.registers[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18951_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01193_),
    .Q(\core.registers[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18952_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01194_),
    .Q(\core.registers[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18953_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_01195_),
    .Q(\core.registers[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18954_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01196_),
    .Q(\core.registers[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18955_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01197_),
    .Q(\core.registers[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18956_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01198_),
    .Q(\core.registers[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18957_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01199_),
    .Q(\core.registers[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18958_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01200_),
    .Q(\core.registers[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18959_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01201_),
    .Q(\core.registers[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18960_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_01202_),
    .Q(\core.registers[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18961_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_01203_),
    .Q(\core.registers[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18962_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_01204_),
    .Q(\core.registers[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18963_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_01205_),
    .Q(\core.registers[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18964_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01206_),
    .Q(\core.registers[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18965_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_01207_),
    .Q(\core.registers[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18966_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01208_),
    .Q(\core.registers[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18967_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01209_),
    .Q(\core.registers[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18968_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01210_),
    .Q(\core.registers[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18969_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_01211_),
    .Q(\core.registers[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18970_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_01212_),
    .Q(\core.registers[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18971_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01213_),
    .Q(\core.registers[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18972_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_01214_),
    .Q(\core.registers[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18973_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_01215_),
    .Q(\core.registers[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18974_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_01216_),
    .Q(\core.registers[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18975_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01217_),
    .Q(\core.registers[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18976_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01218_),
    .Q(\core.registers[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18977_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01219_),
    .Q(\core.registers[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18978_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01220_),
    .Q(\core.registers[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18979_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01221_),
    .Q(\core.registers[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18980_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01222_),
    .Q(\core.registers[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18981_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01223_),
    .Q(\core.registers[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18982_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01224_),
    .Q(\core.registers[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18983_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_01225_),
    .Q(\core.registers[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18984_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01226_),
    .Q(\core.registers[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18985_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01227_),
    .Q(\core.registers[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18986_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01228_),
    .Q(\core.registers[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18987_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_01229_),
    .Q(\core.registers[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18988_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01230_),
    .Q(\core.registers[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18989_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01231_),
    .Q(\core.registers[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18990_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01232_),
    .Q(\core.registers[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18991_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_01233_),
    .Q(\core.registers[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18992_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_01234_),
    .Q(\core.registers[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18993_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_01235_),
    .Q(\core.registers[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18994_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_01236_),
    .Q(\core.registers[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18995_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_01237_),
    .Q(\core.registers[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18996_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_01238_),
    .Q(\core.registers[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18997_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_01239_),
    .Q(\core.registers[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18998_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01240_),
    .Q(\core.registers[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18999_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01241_),
    .Q(\core.registers[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19000_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01242_),
    .Q(\core.registers[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19001_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_01243_),
    .Q(\core.registers[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19002_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_01244_),
    .Q(\core.registers[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19003_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01245_),
    .Q(\core.registers[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19004_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01246_),
    .Q(\core.registers[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19005_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01247_),
    .Q(\core.registers[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19006_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01248_),
    .Q(\core.registers[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19007_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01249_),
    .Q(\core.registers[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19008_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01250_),
    .Q(\core.registers[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19009_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_01251_),
    .Q(\core.registers[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19010_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01252_),
    .Q(\core.registers[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19011_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01253_),
    .Q(\core.registers[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19012_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01254_),
    .Q(\core.registers[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19013_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01255_),
    .Q(\core.registers[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19014_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01256_),
    .Q(\core.registers[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19015_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_01257_),
    .Q(\core.registers[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19016_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01258_),
    .Q(\core.registers[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19017_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_01259_),
    .Q(\core.registers[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19018_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01260_),
    .Q(\core.registers[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19019_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01261_),
    .Q(\core.registers[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19020_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01262_),
    .Q(\core.registers[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19021_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01263_),
    .Q(\core.registers[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19022_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01264_),
    .Q(\core.registers[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19023_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01265_),
    .Q(\core.registers[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19024_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01266_),
    .Q(\core.registers[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19025_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_01267_),
    .Q(\core.registers[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19026_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01268_),
    .Q(\core.registers[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19027_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01269_),
    .Q(\core.registers[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19028_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_01270_),
    .Q(\core.registers[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19029_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01271_),
    .Q(\core.registers[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19030_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01272_),
    .Q(\core.registers[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19031_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01273_),
    .Q(\core.registers[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19032_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01274_),
    .Q(\core.registers[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19033_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01275_),
    .Q(\core.registers[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19034_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01276_),
    .Q(\core.registers[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19035_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01277_),
    .Q(\core.registers[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19036_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01278_),
    .Q(\core.registers[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19037_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01279_),
    .Q(\core.registers[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19038_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01280_),
    .Q(\core.registers[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19039_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01281_),
    .Q(\core.registers[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19040_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01282_),
    .Q(\core.registers[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19041_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_01283_),
    .Q(\core.registers[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19042_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01284_),
    .Q(\core.registers[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19043_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01285_),
    .Q(\core.registers[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19044_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01286_),
    .Q(\core.registers[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19045_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01287_),
    .Q(\core.registers[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19046_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01288_),
    .Q(\core.registers[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19047_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_01289_),
    .Q(\core.registers[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19048_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01290_),
    .Q(\core.registers[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19049_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_01291_),
    .Q(\core.registers[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19050_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01292_),
    .Q(\core.registers[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19051_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01293_),
    .Q(\core.registers[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19052_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01294_),
    .Q(\core.registers[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19053_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01295_),
    .Q(\core.registers[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19054_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01296_),
    .Q(\core.registers[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19055_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01297_),
    .Q(\core.registers[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19056_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01298_),
    .Q(\core.registers[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19057_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01299_),
    .Q(\core.registers[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19058_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01300_),
    .Q(\core.registers[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19059_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_01301_),
    .Q(\core.registers[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19060_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_01302_),
    .Q(\core.registers[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19061_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01303_),
    .Q(\core.registers[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19062_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_01304_),
    .Q(\core.registers[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19063_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01305_),
    .Q(\core.registers[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19064_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01306_),
    .Q(\core.registers[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19065_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01307_),
    .Q(\core.registers[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19066_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01308_),
    .Q(\core.registers[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19067_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01309_),
    .Q(\core.registers[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19068_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01310_),
    .Q(\core.registers[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19069_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01311_),
    .Q(\core.registers[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19070_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_01312_),
    .Q(\core.registers[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19071_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_01313_),
    .Q(\core.registers[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19072_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01314_),
    .Q(\core.registers[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19073_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01315_),
    .Q(\core.registers[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19074_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01316_),
    .Q(\core.registers[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19075_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01317_),
    .Q(\core.registers[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19076_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01318_),
    .Q(\core.registers[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19077_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01319_),
    .Q(\core.registers[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19078_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01320_),
    .Q(\core.registers[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19079_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_01321_),
    .Q(\core.registers[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19080_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01322_),
    .Q(\core.registers[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19081_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01323_),
    .Q(\core.registers[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19082_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_01324_),
    .Q(\core.registers[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19083_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_01325_),
    .Q(\core.registers[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19084_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01326_),
    .Q(\core.registers[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19085_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01327_),
    .Q(\core.registers[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19086_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01328_),
    .Q(\core.registers[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19087_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01329_),
    .Q(\core.registers[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19088_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_01330_),
    .Q(\core.registers[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19089_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01331_),
    .Q(\core.registers[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19090_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_01332_),
    .Q(\core.registers[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19091_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_01333_),
    .Q(\core.registers[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19092_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_01334_),
    .Q(\core.registers[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19093_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_01335_),
    .Q(\core.registers[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19094_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01336_),
    .Q(\core.registers[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19095_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01337_),
    .Q(\core.registers[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19096_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01338_),
    .Q(\core.registers[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19097_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01339_),
    .Q(\core.registers[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19098_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_01340_),
    .Q(\core.registers[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19099_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_01341_),
    .Q(\core.registers[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19100_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01342_),
    .Q(\core.registers[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19101_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01343_),
    .Q(\core.registers[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19102_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_01344_),
    .Q(\core.registers[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19103_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01345_),
    .Q(\core.registers[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19104_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01346_),
    .Q(\core.registers[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19105_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01347_),
    .Q(\core.registers[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19106_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01348_),
    .Q(\core.registers[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19107_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01349_),
    .Q(\core.registers[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19108_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01350_),
    .Q(\core.registers[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19109_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01351_),
    .Q(\core.registers[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19110_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_01352_),
    .Q(\core.registers[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19111_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_01353_),
    .Q(\core.registers[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19112_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01354_),
    .Q(\core.registers[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19113_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_01355_),
    .Q(\core.registers[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19114_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_01356_),
    .Q(\core.registers[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19115_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01357_),
    .Q(\core.registers[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19116_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_01358_),
    .Q(\core.registers[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19117_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01359_),
    .Q(\core.registers[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19118_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01360_),
    .Q(\core.registers[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19119_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01361_),
    .Q(\core.registers[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19120_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_01362_),
    .Q(\core.registers[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19121_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_01363_),
    .Q(\core.registers[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19122_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_01364_),
    .Q(\core.registers[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19123_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_01365_),
    .Q(\core.registers[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19124_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01366_),
    .Q(\core.registers[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19125_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_01367_),
    .Q(\core.registers[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19126_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01368_),
    .Q(\core.registers[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19127_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01369_),
    .Q(\core.registers[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19128_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01370_),
    .Q(\core.registers[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19129_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01371_),
    .Q(\core.registers[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19130_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_01372_),
    .Q(\core.registers[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19131_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01373_),
    .Q(\core.registers[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19132_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01374_),
    .Q(\core.registers[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19133_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01375_),
    .Q(\core.registers[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19134_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_01376_),
    .Q(\core.registers[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19135_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01377_),
    .Q(\core.registers[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19136_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01378_),
    .Q(\core.registers[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19137_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01379_),
    .Q(\core.registers[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19138_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01380_),
    .Q(\core.registers[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19139_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01381_),
    .Q(\core.registers[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19140_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01382_),
    .Q(\core.registers[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19141_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01383_),
    .Q(\core.registers[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19142_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_01384_),
    .Q(\core.registers[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19143_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_01385_),
    .Q(\core.registers[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19144_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01386_),
    .Q(\core.registers[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19145_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_01387_),
    .Q(\core.registers[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19146_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01388_),
    .Q(\core.registers[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19147_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01389_),
    .Q(\core.registers[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19148_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_01390_),
    .Q(\core.registers[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19149_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01391_),
    .Q(\core.registers[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19150_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_01392_),
    .Q(\core.registers[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19151_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01393_),
    .Q(\core.registers[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19152_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_01394_),
    .Q(\core.registers[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19153_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_01395_),
    .Q(\core.registers[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19154_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_01396_),
    .Q(\core.registers[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19155_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_01397_),
    .Q(\core.registers[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19156_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01398_),
    .Q(\core.registers[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19157_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_01399_),
    .Q(\core.registers[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19158_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01400_),
    .Q(\core.registers[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19159_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01401_),
    .Q(\core.registers[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19160_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01402_),
    .Q(\core.registers[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19161_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01403_),
    .Q(\core.registers[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19162_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_01404_),
    .Q(\core.registers[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19163_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_01405_),
    .Q(\core.registers[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19164_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01406_),
    .Q(\core.registers[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19165_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_01407_),
    .Q(\core.registers[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19166_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01408_),
    .Q(\core.registers[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19167_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01409_),
    .Q(\core.registers[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19168_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01410_),
    .Q(\core.registers[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19169_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01411_),
    .Q(\core.registers[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19170_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01412_),
    .Q(\core.registers[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19171_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01413_),
    .Q(\core.registers[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19172_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01414_),
    .Q(\core.registers[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19173_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01415_),
    .Q(\core.registers[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19174_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01416_),
    .Q(\core.registers[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19175_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01417_),
    .Q(\core.registers[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19176_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01418_),
    .Q(\core.registers[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19177_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01419_),
    .Q(\core.registers[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19178_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01420_),
    .Q(\core.registers[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19179_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01421_),
    .Q(\core.registers[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19180_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01422_),
    .Q(\core.registers[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19181_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01423_),
    .Q(\core.registers[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19182_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01424_),
    .Q(\core.registers[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19183_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01425_),
    .Q(\core.registers[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19184_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_01426_),
    .Q(\core.registers[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19185_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01427_),
    .Q(\core.registers[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19186_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01428_),
    .Q(\core.registers[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19187_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01429_),
    .Q(\core.registers[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19188_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_01430_),
    .Q(\core.registers[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19189_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_01431_),
    .Q(\core.registers[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19190_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01432_),
    .Q(\core.registers[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19191_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01433_),
    .Q(\core.registers[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19192_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01434_),
    .Q(\core.registers[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19193_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_01435_),
    .Q(\core.registers[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19194_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_01436_),
    .Q(\core.registers[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19195_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01437_),
    .Q(\core.registers[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19196_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01438_),
    .Q(\core.registers[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19197_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_01439_),
    .Q(\core.registers[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19198_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01440_),
    .Q(\core.registers[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19199_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01441_),
    .Q(\core.registers[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19200_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01442_),
    .Q(\core.registers[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19201_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01443_),
    .Q(\core.registers[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19202_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01444_),
    .Q(\core.registers[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19203_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01445_),
    .Q(\core.registers[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19204_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01446_),
    .Q(\core.registers[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19205_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01447_),
    .Q(\core.registers[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19206_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01448_),
    .Q(\core.registers[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19207_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01449_),
    .Q(\core.registers[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19208_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01450_),
    .Q(\core.registers[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19209_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_01451_),
    .Q(\core.registers[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19210_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01452_),
    .Q(\core.registers[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19211_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01453_),
    .Q(\core.registers[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19212_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01454_),
    .Q(\core.registers[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19213_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01455_),
    .Q(\core.registers[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19214_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01456_),
    .Q(\core.registers[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19215_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_01457_),
    .Q(\core.registers[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19216_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_01458_),
    .Q(\core.registers[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19217_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01459_),
    .Q(\core.registers[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19218_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01460_),
    .Q(\core.registers[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19219_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01461_),
    .Q(\core.registers[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19220_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_01462_),
    .Q(\core.registers[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19221_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_01463_),
    .Q(\core.registers[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19222_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01464_),
    .Q(\core.registers[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19223_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01465_),
    .Q(\core.registers[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19224_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01466_),
    .Q(\core.registers[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19225_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_01467_),
    .Q(\core.registers[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19226_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_01468_),
    .Q(\core.registers[30][31] ));
 sky130_fd_sc_hd__dfxtp_4 _19227_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_01469_),
    .Q(\wbSRAMInterface.currentByteSelect[0] ));
 sky130_fd_sc_hd__dfxtp_4 _19228_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_01470_),
    .Q(\wbSRAMInterface.currentByteSelect[1] ));
 sky130_fd_sc_hd__dfxtp_4 _19229_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_01471_),
    .Q(\wbSRAMInterface.currentByteSelect[2] ));
 sky130_fd_sc_hd__dfxtp_4 _19230_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_01472_),
    .Q(\wbSRAMInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__dfxtp_4 _19231_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_01473_),
    .Q(net482));
 sky130_fd_sc_hd__dfxtp_2 _19232_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01474_),
    .Q(\core.csr.instretTimer.currentValue[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19233_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01475_),
    .Q(\core.csr.instretTimer.currentValue[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19234_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01476_),
    .Q(\core.csr.instretTimer.currentValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19235_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01477_),
    .Q(\core.csr.instretTimer.currentValue[3] ));
 sky130_fd_sc_hd__dfxtp_2 _19236_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_01478_),
    .Q(\core.csr.instretTimer.currentValue[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19237_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_01479_),
    .Q(\core.csr.instretTimer.currentValue[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19238_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_01480_),
    .Q(\core.csr.instretTimer.currentValue[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19239_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_01481_),
    .Q(\core.csr.instretTimer.currentValue[7] ));
 sky130_fd_sc_hd__dfxtp_2 _19240_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_01482_),
    .Q(\core.csr.instretTimer.currentValue[8] ));
 sky130_fd_sc_hd__dfxtp_2 _19241_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01483_),
    .Q(\core.csr.instretTimer.currentValue[9] ));
 sky130_fd_sc_hd__dfxtp_2 _19242_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01484_),
    .Q(\core.csr.instretTimer.currentValue[10] ));
 sky130_fd_sc_hd__dfxtp_2 _19243_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01485_),
    .Q(\core.csr.instretTimer.currentValue[11] ));
 sky130_fd_sc_hd__dfxtp_2 _19244_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01486_),
    .Q(\core.csr.instretTimer.currentValue[12] ));
 sky130_fd_sc_hd__dfxtp_2 _19245_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01487_),
    .Q(\core.csr.instretTimer.currentValue[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19246_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01488_),
    .Q(\core.csr.instretTimer.currentValue[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19247_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01489_),
    .Q(\core.csr.instretTimer.currentValue[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19248_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01490_),
    .Q(\core.csr.instretTimer.currentValue[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19249_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01491_),
    .Q(\core.csr.instretTimer.currentValue[17] ));
 sky130_fd_sc_hd__dfxtp_2 _19250_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01492_),
    .Q(\core.csr.instretTimer.currentValue[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19251_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01493_),
    .Q(\core.csr.instretTimer.currentValue[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19252_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01494_),
    .Q(\core.csr.instretTimer.currentValue[20] ));
 sky130_fd_sc_hd__dfxtp_2 _19253_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01495_),
    .Q(\core.csr.instretTimer.currentValue[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19254_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01496_),
    .Q(\core.csr.instretTimer.currentValue[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19255_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01497_),
    .Q(\core.csr.instretTimer.currentValue[23] ));
 sky130_fd_sc_hd__dfxtp_2 _19256_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01498_),
    .Q(\core.csr.instretTimer.currentValue[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19257_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01499_),
    .Q(\core.csr.instretTimer.currentValue[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19258_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01500_),
    .Q(\core.csr.instretTimer.currentValue[26] ));
 sky130_fd_sc_hd__dfxtp_2 _19259_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01501_),
    .Q(\core.csr.instretTimer.currentValue[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19260_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01502_),
    .Q(\core.csr.instretTimer.currentValue[28] ));
 sky130_fd_sc_hd__dfxtp_2 _19261_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01503_),
    .Q(\core.csr.instretTimer.currentValue[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19262_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01504_),
    .Q(\core.csr.instretTimer.currentValue[30] ));
 sky130_fd_sc_hd__dfxtp_2 _19263_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01505_),
    .Q(\core.csr.instretTimer.currentValue[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19264_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01506_),
    .Q(\core.csr.instretTimer.currentValue[32] ));
 sky130_fd_sc_hd__dfxtp_1 _19265_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01507_),
    .Q(\core.csr.instretTimer.currentValue[33] ));
 sky130_fd_sc_hd__dfxtp_1 _19266_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01508_),
    .Q(\core.csr.instretTimer.currentValue[34] ));
 sky130_fd_sc_hd__dfxtp_1 _19267_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01509_),
    .Q(\core.csr.instretTimer.currentValue[35] ));
 sky130_fd_sc_hd__dfxtp_1 _19268_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01510_),
    .Q(\core.csr.instretTimer.currentValue[36] ));
 sky130_fd_sc_hd__dfxtp_1 _19269_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_01511_),
    .Q(\core.csr.instretTimer.currentValue[37] ));
 sky130_fd_sc_hd__dfxtp_1 _19270_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_01512_),
    .Q(\core.csr.instretTimer.currentValue[38] ));
 sky130_fd_sc_hd__dfxtp_1 _19271_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_01513_),
    .Q(\core.csr.instretTimer.currentValue[39] ));
 sky130_fd_sc_hd__dfxtp_1 _19272_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_01514_),
    .Q(\core.csr.instretTimer.currentValue[40] ));
 sky130_fd_sc_hd__dfxtp_1 _19273_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_01515_),
    .Q(\core.csr.instretTimer.currentValue[41] ));
 sky130_fd_sc_hd__dfxtp_1 _19274_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01516_),
    .Q(\core.csr.instretTimer.currentValue[42] ));
 sky130_fd_sc_hd__dfxtp_1 _19275_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01517_),
    .Q(\core.csr.instretTimer.currentValue[43] ));
 sky130_fd_sc_hd__dfxtp_1 _19276_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01518_),
    .Q(\core.csr.instretTimer.currentValue[44] ));
 sky130_fd_sc_hd__dfxtp_1 _19277_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01519_),
    .Q(\core.csr.instretTimer.currentValue[45] ));
 sky130_fd_sc_hd__dfxtp_1 _19278_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01520_),
    .Q(\core.csr.instretTimer.currentValue[46] ));
 sky130_fd_sc_hd__dfxtp_1 _19279_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01521_),
    .Q(\core.csr.instretTimer.currentValue[47] ));
 sky130_fd_sc_hd__dfxtp_1 _19280_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01522_),
    .Q(\core.csr.instretTimer.currentValue[48] ));
 sky130_fd_sc_hd__dfxtp_1 _19281_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01523_),
    .Q(\core.csr.instretTimer.currentValue[49] ));
 sky130_fd_sc_hd__dfxtp_1 _19282_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01524_),
    .Q(\core.csr.instretTimer.currentValue[50] ));
 sky130_fd_sc_hd__dfxtp_1 _19283_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01525_),
    .Q(\core.csr.instretTimer.currentValue[51] ));
 sky130_fd_sc_hd__dfxtp_1 _19284_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01526_),
    .Q(\core.csr.instretTimer.currentValue[52] ));
 sky130_fd_sc_hd__dfxtp_1 _19285_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01527_),
    .Q(\core.csr.instretTimer.currentValue[53] ));
 sky130_fd_sc_hd__dfxtp_1 _19286_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_01528_),
    .Q(\core.csr.instretTimer.currentValue[54] ));
 sky130_fd_sc_hd__dfxtp_1 _19287_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01529_),
    .Q(\core.csr.instretTimer.currentValue[55] ));
 sky130_fd_sc_hd__dfxtp_1 _19288_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01530_),
    .Q(\core.csr.instretTimer.currentValue[56] ));
 sky130_fd_sc_hd__dfxtp_1 _19289_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01531_),
    .Q(\core.csr.instretTimer.currentValue[57] ));
 sky130_fd_sc_hd__dfxtp_1 _19290_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01532_),
    .Q(\core.csr.instretTimer.currentValue[58] ));
 sky130_fd_sc_hd__dfxtp_1 _19291_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01533_),
    .Q(\core.csr.instretTimer.currentValue[59] ));
 sky130_fd_sc_hd__dfxtp_1 _19292_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01534_),
    .Q(\core.csr.instretTimer.currentValue[60] ));
 sky130_fd_sc_hd__dfxtp_2 _19293_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01535_),
    .Q(\core.csr.instretTimer.currentValue[61] ));
 sky130_fd_sc_hd__dfxtp_1 _19294_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01536_),
    .Q(\core.csr.instretTimer.currentValue[62] ));
 sky130_fd_sc_hd__dfxtp_1 _19295_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01537_),
    .Q(\core.csr.instretTimer.currentValue[63] ));
 sky130_fd_sc_hd__dfxtp_1 _19296_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_01538_),
    .Q(\core.csr.mconfigptr.currentValue[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19297_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_01539_),
    .Q(\core.csr.mconfigptr.currentValue[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19298_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_01540_),
    .Q(\core.csr.mconfigptr.currentValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19299_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_01541_),
    .Q(\core.csr.mconfigptr.currentValue[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19300_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_01542_),
    .Q(\core.csr.mconfigptr.currentValue[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19301_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_01543_),
    .Q(\core.csr.mconfigptr.currentValue[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19302_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01544_),
    .Q(\core.csr.mconfigptr.currentValue[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19303_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_01545_),
    .Q(\core.csr.mconfigptr.currentValue[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19304_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_01546_),
    .Q(\core.csr.mconfigptr.currentValue[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19305_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01547_),
    .Q(\core.csr.mconfigptr.currentValue[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19306_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01548_),
    .Q(\core.csr.mconfigptr.currentValue[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19307_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_01549_),
    .Q(\core.csr.mconfigptr.currentValue[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19308_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_01550_),
    .Q(\core.csr.mconfigptr.currentValue[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19309_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_01551_),
    .Q(\core.csr.mconfigptr.currentValue[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19310_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_01552_),
    .Q(\core.csr.mconfigptr.currentValue[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19311_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_01553_),
    .Q(\core.csr.mconfigptr.currentValue[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19312_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01554_),
    .Q(\core.csr.mconfigptr.currentValue[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19313_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01555_),
    .Q(\core.csr.mconfigptr.currentValue[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19314_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_01556_),
    .Q(\core.csr.mconfigptr.currentValue[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19315_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01557_),
    .Q(\core.csr.mconfigptr.currentValue[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19316_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01558_),
    .Q(\core.csr.mconfigptr.currentValue[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19317_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01559_),
    .Q(\core.csr.mconfigptr.currentValue[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19318_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_01560_),
    .Q(\core.csr.mconfigptr.currentValue[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19319_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_01561_),
    .Q(\core.csr.mconfigptr.currentValue[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19320_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_01562_),
    .Q(\core.csr.mconfigptr.currentValue[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19321_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_01563_),
    .Q(\core.csr.mconfigptr.currentValue[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19322_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_01564_),
    .Q(\core.csr.mconfigptr.currentValue[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19323_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_01565_),
    .Q(\core.csr.mconfigptr.currentValue[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19324_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_01566_),
    .Q(\core.csr.mconfigptr.currentValue[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19325_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01567_),
    .Q(\core.csr.mconfigptr.currentValue[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19326_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_01568_),
    .Q(\core.csr.mconfigptr.currentValue[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19327_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01569_),
    .Q(\core.csr.mconfigptr.currentValue[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19328_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01570_),
    .Q(\core.csr.traps.mscratch.currentValue[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19329_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01571_),
    .Q(\core.csr.traps.mscratch.currentValue[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19330_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01572_),
    .Q(\core.csr.traps.mscratch.currentValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19331_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01573_),
    .Q(\core.csr.traps.mscratch.currentValue[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19332_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01574_),
    .Q(\core.csr.traps.mscratch.currentValue[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19333_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01575_),
    .Q(\core.csr.traps.mscratch.currentValue[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19334_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01576_),
    .Q(\core.csr.traps.mscratch.currentValue[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19335_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01577_),
    .Q(\core.csr.traps.mscratch.currentValue[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19336_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01578_),
    .Q(\core.csr.traps.mscratch.currentValue[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19337_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_01579_),
    .Q(\core.csr.traps.mscratch.currentValue[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19338_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01580_),
    .Q(\core.csr.traps.mscratch.currentValue[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19339_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01581_),
    .Q(\core.csr.traps.mscratch.currentValue[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19340_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01582_),
    .Q(\core.csr.traps.mscratch.currentValue[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19341_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01583_),
    .Q(\core.csr.traps.mscratch.currentValue[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19342_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01584_),
    .Q(\core.csr.traps.mscratch.currentValue[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19343_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_01585_),
    .Q(\core.csr.traps.mscratch.currentValue[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19344_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01586_),
    .Q(\core.csr.traps.mscratch.currentValue[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19345_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_01587_),
    .Q(\core.csr.traps.mscratch.currentValue[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19346_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01588_),
    .Q(\core.csr.traps.mscratch.currentValue[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19347_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01589_),
    .Q(\core.csr.traps.mscratch.currentValue[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19348_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01590_),
    .Q(\core.csr.traps.mscratch.currentValue[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19349_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_01591_),
    .Q(\core.csr.traps.mscratch.currentValue[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19350_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01592_),
    .Q(\core.csr.traps.mscratch.currentValue[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19351_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01593_),
    .Q(\core.csr.traps.mscratch.currentValue[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19352_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01594_),
    .Q(\core.csr.traps.mscratch.currentValue[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19353_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01595_),
    .Q(\core.csr.traps.mscratch.currentValue[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19354_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01596_),
    .Q(\core.csr.traps.mscratch.currentValue[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19355_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01597_),
    .Q(\core.csr.traps.mscratch.currentValue[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19356_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01598_),
    .Q(\core.csr.traps.mscratch.currentValue[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19357_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01599_),
    .Q(\core.csr.traps.mscratch.currentValue[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19358_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01600_),
    .Q(\core.csr.traps.mscratch.currentValue[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19359_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01601_),
    .Q(\core.csr.traps.mscratch.currentValue[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19360_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01602_),
    .Q(\core.csr.traps.mie.currentValue[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19361_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01603_),
    .Q(\core.csr.traps.mie.currentValue[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19362_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01604_),
    .Q(\core.csr.traps.mie.currentValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19363_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01605_),
    .Q(\core.csr.traps.mie.currentValue[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19364_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01606_),
    .Q(\core.csr.traps.mie.currentValue[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19365_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01607_),
    .Q(\core.csr.traps.mie.currentValue[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19366_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01608_),
    .Q(\core.csr.traps.mie.currentValue[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19367_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01609_),
    .Q(\core.csr.traps.mie.currentValue[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19368_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01610_),
    .Q(\core.csr.traps.mie.currentValue[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19369_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_01611_),
    .Q(\core.csr.traps.mie.currentValue[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19370_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01612_),
    .Q(\core.csr.traps.mie.currentValue[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19371_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01613_),
    .Q(\core.csr.traps.mie.currentValue[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19372_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01614_),
    .Q(\core.csr.traps.mie.currentValue[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19373_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01615_),
    .Q(\core.csr.traps.mie.currentValue[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19374_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01616_),
    .Q(\core.csr.traps.mie.currentValue[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19375_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_01617_),
    .Q(\core.csr.traps.mie.currentValue[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19376_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01618_),
    .Q(\core.csr.traps.mie.currentValue[16] ));
 sky130_fd_sc_hd__dfxtp_2 _19377_ (.CLK(clknet_leaf_161_wb_clk_i),
    .D(_01619_),
    .Q(\core.csr.traps.mie.currentValue[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19378_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01620_),
    .Q(\core.csr.traps.mie.currentValue[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19379_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01621_),
    .Q(\core.csr.traps.mie.currentValue[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19380_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01622_),
    .Q(\core.csr.traps.mie.currentValue[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19381_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_01623_),
    .Q(\core.csr.traps.mie.currentValue[21] ));
 sky130_fd_sc_hd__dfxtp_2 _19382_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01624_),
    .Q(\core.csr.traps.mie.currentValue[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19383_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01625_),
    .Q(\core.csr.traps.mie.currentValue[23] ));
 sky130_fd_sc_hd__dfxtp_2 _19384_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01626_),
    .Q(\core.csr.traps.mie.currentValue[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19385_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01627_),
    .Q(\core.csr.traps.mie.currentValue[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19386_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01628_),
    .Q(\core.csr.traps.mie.currentValue[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19387_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01629_),
    .Q(\core.csr.traps.mie.currentValue[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19388_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01630_),
    .Q(\core.csr.traps.mie.currentValue[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19389_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01631_),
    .Q(\core.csr.traps.mie.currentValue[29] ));
 sky130_fd_sc_hd__dfxtp_2 _19390_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01632_),
    .Q(\core.csr.traps.mie.currentValue[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19391_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01633_),
    .Q(\core.csr.traps.mie.currentValue[31] ));
 sky130_fd_sc_hd__dfxtp_2 _19392_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01634_),
    .Q(\core.csr.traps.mcause.csrReadData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19393_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01635_),
    .Q(\core.csr.traps.mcause.csrReadData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19394_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01636_),
    .Q(\core.csr.traps.mcause.csrReadData[2] ));
 sky130_fd_sc_hd__dfxtp_4 _19395_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01637_),
    .Q(\core.csr.traps.mcause.csrReadData[3] ));
 sky130_fd_sc_hd__dfxtp_2 _19396_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01638_),
    .Q(\core.csr.traps.mcause.csrReadData[4] ));
 sky130_fd_sc_hd__dfxtp_2 _19397_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01639_),
    .Q(\core.csr.traps.mcause.csrReadData[5] ));
 sky130_fd_sc_hd__dfxtp_2 _19398_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01640_),
    .Q(\core.csr.traps.mcause.csrReadData[6] ));
 sky130_fd_sc_hd__dfxtp_2 _19399_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01641_),
    .Q(\core.csr.traps.mcause.csrReadData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19400_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_01642_),
    .Q(\core.csr.traps.mcause.csrReadData[8] ));
 sky130_fd_sc_hd__dfxtp_4 _19401_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_01643_),
    .Q(\core.csr.traps.mcause.csrReadData[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19402_ (.CLK(clknet_leaf_151_wb_clk_i),
    .D(_01644_),
    .Q(\core.csr.traps.mcause.csrReadData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19403_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01645_),
    .Q(\core.csr.traps.mcause.csrReadData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19404_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01646_),
    .Q(\core.csr.traps.mcause.csrReadData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19405_ (.CLK(clknet_leaf_151_wb_clk_i),
    .D(_01647_),
    .Q(\core.csr.traps.mcause.csrReadData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19406_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01648_),
    .Q(\core.csr.traps.mcause.csrReadData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19407_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01649_),
    .Q(\core.csr.traps.mcause.csrReadData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19408_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01650_),
    .Q(\core.csr.traps.mcause.csrReadData[16] ));
 sky130_fd_sc_hd__dfxtp_2 _19409_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_01651_),
    .Q(\core.csr.traps.mcause.csrReadData[17] ));
 sky130_fd_sc_hd__dfxtp_2 _19410_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01652_),
    .Q(\core.csr.traps.mcause.csrReadData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19411_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01653_),
    .Q(\core.csr.traps.mcause.csrReadData[19] ));
 sky130_fd_sc_hd__dfxtp_2 _19412_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01654_),
    .Q(\core.csr.traps.mcause.csrReadData[20] ));
 sky130_fd_sc_hd__dfxtp_2 _19413_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_01655_),
    .Q(\core.csr.traps.mcause.csrReadData[21] ));
 sky130_fd_sc_hd__dfxtp_2 _19414_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01656_),
    .Q(\core.csr.traps.mcause.csrReadData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19415_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01657_),
    .Q(\core.csr.traps.mcause.csrReadData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19416_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01658_),
    .Q(\core.csr.traps.mcause.csrReadData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19417_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01659_),
    .Q(\core.csr.traps.mcause.csrReadData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19418_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01660_),
    .Q(\core.csr.traps.mcause.csrReadData[26] ));
 sky130_fd_sc_hd__dfxtp_2 _19419_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01661_),
    .Q(\core.csr.traps.mcause.csrReadData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19420_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01662_),
    .Q(\core.csr.traps.mcause.csrReadData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19421_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_01663_),
    .Q(\core.csr.traps.mcause.csrReadData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19422_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_01664_),
    .Q(\core.csr.traps.mcause.csrReadData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19423_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01665_),
    .Q(\core.csr.traps.mcause.csrReadData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19424_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01666_),
    .Q(\core.csr.trapReturnVector[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19425_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01667_),
    .Q(\core.csr.trapReturnVector[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19426_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_01668_),
    .Q(\core.csr.trapReturnVector[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19427_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_01669_),
    .Q(\core.csr.trapReturnVector[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19428_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_01670_),
    .Q(\core.csr.trapReturnVector[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19429_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01671_),
    .Q(\core.csr.trapReturnVector[5] ));
 sky130_fd_sc_hd__dfxtp_2 _19430_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01672_),
    .Q(\core.csr.trapReturnVector[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19431_ (.CLK(clknet_leaf_151_wb_clk_i),
    .D(_01673_),
    .Q(\core.csr.trapReturnVector[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19432_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_01674_),
    .Q(\core.csr.trapReturnVector[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19433_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_01675_),
    .Q(\core.csr.trapReturnVector[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19434_ (.CLK(clknet_leaf_151_wb_clk_i),
    .D(_01676_),
    .Q(\core.csr.trapReturnVector[10] ));
 sky130_fd_sc_hd__dfxtp_2 _19435_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01677_),
    .Q(\core.csr.trapReturnVector[11] ));
 sky130_fd_sc_hd__dfxtp_2 _19436_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01678_),
    .Q(\core.csr.trapReturnVector[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19437_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01679_),
    .Q(\core.csr.trapReturnVector[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19438_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_01680_),
    .Q(\core.csr.trapReturnVector[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19439_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01681_),
    .Q(\core.csr.trapReturnVector[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19440_ (.CLK(clknet_leaf_161_wb_clk_i),
    .D(_01682_),
    .Q(\core.csr.trapReturnVector[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19441_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_01683_),
    .Q(\core.csr.trapReturnVector[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19442_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01684_),
    .Q(\core.csr.trapReturnVector[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19443_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_01685_),
    .Q(\core.csr.trapReturnVector[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19444_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_01686_),
    .Q(\core.csr.trapReturnVector[20] ));
 sky130_fd_sc_hd__dfxtp_2 _19445_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_01687_),
    .Q(\core.csr.trapReturnVector[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19446_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01688_),
    .Q(\core.csr.trapReturnVector[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19447_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01689_),
    .Q(\core.csr.trapReturnVector[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19448_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01690_),
    .Q(\core.csr.trapReturnVector[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19449_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01691_),
    .Q(\core.csr.trapReturnVector[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19450_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_01692_),
    .Q(\core.csr.trapReturnVector[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19451_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01693_),
    .Q(\core.csr.trapReturnVector[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19452_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_01694_),
    .Q(\core.csr.trapReturnVector[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19453_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_01695_),
    .Q(\core.csr.trapReturnVector[29] ));
 sky130_fd_sc_hd__dfxtp_4 _19454_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_01696_),
    .Q(\core.csr.trapReturnVector[30] ));
 sky130_fd_sc_hd__dfxtp_2 _19455_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_01697_),
    .Q(\core.csr.trapReturnVector[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19456_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01698_),
    .Q(\core.csr.traps.mtvec.csrReadData[0] ));
 sky130_fd_sc_hd__dfxtp_2 _19457_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01699_),
    .Q(\core.csr.traps.mtvec.csrReadData[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19458_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01700_),
    .Q(\core.csr.traps.mtvec.csrReadData[2] ));
 sky130_fd_sc_hd__dfxtp_2 _19459_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01701_),
    .Q(\core.csr.traps.mtvec.csrReadData[3] ));
 sky130_fd_sc_hd__dfxtp_2 _19460_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01702_),
    .Q(\core.csr.traps.mtvec.csrReadData[4] ));
 sky130_fd_sc_hd__dfxtp_4 _19461_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01703_),
    .Q(\core.csr.traps.mtvec.csrReadData[5] ));
 sky130_fd_sc_hd__dfxtp_2 _19462_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01704_),
    .Q(\core.csr.traps.mtvec.csrReadData[6] ));
 sky130_fd_sc_hd__dfxtp_4 _19463_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01705_),
    .Q(\core.csr.traps.mtvec.csrReadData[7] ));
 sky130_fd_sc_hd__dfxtp_2 _19464_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01706_),
    .Q(\core.csr.traps.mtvec.csrReadData[8] ));
 sky130_fd_sc_hd__dfxtp_2 _19465_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_01707_),
    .Q(\core.csr.traps.mtvec.csrReadData[9] ));
 sky130_fd_sc_hd__dfxtp_2 _19466_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01708_),
    .Q(\core.csr.traps.mtvec.csrReadData[10] ));
 sky130_fd_sc_hd__dfxtp_4 _19467_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01709_),
    .Q(\core.csr.traps.mtvec.csrReadData[11] ));
 sky130_fd_sc_hd__dfxtp_2 _19468_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01710_),
    .Q(\core.csr.traps.mtvec.csrReadData[12] ));
 sky130_fd_sc_hd__dfxtp_2 _19469_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01711_),
    .Q(\core.csr.traps.mtvec.csrReadData[13] ));
 sky130_fd_sc_hd__dfxtp_2 _19470_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01712_),
    .Q(\core.csr.traps.mtvec.csrReadData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19471_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_01713_),
    .Q(\core.csr.traps.mtvec.csrReadData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19472_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01714_),
    .Q(\core.csr.traps.mtvec.csrReadData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19473_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_01715_),
    .Q(\core.csr.traps.mtvec.csrReadData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19474_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01716_),
    .Q(\core.csr.traps.mtvec.csrReadData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19475_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01717_),
    .Q(\core.csr.traps.mtvec.csrReadData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19476_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01718_),
    .Q(\core.csr.traps.mtvec.csrReadData[20] ));
 sky130_fd_sc_hd__dfxtp_4 _19477_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_01719_),
    .Q(\core.csr.traps.mtvec.csrReadData[21] ));
 sky130_fd_sc_hd__dfxtp_2 _19478_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01720_),
    .Q(\core.csr.traps.mtvec.csrReadData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19479_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01721_),
    .Q(\core.csr.traps.mtvec.csrReadData[23] ));
 sky130_fd_sc_hd__dfxtp_2 _19480_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01722_),
    .Q(\core.csr.traps.mtvec.csrReadData[24] ));
 sky130_fd_sc_hd__dfxtp_2 _19481_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01723_),
    .Q(\core.csr.traps.mtvec.csrReadData[25] ));
 sky130_fd_sc_hd__dfxtp_2 _19482_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01724_),
    .Q(\core.csr.traps.mtvec.csrReadData[26] ));
 sky130_fd_sc_hd__dfxtp_2 _19483_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01725_),
    .Q(\core.csr.traps.mtvec.csrReadData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19484_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01726_),
    .Q(\core.csr.traps.mtvec.csrReadData[28] ));
 sky130_fd_sc_hd__dfxtp_2 _19485_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01727_),
    .Q(\core.csr.traps.mtvec.csrReadData[29] ));
 sky130_fd_sc_hd__dfxtp_4 _19486_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01728_),
    .Q(\core.csr.traps.mtvec.csrReadData[30] ));
 sky130_fd_sc_hd__dfxtp_2 _19487_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01729_),
    .Q(\core.csr.traps.mtvec.csrReadData[31] ));
 sky130_fd_sc_hd__dfxtp_4 _19488_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01730_),
    .Q(\core.csr.traps.machineInterruptEnable ));
 sky130_fd_sc_hd__dfxtp_2 _19489_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01731_),
    .Q(\core.csr.traps.machinePreviousInterruptEnable ));
 sky130_fd_sc_hd__dfxtp_1 _19490_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_01732_),
    .Q(\core.csr.traps.mtval.csrReadData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19491_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01733_),
    .Q(\core.csr.traps.mtval.csrReadData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19492_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_01734_),
    .Q(\core.csr.traps.mtval.csrReadData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19493_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_01735_),
    .Q(\core.csr.traps.mtval.csrReadData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19494_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01736_),
    .Q(\core.csr.traps.mtval.csrReadData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19495_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01737_),
    .Q(\core.csr.traps.mtval.csrReadData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19496_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01738_),
    .Q(\core.csr.traps.mtval.csrReadData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19497_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01739_),
    .Q(\core.csr.traps.mtval.csrReadData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19498_ (.CLK(clknet_leaf_151_wb_clk_i),
    .D(_01740_),
    .Q(\core.csr.traps.mtval.csrReadData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19499_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_01741_),
    .Q(\core.csr.traps.mtval.csrReadData[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19500_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01742_),
    .Q(\core.csr.traps.mtval.csrReadData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19501_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01743_),
    .Q(\core.csr.traps.mtval.csrReadData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19502_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01744_),
    .Q(\core.csr.traps.mtval.csrReadData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19503_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_01745_),
    .Q(\core.csr.traps.mtval.csrReadData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19504_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_01746_),
    .Q(\core.csr.traps.mtval.csrReadData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19505_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01747_),
    .Q(\core.csr.traps.mtval.csrReadData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19506_ (.CLK(clknet_leaf_161_wb_clk_i),
    .D(_01748_),
    .Q(\core.csr.traps.mtval.csrReadData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19507_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_01749_),
    .Q(\core.csr.traps.mtval.csrReadData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19508_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_01750_),
    .Q(\core.csr.traps.mtval.csrReadData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19509_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_01751_),
    .Q(\core.csr.traps.mtval.csrReadData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19510_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01752_),
    .Q(\core.csr.traps.mtval.csrReadData[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19511_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_01753_),
    .Q(\core.csr.traps.mtval.csrReadData[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19512_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01754_),
    .Q(\core.csr.traps.mtval.csrReadData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19513_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01755_),
    .Q(\core.csr.traps.mtval.csrReadData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19514_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01756_),
    .Q(\core.csr.traps.mtval.csrReadData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19515_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01757_),
    .Q(\core.csr.traps.mtval.csrReadData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19516_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_01758_),
    .Q(\core.csr.traps.mtval.csrReadData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19517_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01759_),
    .Q(\core.csr.traps.mtval.csrReadData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19518_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01760_),
    .Q(\core.csr.traps.mtval.csrReadData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19519_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01761_),
    .Q(\core.csr.traps.mtval.csrReadData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19520_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_01762_),
    .Q(\core.csr.traps.mtval.csrReadData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19521_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_01763_),
    .Q(\core.csr.traps.mtval.csrReadData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19522_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01764_),
    .Q(\core.csr.traps.mip.csrReadData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19523_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01765_),
    .Q(\core.csr.traps.mip.csrReadData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19524_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01766_),
    .Q(\core.csr.traps.mip.csrReadData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19525_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01767_),
    .Q(\core.csr.traps.mip.csrReadData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19526_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_01768_),
    .Q(\core.csr.traps.mip.csrReadData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19527_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01769_),
    .Q(\core.csr.traps.mip.csrReadData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19528_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01770_),
    .Q(\core.csr.traps.mip.csrReadData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19529_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01771_),
    .Q(\core.csr.traps.mip.csrReadData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19530_ (.CLK(clknet_leaf_151_wb_clk_i),
    .D(_01772_),
    .Q(\core.csr.traps.mip.csrReadData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19531_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_01773_),
    .Q(\core.csr.traps.mip.csrReadData[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19532_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01774_),
    .Q(\core.csr.traps.mip.csrReadData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19533_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01775_),
    .Q(\core.csr.traps.mip.csrReadData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19534_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01776_),
    .Q(\core.csr.traps.mip.csrReadData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19535_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_01777_),
    .Q(\core.csr.traps.mip.csrReadData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19536_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_01778_),
    .Q(\core.csr.traps.mip.csrReadData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19537_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01779_),
    .Q(\core.csr.traps.mip.csrReadData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19538_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01780_),
    .Q(\core.csr.traps.mip.csrReadData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19539_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01781_),
    .Q(\core.csr.traps.mip.csrReadData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19540_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01782_),
    .Q(\core.csr.traps.mip.csrReadData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19541_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01783_),
    .Q(\core.csr.traps.mip.csrReadData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19542_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01784_),
    .Q(\core.csr.traps.mip.csrReadData[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19543_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01785_),
    .Q(\core.csr.traps.mip.csrReadData[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19544_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01786_),
    .Q(\core.csr.traps.mip.csrReadData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19545_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01787_),
    .Q(\core.csr.traps.mip.csrReadData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19546_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01788_),
    .Q(\core.csr.traps.mip.csrReadData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19547_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01789_),
    .Q(\core.csr.traps.mip.csrReadData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19548_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01790_),
    .Q(\core.csr.traps.mip.csrReadData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19549_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01791_),
    .Q(\core.csr.traps.mip.csrReadData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19550_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01792_),
    .Q(\core.csr.traps.mip.csrReadData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19551_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01793_),
    .Q(\core.csr.traps.mip.csrReadData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19552_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_01794_),
    .Q(\core.csr.traps.mip.csrReadData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19553_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01795_),
    .Q(\core.csr.traps.mip.csrReadData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19554_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_01796_),
    .Q(\core.registers[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19555_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01797_),
    .Q(\core.registers[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19556_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01798_),
    .Q(\core.registers[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19557_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01799_),
    .Q(\core.registers[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19558_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01800_),
    .Q(\core.registers[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19559_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01801_),
    .Q(\core.registers[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19560_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01802_),
    .Q(\core.registers[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19561_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01803_),
    .Q(\core.registers[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19562_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01804_),
    .Q(\core.registers[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19563_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01805_),
    .Q(\core.registers[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19564_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01806_),
    .Q(\core.registers[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19565_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01807_),
    .Q(\core.registers[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19566_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01808_),
    .Q(\core.registers[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19567_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01809_),
    .Q(\core.registers[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19568_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_01810_),
    .Q(\core.registers[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19569_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01811_),
    .Q(\core.registers[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19570_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_01812_),
    .Q(\core.registers[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19571_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01813_),
    .Q(\core.registers[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19572_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01814_),
    .Q(\core.registers[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19573_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_01815_),
    .Q(\core.registers[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19574_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_01816_),
    .Q(\core.registers[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19575_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_01817_),
    .Q(\core.registers[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19576_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01818_),
    .Q(\core.registers[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19577_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_01819_),
    .Q(\core.registers[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19578_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_01820_),
    .Q(\core.registers[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19579_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_01821_),
    .Q(\core.registers[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19580_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01822_),
    .Q(\core.registers[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19581_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01823_),
    .Q(\core.registers[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19582_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01824_),
    .Q(\core.registers[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19583_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01825_),
    .Q(\core.registers[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19584_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_01826_),
    .Q(\core.registers[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19585_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01827_),
    .Q(\core.registers[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19586_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_01828_),
    .Q(\core.registers[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19587_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01829_),
    .Q(\core.registers[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19588_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01830_),
    .Q(\core.registers[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19589_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01831_),
    .Q(\core.registers[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19590_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01832_),
    .Q(\core.registers[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19591_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01833_),
    .Q(\core.registers[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19592_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01834_),
    .Q(\core.registers[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19593_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01835_),
    .Q(\core.registers[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19594_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01836_),
    .Q(\core.registers[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19595_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01837_),
    .Q(\core.registers[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19596_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01838_),
    .Q(\core.registers[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19597_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01839_),
    .Q(\core.registers[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19598_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01840_),
    .Q(\core.registers[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19599_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01841_),
    .Q(\core.registers[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19600_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_01842_),
    .Q(\core.registers[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19601_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01843_),
    .Q(\core.registers[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19602_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_01844_),
    .Q(\core.registers[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19603_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01845_),
    .Q(\core.registers[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19604_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01846_),
    .Q(\core.registers[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19605_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01847_),
    .Q(\core.registers[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19606_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_01848_),
    .Q(\core.registers[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19607_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01849_),
    .Q(\core.registers[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19608_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01850_),
    .Q(\core.registers[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19609_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_01851_),
    .Q(\core.registers[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19610_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_01852_),
    .Q(\core.registers[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19611_ (.CLK(clknet_leaf_187_wb_clk_i),
    .D(_01853_),
    .Q(\core.registers[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19612_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01854_),
    .Q(\core.registers[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19613_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01855_),
    .Q(\core.registers[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19614_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01856_),
    .Q(\core.registers[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19615_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01857_),
    .Q(\core.registers[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19616_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_01858_),
    .Q(\core.registers[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19617_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01859_),
    .Q(\core.registers[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19618_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01860_),
    .Q(\core.registers[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19619_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01861_),
    .Q(\core.registers[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19620_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01862_),
    .Q(\core.registers[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19621_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01863_),
    .Q(\core.registers[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19622_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01864_),
    .Q(\core.registers[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19623_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01865_),
    .Q(\core.registers[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19624_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_01866_),
    .Q(\core.registers[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19625_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01867_),
    .Q(\core.registers[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19626_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01868_),
    .Q(\core.registers[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19627_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01869_),
    .Q(\core.registers[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19628_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01870_),
    .Q(\core.registers[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19629_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01871_),
    .Q(\core.registers[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19630_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01872_),
    .Q(\core.registers[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19631_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01873_),
    .Q(\core.registers[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19632_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01874_),
    .Q(\core.registers[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19633_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01875_),
    .Q(\core.registers[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19634_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_01876_),
    .Q(\core.registers[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19635_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01877_),
    .Q(\core.registers[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19636_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01878_),
    .Q(\core.registers[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19637_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01879_),
    .Q(\core.registers[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19638_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_01880_),
    .Q(\core.registers[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19639_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01881_),
    .Q(\core.registers[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19640_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01882_),
    .Q(\core.registers[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19641_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_01883_),
    .Q(\core.registers[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19642_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_01884_),
    .Q(\core.registers[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19643_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_01885_),
    .Q(\core.registers[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19644_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_01886_),
    .Q(\core.registers[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19645_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_01887_),
    .Q(\core.registers[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19646_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01888_),
    .Q(\core.registers[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19647_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01889_),
    .Q(\core.registers[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19648_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_01890_),
    .Q(\core.registers[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19649_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_01891_),
    .Q(\core.registers[14][31] ));
 sky130_fd_sc_hd__dfxtp_2 _19650_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_01892_),
    .Q(\core.pipe2_stall ));
 sky130_fd_sc_hd__buf_2 _19652_ (.A(clknet_4_0__leaf_wb_clk_i),
    .X(net303));
 sky130_fd_sc_hd__buf_2 _19653_ (.A(clknet_leaf_45_wb_clk_i),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_4_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_4_10__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_4_11__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_4_12__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_4_13__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_4_14__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_4_15__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_4_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_4_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_4_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_4_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_4_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_4_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_4_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_4_8__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_4_9__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_100_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_101_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_102_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_103_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_104_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_105_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_106_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_107_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_108_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_109_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_110_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_111_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_112_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_113_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_114_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_115_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_116_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_117_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_118_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_119_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_120_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_121_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_122_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_123_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_124_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_125_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_126_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_127_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_128_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_129_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_130_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_131_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_132_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_133_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_134_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_135_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_136_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_137_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_138_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_139_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_140_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_141_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_142_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_143_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_144_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_145_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_146_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_147_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_148_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_149_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_150_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_151_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_152_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_153_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_154_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_155_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_156_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_157_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_158_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_159_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_160_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_161_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_162_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_163_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_164_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_165_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_166_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_167_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_168_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_169_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_170_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_171_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_172_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_173_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_174_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_175_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_176_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_177_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_178_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_179_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_180_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_181_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_182_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_183_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_184_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_185_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_186_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_187_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_188_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_189_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_190_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_191_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_192_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_193_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_194_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_195_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_196_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_197_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_198_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_199_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_200_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_201_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_202_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_51_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_52_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_53_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_54_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_55_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_56_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_57_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_58_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_59_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_60_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_61_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_62_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_63_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_64_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_65_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_66_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_67_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_68_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_69_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_70_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_71_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_72_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_73_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_74_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_75_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_76_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_77_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_78_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_79_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_80_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_81_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_82_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_83_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_84_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_85_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_86_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_87_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_88_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_89_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_90_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_91_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_92_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_93_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_94_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_95_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_96_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_97_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_98_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_99_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_4 fanout1000 (.A(net1001),
    .X(net1000));
 sky130_fd_sc_hd__buf_2 fanout1001 (.A(net1004),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_4 fanout1002 (.A(net1004),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_2 fanout1003 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__buf_12 fanout1004 (.A(_05373_),
    .X(net1004));
 sky130_fd_sc_hd__buf_6 fanout1005 (.A(_05069_),
    .X(net1005));
 sky130_fd_sc_hd__buf_4 fanout1006 (.A(_05069_),
    .X(net1006));
 sky130_fd_sc_hd__buf_8 fanout1007 (.A(net1008),
    .X(net1007));
 sky130_fd_sc_hd__buf_12 fanout1008 (.A(_03124_),
    .X(net1008));
 sky130_fd_sc_hd__buf_12 fanout1009 (.A(net1010),
    .X(net1009));
 sky130_fd_sc_hd__buf_8 fanout1010 (.A(_03124_),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_16 fanout1011 (.A(_02215_),
    .X(net1011));
 sky130_fd_sc_hd__buf_4 fanout1012 (.A(_02215_),
    .X(net1012));
 sky130_fd_sc_hd__buf_12 fanout1013 (.A(net1014),
    .X(net1013));
 sky130_fd_sc_hd__buf_12 fanout1014 (.A(_02215_),
    .X(net1014));
 sky130_fd_sc_hd__buf_12 fanout1015 (.A(net1018),
    .X(net1015));
 sky130_fd_sc_hd__buf_12 fanout1016 (.A(net1017),
    .X(net1016));
 sky130_fd_sc_hd__buf_12 fanout1017 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__buf_12 fanout1018 (.A(_08768_),
    .X(net1018));
 sky130_fd_sc_hd__buf_4 fanout1019 (.A(net1022),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_4 fanout1020 (.A(net1022),
    .X(net1020));
 sky130_fd_sc_hd__buf_6 fanout1021 (.A(net1022),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout1022 (.A(_07160_),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_4 fanout1023 (.A(_06546_),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_2 fanout1024 (.A(net1026),
    .X(net1024));
 sky130_fd_sc_hd__buf_6 fanout1025 (.A(net1026),
    .X(net1025));
 sky130_fd_sc_hd__buf_8 fanout1026 (.A(_06546_),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_4 fanout1027 (.A(net1030),
    .X(net1027));
 sky130_fd_sc_hd__buf_2 fanout1028 (.A(net1030),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_4 fanout1029 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_2 fanout1030 (.A(_04650_),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_4 fanout1031 (.A(net1032),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_4 fanout1032 (.A(net1034),
    .X(net1032));
 sky130_fd_sc_hd__clkbuf_4 fanout1033 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_2 fanout1034 (.A(_04564_),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_4 fanout1035 (.A(net1036),
    .X(net1035));
 sky130_fd_sc_hd__buf_4 fanout1036 (.A(_04479_),
    .X(net1036));
 sky130_fd_sc_hd__clkbuf_4 fanout1037 (.A(net1038),
    .X(net1037));
 sky130_fd_sc_hd__buf_2 fanout1038 (.A(_04479_),
    .X(net1038));
 sky130_fd_sc_hd__buf_4 fanout1039 (.A(net1040),
    .X(net1039));
 sky130_fd_sc_hd__clkbuf_4 fanout1040 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__clkbuf_4 fanout1041 (.A(_04073_),
    .X(net1041));
 sky130_fd_sc_hd__buf_4 fanout1042 (.A(_04072_),
    .X(net1042));
 sky130_fd_sc_hd__buf_12 fanout1043 (.A(_04070_),
    .X(net1043));
 sky130_fd_sc_hd__clkbuf_16 fanout1044 (.A(_03946_),
    .X(net1044));
 sky130_fd_sc_hd__buf_8 fanout1045 (.A(_03946_),
    .X(net1045));
 sky130_fd_sc_hd__buf_12 fanout1046 (.A(_03945_),
    .X(net1046));
 sky130_fd_sc_hd__buf_4 fanout1047 (.A(net1048),
    .X(net1047));
 sky130_fd_sc_hd__buf_4 fanout1048 (.A(net1051),
    .X(net1048));
 sky130_fd_sc_hd__buf_6 fanout1049 (.A(net1051),
    .X(net1049));
 sky130_fd_sc_hd__buf_2 fanout1050 (.A(net1051),
    .X(net1050));
 sky130_fd_sc_hd__buf_6 fanout1051 (.A(net443),
    .X(net1051));
 sky130_fd_sc_hd__buf_6 fanout1052 (.A(net1054),
    .X(net1052));
 sky130_fd_sc_hd__buf_6 fanout1053 (.A(net1054),
    .X(net1053));
 sky130_fd_sc_hd__buf_6 fanout1054 (.A(_03769_),
    .X(net1054));
 sky130_fd_sc_hd__buf_6 fanout1055 (.A(_02277_),
    .X(net1055));
 sky130_fd_sc_hd__clkbuf_4 fanout1056 (.A(_02277_),
    .X(net1056));
 sky130_fd_sc_hd__buf_6 fanout1057 (.A(net1058),
    .X(net1057));
 sky130_fd_sc_hd__buf_8 fanout1058 (.A(_02277_),
    .X(net1058));
 sky130_fd_sc_hd__clkbuf_8 fanout1059 (.A(_08012_),
    .X(net1059));
 sky130_fd_sc_hd__clkbuf_8 fanout1060 (.A(_07444_),
    .X(net1060));
 sky130_fd_sc_hd__buf_4 fanout1061 (.A(_07444_),
    .X(net1061));
 sky130_fd_sc_hd__clkbuf_4 fanout1062 (.A(net1064),
    .X(net1062));
 sky130_fd_sc_hd__buf_2 fanout1063 (.A(net1064),
    .X(net1063));
 sky130_fd_sc_hd__buf_6 fanout1064 (.A(net1067),
    .X(net1064));
 sky130_fd_sc_hd__buf_4 fanout1065 (.A(net1067),
    .X(net1065));
 sky130_fd_sc_hd__buf_2 fanout1066 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_4 fanout1067 (.A(_07443_),
    .X(net1067));
 sky130_fd_sc_hd__buf_4 fanout1068 (.A(_07163_),
    .X(net1068));
 sky130_fd_sc_hd__clkbuf_4 fanout1069 (.A(net1070),
    .X(net1069));
 sky130_fd_sc_hd__buf_4 fanout1070 (.A(net1075),
    .X(net1070));
 sky130_fd_sc_hd__buf_6 fanout1071 (.A(net1075),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_4 fanout1072 (.A(net1075),
    .X(net1072));
 sky130_fd_sc_hd__clkbuf_4 fanout1073 (.A(net1075),
    .X(net1073));
 sky130_fd_sc_hd__clkbuf_2 fanout1074 (.A(net1075),
    .X(net1074));
 sky130_fd_sc_hd__buf_4 fanout1075 (.A(_07162_),
    .X(net1075));
 sky130_fd_sc_hd__clkbuf_4 fanout1076 (.A(net1079),
    .X(net1076));
 sky130_fd_sc_hd__buf_2 fanout1077 (.A(net1079),
    .X(net1077));
 sky130_fd_sc_hd__clkbuf_4 fanout1078 (.A(net1079),
    .X(net1078));
 sky130_fd_sc_hd__buf_6 fanout1079 (.A(_04983_),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_4 fanout1080 (.A(net1084),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_2 fanout1081 (.A(net1084),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_4 fanout1082 (.A(net1084),
    .X(net1082));
 sky130_fd_sc_hd__clkbuf_2 fanout1083 (.A(net1084),
    .X(net1083));
 sky130_fd_sc_hd__clkbuf_8 fanout1084 (.A(_04899_),
    .X(net1084));
 sky130_fd_sc_hd__clkbuf_4 fanout1085 (.A(net1086),
    .X(net1085));
 sky130_fd_sc_hd__clkbuf_4 fanout1086 (.A(net1087),
    .X(net1086));
 sky130_fd_sc_hd__clkbuf_4 fanout1087 (.A(_04813_),
    .X(net1087));
 sky130_fd_sc_hd__clkbuf_4 fanout1088 (.A(_04813_),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_4 fanout1089 (.A(net1090),
    .X(net1089));
 sky130_fd_sc_hd__clkbuf_4 fanout1090 (.A(net1091),
    .X(net1090));
 sky130_fd_sc_hd__buf_2 fanout1091 (.A(net1092),
    .X(net1091));
 sky130_fd_sc_hd__buf_2 fanout1092 (.A(_04730_),
    .X(net1092));
 sky130_fd_sc_hd__buf_6 fanout1093 (.A(_04069_),
    .X(net1093));
 sky130_fd_sc_hd__buf_6 fanout1094 (.A(net1097),
    .X(net1094));
 sky130_fd_sc_hd__clkbuf_16 fanout1095 (.A(net1096),
    .X(net1095));
 sky130_fd_sc_hd__buf_12 fanout1096 (.A(net1097),
    .X(net1096));
 sky130_fd_sc_hd__buf_8 fanout1097 (.A(_04043_),
    .X(net1097));
 sky130_fd_sc_hd__buf_6 fanout1098 (.A(net1099),
    .X(net1098));
 sky130_fd_sc_hd__buf_4 fanout1099 (.A(_03872_),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_8 fanout1100 (.A(_03872_),
    .X(net1100));
 sky130_fd_sc_hd__buf_2 fanout1101 (.A(_03872_),
    .X(net1101));
 sky130_fd_sc_hd__buf_6 fanout1102 (.A(_02238_),
    .X(net1102));
 sky130_fd_sc_hd__buf_4 fanout1103 (.A(_02238_),
    .X(net1103));
 sky130_fd_sc_hd__buf_6 fanout1104 (.A(_07291_),
    .X(net1104));
 sky130_fd_sc_hd__buf_4 fanout1105 (.A(_07291_),
    .X(net1105));
 sky130_fd_sc_hd__buf_6 fanout1106 (.A(_07290_),
    .X(net1106));
 sky130_fd_sc_hd__buf_2 fanout1107 (.A(_07290_),
    .X(net1107));
 sky130_fd_sc_hd__buf_6 fanout1108 (.A(_07289_),
    .X(net1108));
 sky130_fd_sc_hd__clkbuf_8 fanout1109 (.A(net1110),
    .X(net1109));
 sky130_fd_sc_hd__buf_6 fanout1110 (.A(_07288_),
    .X(net1110));
 sky130_fd_sc_hd__buf_6 fanout1111 (.A(_07157_),
    .X(net1111));
 sky130_fd_sc_hd__buf_4 fanout1112 (.A(net1113),
    .X(net1112));
 sky130_fd_sc_hd__clkbuf_8 fanout1113 (.A(_07156_),
    .X(net1113));
 sky130_fd_sc_hd__buf_6 fanout1114 (.A(net1115),
    .X(net1114));
 sky130_fd_sc_hd__buf_4 fanout1115 (.A(_07154_),
    .X(net1115));
 sky130_fd_sc_hd__clkbuf_4 fanout1116 (.A(net1117),
    .X(net1116));
 sky130_fd_sc_hd__buf_4 fanout1117 (.A(_07153_),
    .X(net1117));
 sky130_fd_sc_hd__buf_4 fanout1118 (.A(net1119),
    .X(net1118));
 sky130_fd_sc_hd__buf_4 fanout1119 (.A(_07149_),
    .X(net1119));
 sky130_fd_sc_hd__buf_4 fanout1120 (.A(net1121),
    .X(net1120));
 sky130_fd_sc_hd__buf_4 fanout1121 (.A(_07139_),
    .X(net1121));
 sky130_fd_sc_hd__buf_6 fanout1122 (.A(net1124),
    .X(net1122));
 sky130_fd_sc_hd__buf_2 fanout1123 (.A(net1124),
    .X(net1123));
 sky130_fd_sc_hd__buf_4 fanout1124 (.A(_07138_),
    .X(net1124));
 sky130_fd_sc_hd__buf_6 fanout1125 (.A(net1126),
    .X(net1125));
 sky130_fd_sc_hd__buf_4 fanout1126 (.A(_07058_),
    .X(net1126));
 sky130_fd_sc_hd__buf_4 fanout1127 (.A(net1128),
    .X(net1127));
 sky130_fd_sc_hd__clkbuf_4 fanout1128 (.A(net1129),
    .X(net1128));
 sky130_fd_sc_hd__buf_4 fanout1129 (.A(_07058_),
    .X(net1129));
 sky130_fd_sc_hd__buf_6 fanout1130 (.A(_07057_),
    .X(net1130));
 sky130_fd_sc_hd__buf_6 fanout1131 (.A(_07057_),
    .X(net1131));
 sky130_fd_sc_hd__clkbuf_8 fanout1132 (.A(net1135),
    .X(net1132));
 sky130_fd_sc_hd__buf_4 fanout1133 (.A(net1134),
    .X(net1133));
 sky130_fd_sc_hd__buf_4 fanout1134 (.A(net1135),
    .X(net1134));
 sky130_fd_sc_hd__buf_4 fanout1135 (.A(_07054_),
    .X(net1135));
 sky130_fd_sc_hd__buf_8 fanout1136 (.A(_07053_),
    .X(net1136));
 sky130_fd_sc_hd__clkbuf_4 fanout1137 (.A(net1138),
    .X(net1137));
 sky130_fd_sc_hd__clkbuf_4 fanout1138 (.A(net1139),
    .X(net1138));
 sky130_fd_sc_hd__clkbuf_4 fanout1139 (.A(net1140),
    .X(net1139));
 sky130_fd_sc_hd__buf_6 fanout1140 (.A(_04422_),
    .X(net1140));
 sky130_fd_sc_hd__buf_6 fanout1141 (.A(net1142),
    .X(net1141));
 sky130_fd_sc_hd__buf_8 fanout1142 (.A(net1143),
    .X(net1142));
 sky130_fd_sc_hd__buf_8 fanout1143 (.A(net1147),
    .X(net1143));
 sky130_fd_sc_hd__buf_8 fanout1144 (.A(net1145),
    .X(net1144));
 sky130_fd_sc_hd__clkbuf_4 fanout1145 (.A(net1147),
    .X(net1145));
 sky130_fd_sc_hd__buf_12 fanout1146 (.A(net1147),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_16 fanout1147 (.A(_04092_),
    .X(net1147));
 sky130_fd_sc_hd__buf_12 fanout1148 (.A(_04091_),
    .X(net1148));
 sky130_fd_sc_hd__buf_8 fanout1149 (.A(_04091_),
    .X(net1149));
 sky130_fd_sc_hd__buf_6 fanout1150 (.A(_04068_),
    .X(net1150));
 sky130_fd_sc_hd__buf_6 fanout1151 (.A(_04067_),
    .X(net1151));
 sky130_fd_sc_hd__buf_2 fanout1152 (.A(net1153),
    .X(net1152));
 sky130_fd_sc_hd__buf_8 fanout1153 (.A(_04067_),
    .X(net1153));
 sky130_fd_sc_hd__buf_6 fanout1154 (.A(_04056_),
    .X(net1154));
 sky130_fd_sc_hd__clkbuf_8 fanout1155 (.A(net1158),
    .X(net1155));
 sky130_fd_sc_hd__buf_4 fanout1156 (.A(net1157),
    .X(net1156));
 sky130_fd_sc_hd__clkbuf_8 fanout1157 (.A(net1158),
    .X(net1157));
 sky130_fd_sc_hd__clkbuf_4 fanout1158 (.A(_02993_),
    .X(net1158));
 sky130_fd_sc_hd__clkbuf_8 fanout1159 (.A(net1162),
    .X(net1159));
 sky130_fd_sc_hd__buf_4 fanout1160 (.A(net1161),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_8 fanout1161 (.A(net1162),
    .X(net1161));
 sky130_fd_sc_hd__buf_4 fanout1162 (.A(_02992_),
    .X(net1162));
 sky130_fd_sc_hd__clkbuf_4 fanout1163 (.A(_02923_),
    .X(net1163));
 sky130_fd_sc_hd__buf_2 fanout1164 (.A(_02923_),
    .X(net1164));
 sky130_fd_sc_hd__clkbuf_4 fanout1165 (.A(net1166),
    .X(net1165));
 sky130_fd_sc_hd__clkbuf_2 fanout1166 (.A(_02923_),
    .X(net1166));
 sky130_fd_sc_hd__buf_4 fanout1167 (.A(_02922_),
    .X(net1167));
 sky130_fd_sc_hd__buf_2 fanout1168 (.A(_02922_),
    .X(net1168));
 sky130_fd_sc_hd__buf_4 fanout1169 (.A(net1170),
    .X(net1169));
 sky130_fd_sc_hd__clkbuf_4 fanout1170 (.A(_02922_),
    .X(net1170));
 sky130_fd_sc_hd__buf_4 fanout1171 (.A(net1174),
    .X(net1171));
 sky130_fd_sc_hd__buf_4 fanout1172 (.A(net1174),
    .X(net1172));
 sky130_fd_sc_hd__buf_4 fanout1173 (.A(net1174),
    .X(net1173));
 sky130_fd_sc_hd__buf_2 fanout1174 (.A(_02921_),
    .X(net1174));
 sky130_fd_sc_hd__buf_6 fanout1175 (.A(net1176),
    .X(net1175));
 sky130_fd_sc_hd__buf_6 fanout1176 (.A(_08706_),
    .X(net1176));
 sky130_fd_sc_hd__clkbuf_8 fanout1177 (.A(_07951_),
    .X(net1177));
 sky130_fd_sc_hd__clkbuf_4 fanout1178 (.A(_07951_),
    .X(net1178));
 sky130_fd_sc_hd__buf_4 fanout1179 (.A(net1180),
    .X(net1179));
 sky130_fd_sc_hd__buf_4 fanout1180 (.A(net1184),
    .X(net1180));
 sky130_fd_sc_hd__clkbuf_8 fanout1181 (.A(net1182),
    .X(net1181));
 sky130_fd_sc_hd__buf_4 fanout1182 (.A(net1183),
    .X(net1182));
 sky130_fd_sc_hd__buf_4 fanout1183 (.A(net1184),
    .X(net1183));
 sky130_fd_sc_hd__clkbuf_4 fanout1184 (.A(_07052_),
    .X(net1184));
 sky130_fd_sc_hd__buf_6 fanout1185 (.A(_07051_),
    .X(net1185));
 sky130_fd_sc_hd__buf_4 fanout1186 (.A(_05071_),
    .X(net1186));
 sky130_fd_sc_hd__clkbuf_2 fanout1187 (.A(_05071_),
    .X(net1187));
 sky130_fd_sc_hd__buf_6 fanout1188 (.A(net1189),
    .X(net1188));
 sky130_fd_sc_hd__buf_8 fanout1189 (.A(_03934_),
    .X(net1189));
 sky130_fd_sc_hd__clkbuf_8 fanout1190 (.A(net1193),
    .X(net1190));
 sky130_fd_sc_hd__buf_4 fanout1191 (.A(net1192),
    .X(net1191));
 sky130_fd_sc_hd__buf_4 fanout1192 (.A(net1193),
    .X(net1192));
 sky130_fd_sc_hd__buf_4 fanout1193 (.A(_02991_),
    .X(net1193));
 sky130_fd_sc_hd__buf_4 fanout1194 (.A(net1195),
    .X(net1194));
 sky130_fd_sc_hd__buf_4 fanout1195 (.A(net1196),
    .X(net1195));
 sky130_fd_sc_hd__buf_2 fanout1196 (.A(net1197),
    .X(net1196));
 sky130_fd_sc_hd__buf_6 fanout1197 (.A(_02909_),
    .X(net1197));
 sky130_fd_sc_hd__clkbuf_8 fanout1198 (.A(net1199),
    .X(net1198));
 sky130_fd_sc_hd__buf_6 fanout1199 (.A(_07538_),
    .X(net1199));
 sky130_fd_sc_hd__buf_8 fanout1200 (.A(net1202),
    .X(net1200));
 sky130_fd_sc_hd__buf_6 fanout1201 (.A(_07457_),
    .X(net1201));
 sky130_fd_sc_hd__buf_2 fanout1202 (.A(_07457_),
    .X(net1202));
 sky130_fd_sc_hd__buf_6 fanout1203 (.A(_07456_),
    .X(net1203));
 sky130_fd_sc_hd__buf_4 fanout1204 (.A(_07456_),
    .X(net1204));
 sky130_fd_sc_hd__buf_8 fanout1205 (.A(_07455_),
    .X(net1205));
 sky130_fd_sc_hd__buf_6 fanout1206 (.A(_07455_),
    .X(net1206));
 sky130_fd_sc_hd__clkbuf_8 fanout1207 (.A(_07369_),
    .X(net1207));
 sky130_fd_sc_hd__buf_2 fanout1208 (.A(_07369_),
    .X(net1208));
 sky130_fd_sc_hd__buf_6 fanout1209 (.A(_07369_),
    .X(net1209));
 sky130_fd_sc_hd__buf_4 fanout1210 (.A(net1212),
    .X(net1210));
 sky130_fd_sc_hd__clkbuf_4 fanout1211 (.A(net1212),
    .X(net1211));
 sky130_fd_sc_hd__buf_4 fanout1212 (.A(_07369_),
    .X(net1212));
 sky130_fd_sc_hd__buf_6 fanout1213 (.A(net1214),
    .X(net1213));
 sky130_fd_sc_hd__buf_6 fanout1214 (.A(_07368_),
    .X(net1214));
 sky130_fd_sc_hd__buf_6 fanout1215 (.A(net1216),
    .X(net1215));
 sky130_fd_sc_hd__clkbuf_8 fanout1216 (.A(net1218),
    .X(net1216));
 sky130_fd_sc_hd__clkbuf_4 fanout1217 (.A(net1218),
    .X(net1217));
 sky130_fd_sc_hd__buf_4 fanout1218 (.A(_07143_),
    .X(net1218));
 sky130_fd_sc_hd__buf_6 fanout1219 (.A(net1220),
    .X(net1219));
 sky130_fd_sc_hd__buf_8 fanout1220 (.A(_07141_),
    .X(net1220));
 sky130_fd_sc_hd__buf_8 fanout1221 (.A(net1223),
    .X(net1221));
 sky130_fd_sc_hd__buf_4 fanout1222 (.A(net1223),
    .X(net1222));
 sky130_fd_sc_hd__buf_4 fanout1223 (.A(_07049_),
    .X(net1223));
 sky130_fd_sc_hd__buf_4 fanout1224 (.A(net1225),
    .X(net1224));
 sky130_fd_sc_hd__buf_4 fanout1225 (.A(net1226),
    .X(net1225));
 sky130_fd_sc_hd__clkbuf_4 fanout1226 (.A(_07049_),
    .X(net1226));
 sky130_fd_sc_hd__buf_4 fanout1227 (.A(net1228),
    .X(net1227));
 sky130_fd_sc_hd__buf_2 fanout1228 (.A(net1229),
    .X(net1228));
 sky130_fd_sc_hd__buf_6 fanout1229 (.A(_07048_),
    .X(net1229));
 sky130_fd_sc_hd__buf_6 fanout1230 (.A(net1232),
    .X(net1230));
 sky130_fd_sc_hd__buf_6 fanout1231 (.A(net1232),
    .X(net1231));
 sky130_fd_sc_hd__buf_4 fanout1232 (.A(_07012_),
    .X(net1232));
 sky130_fd_sc_hd__clkbuf_8 fanout1233 (.A(_07000_),
    .X(net1233));
 sky130_fd_sc_hd__buf_6 fanout1234 (.A(_07000_),
    .X(net1234));
 sky130_fd_sc_hd__clkbuf_4 fanout1235 (.A(_07000_),
    .X(net1235));
 sky130_fd_sc_hd__buf_4 fanout1237 (.A(_04887_),
    .X(net1237));
 sky130_fd_sc_hd__buf_4 fanout1238 (.A(_04887_),
    .X(net1238));
 sky130_fd_sc_hd__clkbuf_16 fanout1239 (.A(net1240),
    .X(net1239));
 sky130_fd_sc_hd__buf_12 fanout1240 (.A(_04096_),
    .X(net1240));
 sky130_fd_sc_hd__clkbuf_8 fanout1241 (.A(_04096_),
    .X(net1241));
 sky130_fd_sc_hd__buf_4 fanout1242 (.A(_04030_),
    .X(net1242));
 sky130_fd_sc_hd__clkbuf_8 fanout1243 (.A(_04021_),
    .X(net1243));
 sky130_fd_sc_hd__buf_8 fanout1244 (.A(_03932_),
    .X(net1244));
 sky130_fd_sc_hd__buf_4 fanout1245 (.A(net1246),
    .X(net1245));
 sky130_fd_sc_hd__buf_6 fanout1246 (.A(_03932_),
    .X(net1246));
 sky130_fd_sc_hd__buf_6 fanout1247 (.A(net1248),
    .X(net1247));
 sky130_fd_sc_hd__buf_4 fanout1248 (.A(_03918_),
    .X(net1248));
 sky130_fd_sc_hd__clkbuf_8 fanout1249 (.A(_03918_),
    .X(net1249));
 sky130_fd_sc_hd__buf_4 fanout1250 (.A(_03918_),
    .X(net1250));
 sky130_fd_sc_hd__buf_12 fanout1251 (.A(net1256),
    .X(net1251));
 sky130_fd_sc_hd__buf_6 fanout1252 (.A(net1253),
    .X(net1252));
 sky130_fd_sc_hd__buf_4 fanout1253 (.A(net1256),
    .X(net1253));
 sky130_fd_sc_hd__buf_6 fanout1254 (.A(net1256),
    .X(net1254));
 sky130_fd_sc_hd__buf_2 fanout1255 (.A(net1256),
    .X(net1255));
 sky130_fd_sc_hd__buf_8 fanout1256 (.A(_03879_),
    .X(net1256));
 sky130_fd_sc_hd__clkbuf_8 fanout1257 (.A(net1258),
    .X(net1257));
 sky130_fd_sc_hd__buf_4 fanout1258 (.A(net1259),
    .X(net1258));
 sky130_fd_sc_hd__buf_4 fanout1259 (.A(_03879_),
    .X(net1259));
 sky130_fd_sc_hd__buf_8 fanout1260 (.A(net1261),
    .X(net1260));
 sky130_fd_sc_hd__buf_6 fanout1261 (.A(net1262),
    .X(net1261));
 sky130_fd_sc_hd__clkbuf_4 fanout1262 (.A(_03879_),
    .X(net1262));
 sky130_fd_sc_hd__buf_12 fanout1263 (.A(_03878_),
    .X(net1263));
 sky130_fd_sc_hd__clkbuf_4 fanout1264 (.A(_03878_),
    .X(net1264));
 sky130_fd_sc_hd__buf_8 fanout1265 (.A(net1267),
    .X(net1265));
 sky130_fd_sc_hd__buf_6 fanout1266 (.A(net1267),
    .X(net1266));
 sky130_fd_sc_hd__buf_6 fanout1267 (.A(_03878_),
    .X(net1267));
 sky130_fd_sc_hd__buf_4 fanout1268 (.A(net1271),
    .X(net1268));
 sky130_fd_sc_hd__buf_4 fanout1269 (.A(net1271),
    .X(net1269));
 sky130_fd_sc_hd__buf_4 fanout1270 (.A(net1271),
    .X(net1270));
 sky130_fd_sc_hd__buf_4 fanout1271 (.A(_08776_),
    .X(net1271));
 sky130_fd_sc_hd__buf_8 fanout1272 (.A(net1273),
    .X(net1272));
 sky130_fd_sc_hd__buf_6 fanout1273 (.A(_07011_),
    .X(net1273));
 sky130_fd_sc_hd__buf_6 fanout1274 (.A(_06999_),
    .X(net1274));
 sky130_fd_sc_hd__buf_8 fanout1275 (.A(_06999_),
    .X(net1275));
 sky130_fd_sc_hd__buf_8 fanout1276 (.A(net1277),
    .X(net1276));
 sky130_fd_sc_hd__buf_6 fanout1277 (.A(net1279),
    .X(net1277));
 sky130_fd_sc_hd__buf_6 fanout1278 (.A(net1279),
    .X(net1278));
 sky130_fd_sc_hd__buf_6 fanout1279 (.A(_06698_),
    .X(net1279));
 sky130_fd_sc_hd__buf_4 fanout1280 (.A(net1286),
    .X(net1280));
 sky130_fd_sc_hd__buf_4 fanout1281 (.A(_02919_),
    .X(net1281));
 sky130_fd_sc_hd__buf_4 fanout1282 (.A(net1284),
    .X(net1282));
 sky130_fd_sc_hd__buf_4 fanout1283 (.A(net1284),
    .X(net1283));
 sky130_fd_sc_hd__clkbuf_4 fanout1284 (.A(net1285),
    .X(net1284));
 sky130_fd_sc_hd__buf_4 fanout1285 (.A(net1286),
    .X(net1285));
 sky130_fd_sc_hd__buf_6 fanout1286 (.A(_02919_),
    .X(net1286));
 sky130_fd_sc_hd__buf_6 fanout1287 (.A(net1290),
    .X(net1287));
 sky130_fd_sc_hd__buf_2 fanout1288 (.A(net1290),
    .X(net1288));
 sky130_fd_sc_hd__buf_6 fanout1289 (.A(net1290),
    .X(net1289));
 sky130_fd_sc_hd__buf_6 fanout1290 (.A(_02210_),
    .X(net1290));
 sky130_fd_sc_hd__buf_4 fanout1291 (.A(net1294),
    .X(net1291));
 sky130_fd_sc_hd__buf_4 fanout1292 (.A(net1294),
    .X(net1292));
 sky130_fd_sc_hd__buf_4 fanout1293 (.A(net1294),
    .X(net1293));
 sky130_fd_sc_hd__clkbuf_4 fanout1294 (.A(_08777_),
    .X(net1294));
 sky130_fd_sc_hd__buf_4 fanout1295 (.A(net1298),
    .X(net1295));
 sky130_fd_sc_hd__clkbuf_4 fanout1296 (.A(net1298),
    .X(net1296));
 sky130_fd_sc_hd__clkbuf_4 fanout1297 (.A(net1298),
    .X(net1297));
 sky130_fd_sc_hd__buf_4 fanout1298 (.A(_08774_),
    .X(net1298));
 sky130_fd_sc_hd__buf_6 fanout1299 (.A(_07487_),
    .X(net1299));
 sky130_fd_sc_hd__buf_6 fanout1300 (.A(_07487_),
    .X(net1300));
 sky130_fd_sc_hd__buf_4 fanout1301 (.A(net1302),
    .X(net1301));
 sky130_fd_sc_hd__clkbuf_2 fanout1302 (.A(net1303),
    .X(net1302));
 sky130_fd_sc_hd__buf_2 fanout1303 (.A(net1304),
    .X(net1303));
 sky130_fd_sc_hd__buf_2 fanout1304 (.A(_07007_),
    .X(net1304));
 sky130_fd_sc_hd__buf_6 fanout1305 (.A(_07007_),
    .X(net1305));
 sky130_fd_sc_hd__clkbuf_4 fanout1306 (.A(net1308),
    .X(net1306));
 sky130_fd_sc_hd__buf_4 fanout1307 (.A(net1308),
    .X(net1307));
 sky130_fd_sc_hd__buf_4 fanout1308 (.A(net1309),
    .X(net1308));
 sky130_fd_sc_hd__clkbuf_2 fanout1309 (.A(_06837_),
    .X(net1309));
 sky130_fd_sc_hd__buf_4 fanout1310 (.A(net1312),
    .X(net1310));
 sky130_fd_sc_hd__clkbuf_4 fanout1311 (.A(net1312),
    .X(net1311));
 sky130_fd_sc_hd__buf_4 fanout1312 (.A(_06707_),
    .X(net1312));
 sky130_fd_sc_hd__buf_6 fanout1313 (.A(_06707_),
    .X(net1313));
 sky130_fd_sc_hd__clkbuf_4 fanout1314 (.A(_06707_),
    .X(net1314));
 sky130_fd_sc_hd__buf_6 fanout1315 (.A(net1318),
    .X(net1315));
 sky130_fd_sc_hd__buf_6 fanout1316 (.A(net1317),
    .X(net1316));
 sky130_fd_sc_hd__buf_8 fanout1317 (.A(net1318),
    .X(net1317));
 sky130_fd_sc_hd__buf_6 fanout1318 (.A(_06681_),
    .X(net1318));
 sky130_fd_sc_hd__buf_12 fanout1319 (.A(_04445_),
    .X(net1319));
 sky130_fd_sc_hd__buf_8 fanout1320 (.A(net1321),
    .X(net1320));
 sky130_fd_sc_hd__clkbuf_16 fanout1321 (.A(_04087_),
    .X(net1321));
 sky130_fd_sc_hd__clkbuf_16 fanout1322 (.A(net1323),
    .X(net1322));
 sky130_fd_sc_hd__buf_8 fanout1323 (.A(_04087_),
    .X(net1323));
 sky130_fd_sc_hd__clkbuf_16 fanout1324 (.A(_04086_),
    .X(net1324));
 sky130_fd_sc_hd__buf_4 fanout1325 (.A(_04086_),
    .X(net1325));
 sky130_fd_sc_hd__buf_12 fanout1326 (.A(net1327),
    .X(net1326));
 sky130_fd_sc_hd__clkbuf_16 fanout1327 (.A(_04086_),
    .X(net1327));
 sky130_fd_sc_hd__buf_8 fanout1328 (.A(net1329),
    .X(net1328));
 sky130_fd_sc_hd__clkbuf_16 fanout1329 (.A(net1340),
    .X(net1329));
 sky130_fd_sc_hd__buf_6 fanout1330 (.A(net1331),
    .X(net1330));
 sky130_fd_sc_hd__buf_6 fanout1331 (.A(net1340),
    .X(net1331));
 sky130_fd_sc_hd__buf_6 fanout1332 (.A(net1334),
    .X(net1332));
 sky130_fd_sc_hd__buf_6 fanout1333 (.A(net1334),
    .X(net1333));
 sky130_fd_sc_hd__buf_6 fanout1334 (.A(net1340),
    .X(net1334));
 sky130_fd_sc_hd__buf_6 fanout1335 (.A(net1339),
    .X(net1335));
 sky130_fd_sc_hd__buf_4 fanout1336 (.A(net1339),
    .X(net1336));
 sky130_fd_sc_hd__buf_6 fanout1337 (.A(net1338),
    .X(net1337));
 sky130_fd_sc_hd__buf_8 fanout1338 (.A(net1339),
    .X(net1338));
 sky130_fd_sc_hd__buf_6 fanout1339 (.A(net1340),
    .X(net1339));
 sky130_fd_sc_hd__clkbuf_16 fanout1340 (.A(_04084_),
    .X(net1340));
 sky130_fd_sc_hd__buf_8 fanout1341 (.A(net1343),
    .X(net1341));
 sky130_fd_sc_hd__buf_4 fanout1342 (.A(net1343),
    .X(net1342));
 sky130_fd_sc_hd__clkbuf_16 fanout1343 (.A(net1356),
    .X(net1343));
 sky130_fd_sc_hd__buf_8 fanout1344 (.A(net1346),
    .X(net1344));
 sky130_fd_sc_hd__buf_4 fanout1345 (.A(net1346),
    .X(net1345));
 sky130_fd_sc_hd__buf_8 fanout1346 (.A(net1356),
    .X(net1346));
 sky130_fd_sc_hd__buf_8 fanout1347 (.A(net1348),
    .X(net1347));
 sky130_fd_sc_hd__buf_6 fanout1348 (.A(net1355),
    .X(net1348));
 sky130_fd_sc_hd__buf_8 fanout1349 (.A(net1355),
    .X(net1349));
 sky130_fd_sc_hd__buf_8 fanout1350 (.A(net1355),
    .X(net1350));
 sky130_fd_sc_hd__clkbuf_4 fanout1351 (.A(net1355),
    .X(net1351));
 sky130_fd_sc_hd__buf_6 fanout1352 (.A(net1354),
    .X(net1352));
 sky130_fd_sc_hd__buf_6 fanout1353 (.A(net1354),
    .X(net1353));
 sky130_fd_sc_hd__buf_4 fanout1354 (.A(net1355),
    .X(net1354));
 sky130_fd_sc_hd__clkbuf_16 fanout1355 (.A(net1356),
    .X(net1355));
 sky130_fd_sc_hd__buf_6 fanout1356 (.A(_04083_),
    .X(net1356));
 sky130_fd_sc_hd__buf_6 fanout1357 (.A(net1358),
    .X(net1357));
 sky130_fd_sc_hd__buf_4 fanout1358 (.A(net1359),
    .X(net1358));
 sky130_fd_sc_hd__buf_6 fanout1359 (.A(_04081_),
    .X(net1359));
 sky130_fd_sc_hd__buf_6 fanout1360 (.A(net1361),
    .X(net1360));
 sky130_fd_sc_hd__buf_6 fanout1361 (.A(net1362),
    .X(net1361));
 sky130_fd_sc_hd__buf_8 fanout1362 (.A(_04081_),
    .X(net1362));
 sky130_fd_sc_hd__buf_6 fanout1363 (.A(net1364),
    .X(net1363));
 sky130_fd_sc_hd__buf_6 fanout1364 (.A(net1365),
    .X(net1364));
 sky130_fd_sc_hd__buf_6 fanout1365 (.A(net1371),
    .X(net1365));
 sky130_fd_sc_hd__buf_4 fanout1366 (.A(net1367),
    .X(net1366));
 sky130_fd_sc_hd__clkbuf_8 fanout1367 (.A(net1370),
    .X(net1367));
 sky130_fd_sc_hd__buf_6 fanout1368 (.A(net1370),
    .X(net1368));
 sky130_fd_sc_hd__clkbuf_4 fanout1369 (.A(net1370),
    .X(net1369));
 sky130_fd_sc_hd__buf_4 fanout1370 (.A(net1371),
    .X(net1370));
 sky130_fd_sc_hd__buf_4 fanout1371 (.A(net1390),
    .X(net1371));
 sky130_fd_sc_hd__buf_6 fanout1372 (.A(net1373),
    .X(net1372));
 sky130_fd_sc_hd__buf_6 fanout1373 (.A(net1374),
    .X(net1373));
 sky130_fd_sc_hd__buf_4 fanout1374 (.A(net1390),
    .X(net1374));
 sky130_fd_sc_hd__buf_6 fanout1375 (.A(net1376),
    .X(net1375));
 sky130_fd_sc_hd__clkbuf_4 fanout1376 (.A(net1390),
    .X(net1376));
 sky130_fd_sc_hd__clkbuf_8 fanout1377 (.A(net1381),
    .X(net1377));
 sky130_fd_sc_hd__clkbuf_8 fanout1378 (.A(net1381),
    .X(net1378));
 sky130_fd_sc_hd__buf_6 fanout1379 (.A(net1381),
    .X(net1379));
 sky130_fd_sc_hd__buf_4 fanout1380 (.A(net1381),
    .X(net1380));
 sky130_fd_sc_hd__clkbuf_8 fanout1381 (.A(net1386),
    .X(net1381));
 sky130_fd_sc_hd__buf_6 fanout1382 (.A(net1386),
    .X(net1382));
 sky130_fd_sc_hd__buf_6 fanout1383 (.A(net1386),
    .X(net1383));
 sky130_fd_sc_hd__buf_6 fanout1384 (.A(net1386),
    .X(net1384));
 sky130_fd_sc_hd__buf_4 fanout1385 (.A(net1386),
    .X(net1385));
 sky130_fd_sc_hd__buf_4 fanout1386 (.A(net1390),
    .X(net1386));
 sky130_fd_sc_hd__buf_6 fanout1387 (.A(net1388),
    .X(net1387));
 sky130_fd_sc_hd__buf_6 fanout1388 (.A(net1390),
    .X(net1388));
 sky130_fd_sc_hd__buf_6 fanout1389 (.A(net1390),
    .X(net1389));
 sky130_fd_sc_hd__buf_8 fanout1390 (.A(_04080_),
    .X(net1390));
 sky130_fd_sc_hd__buf_6 fanout1391 (.A(net1392),
    .X(net1391));
 sky130_fd_sc_hd__buf_6 fanout1392 (.A(net1395),
    .X(net1392));
 sky130_fd_sc_hd__buf_6 fanout1393 (.A(net1395),
    .X(net1393));
 sky130_fd_sc_hd__buf_4 fanout1394 (.A(net1395),
    .X(net1394));
 sky130_fd_sc_hd__clkbuf_8 fanout1395 (.A(net1407),
    .X(net1395));
 sky130_fd_sc_hd__buf_6 fanout1396 (.A(net1398),
    .X(net1396));
 sky130_fd_sc_hd__buf_6 fanout1397 (.A(net1398),
    .X(net1397));
 sky130_fd_sc_hd__clkbuf_4 fanout1398 (.A(net1407),
    .X(net1398));
 sky130_fd_sc_hd__buf_6 fanout1399 (.A(net1407),
    .X(net1399));
 sky130_fd_sc_hd__buf_4 fanout1400 (.A(net1407),
    .X(net1400));
 sky130_fd_sc_hd__buf_6 fanout1401 (.A(net1403),
    .X(net1401));
 sky130_fd_sc_hd__clkbuf_4 fanout1402 (.A(net1403),
    .X(net1402));
 sky130_fd_sc_hd__clkbuf_4 fanout1403 (.A(net1406),
    .X(net1403));
 sky130_fd_sc_hd__buf_6 fanout1404 (.A(net1406),
    .X(net1404));
 sky130_fd_sc_hd__buf_2 fanout1405 (.A(net1406),
    .X(net1405));
 sky130_fd_sc_hd__buf_4 fanout1406 (.A(net1407),
    .X(net1406));
 sky130_fd_sc_hd__buf_4 fanout1407 (.A(_04080_),
    .X(net1407));
 sky130_fd_sc_hd__buf_6 fanout1408 (.A(net1415),
    .X(net1408));
 sky130_fd_sc_hd__clkbuf_4 fanout1409 (.A(net1415),
    .X(net1409));
 sky130_fd_sc_hd__buf_6 fanout1410 (.A(net1415),
    .X(net1410));
 sky130_fd_sc_hd__buf_4 fanout1411 (.A(net1415),
    .X(net1411));
 sky130_fd_sc_hd__buf_6 fanout1412 (.A(net1415),
    .X(net1412));
 sky130_fd_sc_hd__clkbuf_4 fanout1413 (.A(net1415),
    .X(net1413));
 sky130_fd_sc_hd__buf_6 fanout1414 (.A(net1415),
    .X(net1414));
 sky130_fd_sc_hd__buf_6 fanout1415 (.A(_04080_),
    .X(net1415));
 sky130_fd_sc_hd__clkbuf_8 fanout1416 (.A(net1417),
    .X(net1416));
 sky130_fd_sc_hd__clkbuf_8 fanout1417 (.A(net1426),
    .X(net1417));
 sky130_fd_sc_hd__buf_6 fanout1418 (.A(net1419),
    .X(net1418));
 sky130_fd_sc_hd__buf_4 fanout1419 (.A(net1426),
    .X(net1419));
 sky130_fd_sc_hd__buf_4 fanout1420 (.A(net1422),
    .X(net1420));
 sky130_fd_sc_hd__buf_6 fanout1421 (.A(net1426),
    .X(net1421));
 sky130_fd_sc_hd__buf_2 fanout1422 (.A(net1426),
    .X(net1422));
 sky130_fd_sc_hd__buf_4 fanout1423 (.A(net1425),
    .X(net1423));
 sky130_fd_sc_hd__buf_4 fanout1424 (.A(net1426),
    .X(net1424));
 sky130_fd_sc_hd__clkbuf_4 fanout1425 (.A(net1426),
    .X(net1425));
 sky130_fd_sc_hd__buf_6 fanout1426 (.A(_04080_),
    .X(net1426));
 sky130_fd_sc_hd__buf_12 fanout1427 (.A(net1428),
    .X(net1427));
 sky130_fd_sc_hd__buf_12 fanout1428 (.A(_04077_),
    .X(net1428));
 sky130_fd_sc_hd__clkbuf_16 fanout1429 (.A(net1431),
    .X(net1429));
 sky130_fd_sc_hd__buf_4 fanout1430 (.A(net1431),
    .X(net1430));
 sky130_fd_sc_hd__buf_12 fanout1431 (.A(_04076_),
    .X(net1431));
 sky130_fd_sc_hd__buf_8 fanout1432 (.A(net1433),
    .X(net1432));
 sky130_fd_sc_hd__buf_12 fanout1433 (.A(_04076_),
    .X(net1433));
 sky130_fd_sc_hd__buf_6 fanout1434 (.A(net1436),
    .X(net1434));
 sky130_fd_sc_hd__buf_6 fanout1435 (.A(net1436),
    .X(net1435));
 sky130_fd_sc_hd__clkbuf_8 fanout1436 (.A(net1437),
    .X(net1436));
 sky130_fd_sc_hd__buf_4 fanout1437 (.A(_04075_),
    .X(net1437));
 sky130_fd_sc_hd__buf_6 fanout1438 (.A(net1440),
    .X(net1438));
 sky130_fd_sc_hd__clkbuf_4 fanout1439 (.A(net1440),
    .X(net1439));
 sky130_fd_sc_hd__buf_4 fanout1440 (.A(_04075_),
    .X(net1440));
 sky130_fd_sc_hd__buf_8 fanout1441 (.A(net1442),
    .X(net1441));
 sky130_fd_sc_hd__clkbuf_8 fanout1442 (.A(net1446),
    .X(net1442));
 sky130_fd_sc_hd__buf_8 fanout1443 (.A(net1446),
    .X(net1443));
 sky130_fd_sc_hd__buf_6 fanout1444 (.A(net1445),
    .X(net1444));
 sky130_fd_sc_hd__buf_4 fanout1445 (.A(net1446),
    .X(net1445));
 sky130_fd_sc_hd__buf_6 fanout1446 (.A(_04075_),
    .X(net1446));
 sky130_fd_sc_hd__buf_6 fanout1447 (.A(net1448),
    .X(net1447));
 sky130_fd_sc_hd__buf_8 fanout1448 (.A(net1449),
    .X(net1448));
 sky130_fd_sc_hd__buf_6 fanout1449 (.A(_04074_),
    .X(net1449));
 sky130_fd_sc_hd__buf_6 fanout1450 (.A(net1452),
    .X(net1450));
 sky130_fd_sc_hd__buf_4 fanout1451 (.A(net1452),
    .X(net1451));
 sky130_fd_sc_hd__buf_4 fanout1452 (.A(_04074_),
    .X(net1452));
 sky130_fd_sc_hd__buf_6 fanout1453 (.A(net1457),
    .X(net1453));
 sky130_fd_sc_hd__buf_6 fanout1454 (.A(net1457),
    .X(net1454));
 sky130_fd_sc_hd__buf_6 fanout1455 (.A(net1456),
    .X(net1455));
 sky130_fd_sc_hd__buf_4 fanout1456 (.A(net1457),
    .X(net1456));
 sky130_fd_sc_hd__buf_12 fanout1457 (.A(_04074_),
    .X(net1457));
 sky130_fd_sc_hd__buf_4 fanout1458 (.A(_03988_),
    .X(net1458));
 sky130_fd_sc_hd__buf_12 fanout1459 (.A(net1461),
    .X(net1459));
 sky130_fd_sc_hd__buf_12 fanout1460 (.A(net1461),
    .X(net1460));
 sky130_fd_sc_hd__buf_8 fanout1461 (.A(_03890_),
    .X(net1461));
 sky130_fd_sc_hd__buf_6 fanout1462 (.A(net1463),
    .X(net1462));
 sky130_fd_sc_hd__buf_6 fanout1463 (.A(net1464),
    .X(net1463));
 sky130_fd_sc_hd__buf_6 fanout1464 (.A(net1469),
    .X(net1464));
 sky130_fd_sc_hd__buf_6 fanout1465 (.A(net1469),
    .X(net1465));
 sky130_fd_sc_hd__buf_4 fanout1466 (.A(net1469),
    .X(net1466));
 sky130_fd_sc_hd__buf_6 fanout1467 (.A(net1469),
    .X(net1467));
 sky130_fd_sc_hd__clkbuf_4 fanout1468 (.A(net1469),
    .X(net1468));
 sky130_fd_sc_hd__clkbuf_8 fanout1469 (.A(net1525),
    .X(net1469));
 sky130_fd_sc_hd__buf_6 fanout1470 (.A(net1472),
    .X(net1470));
 sky130_fd_sc_hd__clkbuf_4 fanout1471 (.A(net1472),
    .X(net1471));
 sky130_fd_sc_hd__buf_6 fanout1472 (.A(net1475),
    .X(net1472));
 sky130_fd_sc_hd__buf_6 fanout1473 (.A(net1475),
    .X(net1473));
 sky130_fd_sc_hd__buf_4 fanout1474 (.A(net1475),
    .X(net1474));
 sky130_fd_sc_hd__buf_6 fanout1475 (.A(net1525),
    .X(net1475));
 sky130_fd_sc_hd__buf_6 fanout1476 (.A(net1477),
    .X(net1476));
 sky130_fd_sc_hd__buf_6 fanout1477 (.A(net1480),
    .X(net1477));
 sky130_fd_sc_hd__buf_6 fanout1478 (.A(net1480),
    .X(net1478));
 sky130_fd_sc_hd__buf_4 fanout1479 (.A(net1480),
    .X(net1479));
 sky130_fd_sc_hd__buf_4 fanout1480 (.A(net1485),
    .X(net1480));
 sky130_fd_sc_hd__buf_6 fanout1481 (.A(net1485),
    .X(net1481));
 sky130_fd_sc_hd__clkbuf_8 fanout1482 (.A(net1485),
    .X(net1482));
 sky130_fd_sc_hd__buf_6 fanout1483 (.A(net1485),
    .X(net1483));
 sky130_fd_sc_hd__buf_6 fanout1484 (.A(net1485),
    .X(net1484));
 sky130_fd_sc_hd__buf_4 fanout1485 (.A(net1525),
    .X(net1485));
 sky130_fd_sc_hd__buf_6 fanout1486 (.A(net1489),
    .X(net1486));
 sky130_fd_sc_hd__buf_6 fanout1487 (.A(net1488),
    .X(net1487));
 sky130_fd_sc_hd__buf_4 fanout1488 (.A(net1489),
    .X(net1488));
 sky130_fd_sc_hd__clkbuf_4 fanout1489 (.A(net1525),
    .X(net1489));
 sky130_fd_sc_hd__buf_6 fanout1490 (.A(net1494),
    .X(net1490));
 sky130_fd_sc_hd__buf_6 fanout1491 (.A(net1494),
    .X(net1491));
 sky130_fd_sc_hd__buf_6 fanout1492 (.A(net1494),
    .X(net1492));
 sky130_fd_sc_hd__clkbuf_4 fanout1493 (.A(net1494),
    .X(net1493));
 sky130_fd_sc_hd__buf_6 fanout1494 (.A(net1525),
    .X(net1494));
 sky130_fd_sc_hd__buf_6 fanout1495 (.A(net1496),
    .X(net1495));
 sky130_fd_sc_hd__buf_6 fanout1496 (.A(net1499),
    .X(net1496));
 sky130_fd_sc_hd__buf_6 fanout1497 (.A(net1499),
    .X(net1497));
 sky130_fd_sc_hd__clkbuf_4 fanout1498 (.A(net1499),
    .X(net1498));
 sky130_fd_sc_hd__buf_4 fanout1499 (.A(net1525),
    .X(net1499));
 sky130_fd_sc_hd__buf_6 fanout1500 (.A(net1502),
    .X(net1500));
 sky130_fd_sc_hd__buf_4 fanout1501 (.A(net1502),
    .X(net1501));
 sky130_fd_sc_hd__clkbuf_4 fanout1502 (.A(net1505),
    .X(net1502));
 sky130_fd_sc_hd__buf_6 fanout1503 (.A(net1505),
    .X(net1503));
 sky130_fd_sc_hd__clkbuf_8 fanout1504 (.A(net1505),
    .X(net1504));
 sky130_fd_sc_hd__buf_4 fanout1505 (.A(net1525),
    .X(net1505));
 sky130_fd_sc_hd__buf_6 fanout1506 (.A(net1514),
    .X(net1506));
 sky130_fd_sc_hd__clkbuf_4 fanout1507 (.A(net1514),
    .X(net1507));
 sky130_fd_sc_hd__buf_6 fanout1508 (.A(net1514),
    .X(net1508));
 sky130_fd_sc_hd__buf_6 fanout1509 (.A(net1514),
    .X(net1509));
 sky130_fd_sc_hd__buf_6 fanout1510 (.A(net1513),
    .X(net1510));
 sky130_fd_sc_hd__buf_6 fanout1511 (.A(net1513),
    .X(net1511));
 sky130_fd_sc_hd__clkbuf_8 fanout1512 (.A(net1513),
    .X(net1512));
 sky130_fd_sc_hd__buf_4 fanout1513 (.A(net1514),
    .X(net1513));
 sky130_fd_sc_hd__clkbuf_8 fanout1514 (.A(net1524),
    .X(net1514));
 sky130_fd_sc_hd__buf_6 fanout1515 (.A(net1524),
    .X(net1515));
 sky130_fd_sc_hd__clkbuf_4 fanout1516 (.A(net1524),
    .X(net1516));
 sky130_fd_sc_hd__buf_6 fanout1517 (.A(net1518),
    .X(net1517));
 sky130_fd_sc_hd__buf_4 fanout1518 (.A(net1524),
    .X(net1518));
 sky130_fd_sc_hd__buf_6 fanout1519 (.A(net1520),
    .X(net1519));
 sky130_fd_sc_hd__buf_6 fanout1520 (.A(net1523),
    .X(net1520));
 sky130_fd_sc_hd__buf_6 fanout1521 (.A(net1522),
    .X(net1521));
 sky130_fd_sc_hd__buf_6 fanout1522 (.A(net1523),
    .X(net1522));
 sky130_fd_sc_hd__buf_4 fanout1523 (.A(net1524),
    .X(net1523));
 sky130_fd_sc_hd__buf_4 fanout1524 (.A(net1525),
    .X(net1524));
 sky130_fd_sc_hd__buf_12 fanout1525 (.A(_03889_),
    .X(net1525));
 sky130_fd_sc_hd__buf_6 fanout1526 (.A(net1527),
    .X(net1526));
 sky130_fd_sc_hd__buf_6 fanout1527 (.A(net1529),
    .X(net1527));
 sky130_fd_sc_hd__clkbuf_4 fanout1528 (.A(net1529),
    .X(net1528));
 sky130_fd_sc_hd__buf_6 fanout1529 (.A(net1541),
    .X(net1529));
 sky130_fd_sc_hd__buf_6 fanout1530 (.A(net1532),
    .X(net1530));
 sky130_fd_sc_hd__buf_4 fanout1531 (.A(net1532),
    .X(net1531));
 sky130_fd_sc_hd__buf_6 fanout1532 (.A(net1541),
    .X(net1532));
 sky130_fd_sc_hd__buf_6 fanout1533 (.A(net1534),
    .X(net1533));
 sky130_fd_sc_hd__buf_8 fanout1534 (.A(net1541),
    .X(net1534));
 sky130_fd_sc_hd__buf_4 fanout1535 (.A(net1541),
    .X(net1535));
 sky130_fd_sc_hd__buf_6 fanout1536 (.A(net1537),
    .X(net1536));
 sky130_fd_sc_hd__buf_6 fanout1537 (.A(net1541),
    .X(net1537));
 sky130_fd_sc_hd__buf_6 fanout1538 (.A(net1540),
    .X(net1538));
 sky130_fd_sc_hd__buf_4 fanout1539 (.A(net1540),
    .X(net1539));
 sky130_fd_sc_hd__buf_8 fanout1540 (.A(net1541),
    .X(net1540));
 sky130_fd_sc_hd__buf_12 fanout1541 (.A(_03888_),
    .X(net1541));
 sky130_fd_sc_hd__buf_6 fanout1542 (.A(net1543),
    .X(net1542));
 sky130_fd_sc_hd__buf_8 fanout1543 (.A(net1545),
    .X(net1543));
 sky130_fd_sc_hd__buf_8 fanout1544 (.A(net1545),
    .X(net1544));
 sky130_fd_sc_hd__buf_4 fanout1545 (.A(_03887_),
    .X(net1545));
 sky130_fd_sc_hd__buf_6 fanout1546 (.A(net1548),
    .X(net1546));
 sky130_fd_sc_hd__buf_6 fanout1547 (.A(net1548),
    .X(net1547));
 sky130_fd_sc_hd__clkbuf_8 fanout1548 (.A(net1549),
    .X(net1548));
 sky130_fd_sc_hd__buf_6 fanout1549 (.A(_03887_),
    .X(net1549));
 sky130_fd_sc_hd__buf_6 fanout1550 (.A(net1554),
    .X(net1550));
 sky130_fd_sc_hd__buf_8 fanout1551 (.A(net1554),
    .X(net1551));
 sky130_fd_sc_hd__buf_8 fanout1552 (.A(net1554),
    .X(net1552));
 sky130_fd_sc_hd__clkbuf_4 fanout1553 (.A(net1554),
    .X(net1553));
 sky130_fd_sc_hd__buf_6 fanout1554 (.A(_03887_),
    .X(net1554));
 sky130_fd_sc_hd__buf_6 fanout1555 (.A(net1560),
    .X(net1555));
 sky130_fd_sc_hd__buf_6 fanout1556 (.A(net1560),
    .X(net1556));
 sky130_fd_sc_hd__buf_6 fanout1557 (.A(net1560),
    .X(net1557));
 sky130_fd_sc_hd__clkbuf_4 fanout1558 (.A(net1559),
    .X(net1558));
 sky130_fd_sc_hd__buf_8 fanout1559 (.A(net1560),
    .X(net1559));
 sky130_fd_sc_hd__buf_8 fanout1560 (.A(_03887_),
    .X(net1560));
 sky130_fd_sc_hd__buf_6 fanout1561 (.A(net1562),
    .X(net1561));
 sky130_fd_sc_hd__buf_12 fanout1562 (.A(_03886_),
    .X(net1562));
 sky130_fd_sc_hd__buf_8 fanout1563 (.A(net1565),
    .X(net1563));
 sky130_fd_sc_hd__buf_8 fanout1564 (.A(net1565),
    .X(net1564));
 sky130_fd_sc_hd__clkbuf_16 fanout1565 (.A(_03886_),
    .X(net1565));
 sky130_fd_sc_hd__buf_6 fanout1566 (.A(net1567),
    .X(net1566));
 sky130_fd_sc_hd__clkbuf_16 fanout1567 (.A(net1570),
    .X(net1567));
 sky130_fd_sc_hd__buf_12 fanout1568 (.A(net1569),
    .X(net1568));
 sky130_fd_sc_hd__buf_12 fanout1569 (.A(net1570),
    .X(net1569));
 sky130_fd_sc_hd__buf_12 fanout1570 (.A(_03885_),
    .X(net1570));
 sky130_fd_sc_hd__buf_8 fanout1571 (.A(net1572),
    .X(net1571));
 sky130_fd_sc_hd__clkbuf_16 fanout1572 (.A(net1573),
    .X(net1572));
 sky130_fd_sc_hd__buf_6 fanout1573 (.A(net1581),
    .X(net1573));
 sky130_fd_sc_hd__buf_8 fanout1574 (.A(net1575),
    .X(net1574));
 sky130_fd_sc_hd__buf_8 fanout1575 (.A(net1581),
    .X(net1575));
 sky130_fd_sc_hd__buf_8 fanout1576 (.A(net1581),
    .X(net1576));
 sky130_fd_sc_hd__buf_4 fanout1577 (.A(net1581),
    .X(net1577));
 sky130_fd_sc_hd__buf_8 fanout1578 (.A(net1579),
    .X(net1578));
 sky130_fd_sc_hd__buf_8 fanout1579 (.A(net1581),
    .X(net1579));
 sky130_fd_sc_hd__buf_6 fanout1580 (.A(net1581),
    .X(net1580));
 sky130_fd_sc_hd__buf_12 fanout1581 (.A(_03884_),
    .X(net1581));
 sky130_fd_sc_hd__buf_8 fanout1582 (.A(net1584),
    .X(net1582));
 sky130_fd_sc_hd__buf_4 fanout1583 (.A(net1584),
    .X(net1583));
 sky130_fd_sc_hd__buf_6 fanout1584 (.A(net1592),
    .X(net1584));
 sky130_fd_sc_hd__buf_6 fanout1585 (.A(net1586),
    .X(net1585));
 sky130_fd_sc_hd__buf_6 fanout1586 (.A(net1592),
    .X(net1586));
 sky130_fd_sc_hd__buf_8 fanout1587 (.A(net1588),
    .X(net1587));
 sky130_fd_sc_hd__buf_8 fanout1588 (.A(net1592),
    .X(net1588));
 sky130_fd_sc_hd__buf_8 fanout1589 (.A(net1592),
    .X(net1589));
 sky130_fd_sc_hd__buf_6 fanout1590 (.A(net1591),
    .X(net1590));
 sky130_fd_sc_hd__buf_6 fanout1591 (.A(net1592),
    .X(net1591));
 sky130_fd_sc_hd__buf_12 fanout1592 (.A(_03883_),
    .X(net1592));
 sky130_fd_sc_hd__buf_12 fanout1593 (.A(_03882_),
    .X(net1593));
 sky130_fd_sc_hd__clkbuf_8 fanout1594 (.A(_03882_),
    .X(net1594));
 sky130_fd_sc_hd__clkbuf_16 fanout1595 (.A(net1596),
    .X(net1595));
 sky130_fd_sc_hd__buf_12 fanout1596 (.A(_03882_),
    .X(net1596));
 sky130_fd_sc_hd__clkbuf_16 fanout1597 (.A(_03881_),
    .X(net1597));
 sky130_fd_sc_hd__buf_6 fanout1598 (.A(_03881_),
    .X(net1598));
 sky130_fd_sc_hd__buf_8 fanout1599 (.A(net1600),
    .X(net1599));
 sky130_fd_sc_hd__clkbuf_16 fanout1600 (.A(_03881_),
    .X(net1600));
 sky130_fd_sc_hd__clkbuf_16 fanout1601 (.A(_03875_),
    .X(net1601));
 sky130_fd_sc_hd__buf_4 fanout1602 (.A(_03875_),
    .X(net1602));
 sky130_fd_sc_hd__buf_4 fanout1603 (.A(net1604),
    .X(net1603));
 sky130_fd_sc_hd__buf_4 fanout1604 (.A(_02240_),
    .X(net1604));
 sky130_fd_sc_hd__buf_4 fanout1605 (.A(_02240_),
    .X(net1605));
 sky130_fd_sc_hd__buf_2 fanout1606 (.A(_02240_),
    .X(net1606));
 sky130_fd_sc_hd__buf_4 fanout1607 (.A(net1608),
    .X(net1607));
 sky130_fd_sc_hd__buf_4 fanout1608 (.A(_02239_),
    .X(net1608));
 sky130_fd_sc_hd__buf_6 fanout1609 (.A(_02239_),
    .X(net1609));
 sky130_fd_sc_hd__buf_6 fanout1610 (.A(_07009_),
    .X(net1610));
 sky130_fd_sc_hd__buf_4 fanout1611 (.A(net1613),
    .X(net1611));
 sky130_fd_sc_hd__buf_4 fanout1612 (.A(net1613),
    .X(net1612));
 sky130_fd_sc_hd__clkbuf_4 fanout1613 (.A(_07009_),
    .X(net1613));
 sky130_fd_sc_hd__buf_6 fanout1614 (.A(net1615),
    .X(net1614));
 sky130_fd_sc_hd__buf_6 fanout1615 (.A(_06693_),
    .X(net1615));
 sky130_fd_sc_hd__clkbuf_8 fanout1616 (.A(_04002_),
    .X(net1616));
 sky130_fd_sc_hd__clkbuf_8 fanout1617 (.A(_04001_),
    .X(net1617));
 sky130_fd_sc_hd__clkbuf_2 fanout1618 (.A(_04001_),
    .X(net1618));
 sky130_fd_sc_hd__buf_6 fanout1619 (.A(_03998_),
    .X(net1619));
 sky130_fd_sc_hd__clkbuf_4 fanout1620 (.A(_03998_),
    .X(net1620));
 sky130_fd_sc_hd__buf_6 fanout1621 (.A(net1622),
    .X(net1621));
 sky130_fd_sc_hd__buf_4 fanout1622 (.A(_03995_),
    .X(net1622));
 sky130_fd_sc_hd__buf_6 fanout1623 (.A(net1624),
    .X(net1623));
 sky130_fd_sc_hd__buf_4 fanout1624 (.A(_03975_),
    .X(net1624));
 sky130_fd_sc_hd__buf_4 fanout1625 (.A(net1628),
    .X(net1625));
 sky130_fd_sc_hd__clkbuf_4 fanout1626 (.A(net1627),
    .X(net1626));
 sky130_fd_sc_hd__buf_4 fanout1627 (.A(net1628),
    .X(net1627));
 sky130_fd_sc_hd__clkbuf_4 fanout1628 (.A(_03974_),
    .X(net1628));
 sky130_fd_sc_hd__buf_12 fanout1629 (.A(net1632),
    .X(net1629));
 sky130_fd_sc_hd__buf_6 fanout1630 (.A(net1632),
    .X(net1630));
 sky130_fd_sc_hd__buf_12 fanout1631 (.A(net1632),
    .X(net1631));
 sky130_fd_sc_hd__clkbuf_16 fanout1632 (.A(_03856_),
    .X(net1632));
 sky130_fd_sc_hd__buf_12 fanout1633 (.A(net1634),
    .X(net1633));
 sky130_fd_sc_hd__buf_6 fanout1634 (.A(_03855_),
    .X(net1634));
 sky130_fd_sc_hd__buf_6 fanout1635 (.A(net1637),
    .X(net1635));
 sky130_fd_sc_hd__buf_12 fanout1636 (.A(net1637),
    .X(net1636));
 sky130_fd_sc_hd__buf_8 fanout1637 (.A(_03850_),
    .X(net1637));
 sky130_fd_sc_hd__buf_4 fanout1638 (.A(net1640),
    .X(net1638));
 sky130_fd_sc_hd__buf_4 fanout1639 (.A(net1640),
    .X(net1639));
 sky130_fd_sc_hd__clkbuf_4 fanout1640 (.A(_03849_),
    .X(net1640));
 sky130_fd_sc_hd__clkbuf_8 fanout1641 (.A(net1642),
    .X(net1641));
 sky130_fd_sc_hd__buf_6 fanout1642 (.A(net1646),
    .X(net1642));
 sky130_fd_sc_hd__clkbuf_8 fanout1643 (.A(net1644),
    .X(net1643));
 sky130_fd_sc_hd__clkbuf_8 fanout1644 (.A(net1646),
    .X(net1644));
 sky130_fd_sc_hd__buf_6 fanout1645 (.A(net1646),
    .X(net1645));
 sky130_fd_sc_hd__clkbuf_8 fanout1646 (.A(net1662),
    .X(net1646));
 sky130_fd_sc_hd__buf_6 fanout1647 (.A(net1649),
    .X(net1647));
 sky130_fd_sc_hd__buf_6 fanout1648 (.A(net1649),
    .X(net1648));
 sky130_fd_sc_hd__buf_8 fanout1649 (.A(net1650),
    .X(net1649));
 sky130_fd_sc_hd__buf_8 fanout1650 (.A(net1662),
    .X(net1650));
 sky130_fd_sc_hd__buf_6 fanout1651 (.A(net1652),
    .X(net1651));
 sky130_fd_sc_hd__buf_6 fanout1652 (.A(net1655),
    .X(net1652));
 sky130_fd_sc_hd__buf_6 fanout1653 (.A(net1655),
    .X(net1653));
 sky130_fd_sc_hd__clkbuf_4 fanout1654 (.A(net1655),
    .X(net1654));
 sky130_fd_sc_hd__buf_6 fanout1655 (.A(net1662),
    .X(net1655));
 sky130_fd_sc_hd__buf_8 fanout1656 (.A(net1662),
    .X(net1656));
 sky130_fd_sc_hd__buf_4 fanout1657 (.A(net1662),
    .X(net1657));
 sky130_fd_sc_hd__clkbuf_8 fanout1658 (.A(net1660),
    .X(net1658));
 sky130_fd_sc_hd__clkbuf_8 fanout1659 (.A(net1660),
    .X(net1659));
 sky130_fd_sc_hd__clkbuf_8 fanout1660 (.A(net1661),
    .X(net1660));
 sky130_fd_sc_hd__buf_6 fanout1661 (.A(net1662),
    .X(net1661));
 sky130_fd_sc_hd__buf_12 fanout1662 (.A(_03842_),
    .X(net1662));
 sky130_fd_sc_hd__buf_12 fanout1663 (.A(net1667),
    .X(net1663));
 sky130_fd_sc_hd__buf_6 fanout1664 (.A(net1665),
    .X(net1664));
 sky130_fd_sc_hd__buf_6 fanout1665 (.A(net1667),
    .X(net1665));
 sky130_fd_sc_hd__clkbuf_16 fanout1666 (.A(net1667),
    .X(net1666));
 sky130_fd_sc_hd__clkbuf_16 fanout1667 (.A(_03841_),
    .X(net1667));
 sky130_fd_sc_hd__buf_6 fanout1668 (.A(net1669),
    .X(net1668));
 sky130_fd_sc_hd__clkbuf_16 fanout1669 (.A(net1671),
    .X(net1669));
 sky130_fd_sc_hd__buf_12 fanout1670 (.A(net1671),
    .X(net1670));
 sky130_fd_sc_hd__buf_12 fanout1671 (.A(_03840_),
    .X(net1671));
 sky130_fd_sc_hd__buf_12 fanout1672 (.A(net1673),
    .X(net1672));
 sky130_fd_sc_hd__buf_12 fanout1673 (.A(net1674),
    .X(net1673));
 sky130_fd_sc_hd__buf_12 fanout1674 (.A(_03838_),
    .X(net1674));
 sky130_fd_sc_hd__buf_6 fanout1675 (.A(net1676),
    .X(net1675));
 sky130_fd_sc_hd__buf_6 fanout1676 (.A(net1679),
    .X(net1676));
 sky130_fd_sc_hd__clkbuf_8 fanout1677 (.A(net1679),
    .X(net1677));
 sky130_fd_sc_hd__clkbuf_8 fanout1678 (.A(net1679),
    .X(net1678));
 sky130_fd_sc_hd__buf_8 fanout1679 (.A(net1685),
    .X(net1679));
 sky130_fd_sc_hd__buf_6 fanout1680 (.A(net1684),
    .X(net1680));
 sky130_fd_sc_hd__buf_4 fanout1681 (.A(net1684),
    .X(net1681));
 sky130_fd_sc_hd__buf_6 fanout1682 (.A(net1684),
    .X(net1682));
 sky130_fd_sc_hd__buf_6 fanout1683 (.A(net1684),
    .X(net1683));
 sky130_fd_sc_hd__buf_12 fanout1684 (.A(net1685),
    .X(net1684));
 sky130_fd_sc_hd__buf_8 fanout1685 (.A(_03837_),
    .X(net1685));
 sky130_fd_sc_hd__buf_6 fanout1686 (.A(net1687),
    .X(net1686));
 sky130_fd_sc_hd__buf_6 fanout1687 (.A(net1690),
    .X(net1687));
 sky130_fd_sc_hd__buf_6 fanout1688 (.A(net1689),
    .X(net1688));
 sky130_fd_sc_hd__buf_6 fanout1689 (.A(net1690),
    .X(net1689));
 sky130_fd_sc_hd__buf_8 fanout1690 (.A(_03837_),
    .X(net1690));
 sky130_fd_sc_hd__buf_6 fanout1691 (.A(net1695),
    .X(net1691));
 sky130_fd_sc_hd__buf_6 fanout1692 (.A(net1695),
    .X(net1692));
 sky130_fd_sc_hd__buf_2 fanout1693 (.A(net1695),
    .X(net1693));
 sky130_fd_sc_hd__clkbuf_8 fanout1694 (.A(net1695),
    .X(net1694));
 sky130_fd_sc_hd__buf_6 fanout1695 (.A(_03837_),
    .X(net1695));
 sky130_fd_sc_hd__buf_4 fanout1696 (.A(net1697),
    .X(net1696));
 sky130_fd_sc_hd__clkbuf_4 fanout1697 (.A(net1698),
    .X(net1697));
 sky130_fd_sc_hd__buf_4 fanout1698 (.A(_03837_),
    .X(net1698));
 sky130_fd_sc_hd__buf_8 fanout1699 (.A(net1700),
    .X(net1699));
 sky130_fd_sc_hd__buf_12 fanout1700 (.A(net1703),
    .X(net1700));
 sky130_fd_sc_hd__buf_8 fanout1701 (.A(net1702),
    .X(net1701));
 sky130_fd_sc_hd__buf_12 fanout1702 (.A(net1703),
    .X(net1702));
 sky130_fd_sc_hd__buf_12 fanout1703 (.A(_03836_),
    .X(net1703));
 sky130_fd_sc_hd__clkbuf_16 fanout1704 (.A(net1705),
    .X(net1704));
 sky130_fd_sc_hd__buf_12 fanout1705 (.A(_03835_),
    .X(net1705));
 sky130_fd_sc_hd__buf_12 fanout1706 (.A(net1707),
    .X(net1706));
 sky130_fd_sc_hd__buf_12 fanout1707 (.A(_03835_),
    .X(net1707));
 sky130_fd_sc_hd__buf_8 fanout1708 (.A(net1709),
    .X(net1708));
 sky130_fd_sc_hd__buf_8 fanout1709 (.A(net1711),
    .X(net1709));
 sky130_fd_sc_hd__buf_12 fanout1710 (.A(net1711),
    .X(net1710));
 sky130_fd_sc_hd__buf_12 fanout1711 (.A(_03834_),
    .X(net1711));
 sky130_fd_sc_hd__buf_6 fanout1712 (.A(_03829_),
    .X(net1712));
 sky130_fd_sc_hd__buf_8 fanout1713 (.A(_03820_),
    .X(net1713));
 sky130_fd_sc_hd__buf_6 fanout1714 (.A(_03820_),
    .X(net1714));
 sky130_fd_sc_hd__buf_8 fanout1715 (.A(net1716),
    .X(net1715));
 sky130_fd_sc_hd__clkbuf_4 fanout1716 (.A(net1718),
    .X(net1716));
 sky130_fd_sc_hd__buf_8 fanout1717 (.A(net1718),
    .X(net1717));
 sky130_fd_sc_hd__buf_4 fanout1718 (.A(_03820_),
    .X(net1718));
 sky130_fd_sc_hd__buf_12 fanout1719 (.A(net482),
    .X(net1719));
 sky130_fd_sc_hd__buf_4 fanout1720 (.A(\jtag.state[1] ),
    .X(net1720));
 sky130_fd_sc_hd__buf_6 fanout1721 (.A(\jtag.state[0] ),
    .X(net1721));
 sky130_fd_sc_hd__buf_4 fanout1722 (.A(net1723),
    .X(net1722));
 sky130_fd_sc_hd__clkbuf_4 fanout1723 (.A(\jtag.tckRisingEdge ),
    .X(net1723));
 sky130_fd_sc_hd__buf_4 fanout1724 (.A(net1725),
    .X(net1724));
 sky130_fd_sc_hd__buf_6 fanout1725 (.A(net1730),
    .X(net1725));
 sky130_fd_sc_hd__buf_6 fanout1726 (.A(net1730),
    .X(net1726));
 sky130_fd_sc_hd__buf_4 fanout1727 (.A(net1728),
    .X(net1727));
 sky130_fd_sc_hd__clkbuf_4 fanout1728 (.A(net1730),
    .X(net1728));
 sky130_fd_sc_hd__buf_6 fanout1729 (.A(net1730),
    .X(net1729));
 sky130_fd_sc_hd__buf_6 fanout1730 (.A(\core.management_run ),
    .X(net1730));
 sky130_fd_sc_hd__buf_4 fanout1731 (.A(net1733),
    .X(net1731));
 sky130_fd_sc_hd__clkbuf_4 fanout1732 (.A(net1733),
    .X(net1732));
 sky130_fd_sc_hd__clkbuf_4 fanout1733 (.A(\core.management_interruptEnable ),
    .X(net1733));
 sky130_fd_sc_hd__buf_12 fanout1734 (.A(\localMemoryInterface.lastRBankSelect ),
    .X(net1734));
 sky130_fd_sc_hd__buf_4 fanout1735 (.A(\localMemoryInterface.lastRBankSelect ),
    .X(net1735));
 sky130_fd_sc_hd__buf_12 fanout1736 (.A(\localMemoryInterface.lastRBankSelect ),
    .X(net1736));
 sky130_fd_sc_hd__buf_6 fanout1737 (.A(\localMemoryInterface.lastRBankSelect ),
    .X(net1737));
 sky130_fd_sc_hd__buf_6 fanout1738 (.A(net1740),
    .X(net1738));
 sky130_fd_sc_hd__buf_4 fanout1739 (.A(net1740),
    .X(net1739));
 sky130_fd_sc_hd__clkbuf_4 fanout1740 (.A(\localMemoryInterface.wbReadReady ),
    .X(net1740));
 sky130_fd_sc_hd__buf_12 fanout1741 (.A(\localMemoryInterface.lastRWBankSelect ),
    .X(net1741));
 sky130_fd_sc_hd__clkbuf_4 fanout1742 (.A(\localMemoryInterface.lastRWBankSelect ),
    .X(net1742));
 sky130_fd_sc_hd__buf_4 fanout1743 (.A(\localMemoryInterface.lastRWBankSelect ),
    .X(net1743));
 sky130_fd_sc_hd__buf_2 fanout1744 (.A(\localMemoryInterface.lastRWBankSelect ),
    .X(net1744));
 sky130_fd_sc_hd__buf_4 fanout1745 (.A(\memoryController.last_data_enableLocalMemory ),
    .X(net1745));
 sky130_fd_sc_hd__buf_4 fanout1746 (.A(\memoryController.last_instruction_enableLocalMemory ),
    .X(net1746));
 sky130_fd_sc_hd__buf_12 fanout1747 (.A(net457),
    .X(net1747));
 sky130_fd_sc_hd__buf_12 fanout1748 (.A(net476),
    .X(net1748));
 sky130_fd_sc_hd__buf_6 fanout1749 (.A(\core.pipe1_resultRegister[1] ),
    .X(net1749));
 sky130_fd_sc_hd__buf_8 fanout1750 (.A(\core.pipe1_resultRegister[0] ),
    .X(net1750));
 sky130_fd_sc_hd__buf_12 fanout1751 (.A(\core.pipe0_currentInstruction[31] ),
    .X(net1751));
 sky130_fd_sc_hd__buf_12 fanout1752 (.A(\core.pipe0_currentInstruction[30] ),
    .X(net1752));
 sky130_fd_sc_hd__buf_8 fanout1753 (.A(net1754),
    .X(net1753));
 sky130_fd_sc_hd__buf_12 fanout1754 (.A(net1755),
    .X(net1754));
 sky130_fd_sc_hd__buf_12 fanout1755 (.A(\core.pipe0_currentInstruction[24] ),
    .X(net1755));
 sky130_fd_sc_hd__buf_6 fanout1756 (.A(net1757),
    .X(net1756));
 sky130_fd_sc_hd__buf_6 fanout1757 (.A(net1758),
    .X(net1757));
 sky130_fd_sc_hd__clkbuf_4 fanout1758 (.A(net1760),
    .X(net1758));
 sky130_fd_sc_hd__buf_12 fanout1759 (.A(net1760),
    .X(net1759));
 sky130_fd_sc_hd__clkbuf_16 fanout1760 (.A(\core.pipe0_currentInstruction[24] ),
    .X(net1760));
 sky130_fd_sc_hd__buf_12 fanout1761 (.A(net1762),
    .X(net1761));
 sky130_fd_sc_hd__buf_12 fanout1762 (.A(\core.pipe0_currentInstruction[23] ),
    .X(net1762));
 sky130_fd_sc_hd__buf_12 fanout1763 (.A(net1764),
    .X(net1763));
 sky130_fd_sc_hd__buf_12 fanout1764 (.A(net1767),
    .X(net1764));
 sky130_fd_sc_hd__buf_12 fanout1765 (.A(net1766),
    .X(net1765));
 sky130_fd_sc_hd__buf_12 fanout1766 (.A(net1767),
    .X(net1766));
 sky130_fd_sc_hd__clkbuf_16 fanout1767 (.A(\core.pipe0_currentInstruction[22] ),
    .X(net1767));
 sky130_fd_sc_hd__buf_6 fanout1768 (.A(net1771),
    .X(net1768));
 sky130_fd_sc_hd__buf_4 fanout1769 (.A(net1771),
    .X(net1769));
 sky130_fd_sc_hd__buf_6 fanout1770 (.A(net1771),
    .X(net1770));
 sky130_fd_sc_hd__buf_12 fanout1771 (.A(\core.pipe0_currentInstruction[21] ),
    .X(net1771));
 sky130_fd_sc_hd__buf_8 fanout1772 (.A(net1775),
    .X(net1772));
 sky130_fd_sc_hd__buf_6 fanout1773 (.A(net1775),
    .X(net1773));
 sky130_fd_sc_hd__buf_6 fanout1774 (.A(net1775),
    .X(net1774));
 sky130_fd_sc_hd__buf_12 fanout1775 (.A(\core.pipe0_currentInstruction[21] ),
    .X(net1775));
 sky130_fd_sc_hd__buf_12 fanout1776 (.A(\core.pipe0_currentInstruction[20] ),
    .X(net1776));
 sky130_fd_sc_hd__buf_12 fanout1777 (.A(\core.pipe0_currentInstruction[20] ),
    .X(net1777));
 sky130_fd_sc_hd__buf_6 fanout1778 (.A(net1779),
    .X(net1778));
 sky130_fd_sc_hd__clkbuf_16 fanout1779 (.A(net1780),
    .X(net1779));
 sky130_fd_sc_hd__buf_12 fanout1780 (.A(\core.pipe0_currentInstruction[19] ),
    .X(net1780));
 sky130_fd_sc_hd__buf_6 fanout1781 (.A(net1782),
    .X(net1781));
 sky130_fd_sc_hd__buf_12 fanout1782 (.A(net1783),
    .X(net1782));
 sky130_fd_sc_hd__buf_8 fanout1783 (.A(\core.pipe0_currentInstruction[19] ),
    .X(net1783));
 sky130_fd_sc_hd__buf_12 fanout1784 (.A(\core.pipe0_currentInstruction[17] ),
    .X(net1784));
 sky130_fd_sc_hd__buf_12 fanout1785 (.A(net1786),
    .X(net1785));
 sky130_fd_sc_hd__clkbuf_16 fanout1786 (.A(\core.pipe0_currentInstruction[17] ),
    .X(net1786));
 sky130_fd_sc_hd__buf_8 fanout1787 (.A(net1789),
    .X(net1787));
 sky130_fd_sc_hd__buf_6 fanout1788 (.A(net1789),
    .X(net1788));
 sky130_fd_sc_hd__buf_12 fanout1789 (.A(\core.pipe0_currentInstruction[16] ),
    .X(net1789));
 sky130_fd_sc_hd__buf_6 fanout1790 (.A(net1791),
    .X(net1790));
 sky130_fd_sc_hd__buf_12 fanout1791 (.A(net1792),
    .X(net1791));
 sky130_fd_sc_hd__buf_12 fanout1792 (.A(\core.pipe0_currentInstruction[16] ),
    .X(net1792));
 sky130_fd_sc_hd__buf_12 fanout1793 (.A(\core.pipe0_currentInstruction[15] ),
    .X(net1793));
 sky130_fd_sc_hd__buf_12 fanout1794 (.A(\core.pipe0_currentInstruction[14] ),
    .X(net1794));
 sky130_fd_sc_hd__buf_4 fanout1795 (.A(\core.pipe0_currentInstruction[14] ),
    .X(net1795));
 sky130_fd_sc_hd__clkbuf_4 fanout1796 (.A(net1798),
    .X(net1796));
 sky130_fd_sc_hd__clkbuf_2 fanout1797 (.A(net1798),
    .X(net1797));
 sky130_fd_sc_hd__buf_4 fanout1798 (.A(\core.pipe1_operation.currentPipeStall ),
    .X(net1798));
 sky130_fd_sc_hd__buf_8 fanout1799 (.A(\core.csr.currentInstruction[14] ),
    .X(net1799));
 sky130_fd_sc_hd__buf_4 fanout1800 (.A(\core.csr.currentInstruction[13] ),
    .X(net1800));
 sky130_fd_sc_hd__buf_6 fanout1801 (.A(\core.csr.currentInstruction[9] ),
    .X(net1801));
 sky130_fd_sc_hd__clkbuf_4 fanout1802 (.A(net1804),
    .X(net1802));
 sky130_fd_sc_hd__buf_4 fanout1803 (.A(net1804),
    .X(net1803));
 sky130_fd_sc_hd__clkbuf_4 fanout1804 (.A(net1805),
    .X(net1804));
 sky130_fd_sc_hd__clkbuf_8 fanout1805 (.A(net1870),
    .X(net1805));
 sky130_fd_sc_hd__clkbuf_4 fanout1806 (.A(net1809),
    .X(net1806));
 sky130_fd_sc_hd__clkbuf_4 fanout1807 (.A(net1809),
    .X(net1807));
 sky130_fd_sc_hd__clkbuf_2 fanout1808 (.A(net1809),
    .X(net1808));
 sky130_fd_sc_hd__clkbuf_4 fanout1809 (.A(net1810),
    .X(net1809));
 sky130_fd_sc_hd__buf_4 fanout1810 (.A(net1820),
    .X(net1810));
 sky130_fd_sc_hd__clkbuf_4 fanout1811 (.A(net1812),
    .X(net1811));
 sky130_fd_sc_hd__buf_2 fanout1812 (.A(net1813),
    .X(net1812));
 sky130_fd_sc_hd__buf_2 fanout1813 (.A(net1820),
    .X(net1813));
 sky130_fd_sc_hd__buf_4 fanout1814 (.A(net1815),
    .X(net1814));
 sky130_fd_sc_hd__buf_4 fanout1815 (.A(net1820),
    .X(net1815));
 sky130_fd_sc_hd__buf_4 fanout1816 (.A(net1819),
    .X(net1816));
 sky130_fd_sc_hd__buf_2 fanout1817 (.A(net1819),
    .X(net1817));
 sky130_fd_sc_hd__buf_4 fanout1818 (.A(net1819),
    .X(net1818));
 sky130_fd_sc_hd__clkbuf_4 fanout1819 (.A(net1820),
    .X(net1819));
 sky130_fd_sc_hd__clkbuf_8 fanout1820 (.A(net1870),
    .X(net1820));
 sky130_fd_sc_hd__clkbuf_4 fanout1821 (.A(net1823),
    .X(net1821));
 sky130_fd_sc_hd__buf_2 fanout1822 (.A(net1823),
    .X(net1822));
 sky130_fd_sc_hd__buf_6 fanout1823 (.A(net1824),
    .X(net1823));
 sky130_fd_sc_hd__buf_6 fanout1824 (.A(net1870),
    .X(net1824));
 sky130_fd_sc_hd__buf_4 fanout1825 (.A(net1826),
    .X(net1825));
 sky130_fd_sc_hd__clkbuf_4 fanout1826 (.A(net1833),
    .X(net1826));
 sky130_fd_sc_hd__buf_4 fanout1827 (.A(net1833),
    .X(net1827));
 sky130_fd_sc_hd__buf_4 fanout1828 (.A(net1833),
    .X(net1828));
 sky130_fd_sc_hd__buf_4 fanout1829 (.A(net1832),
    .X(net1829));
 sky130_fd_sc_hd__buf_4 fanout1830 (.A(net1832),
    .X(net1830));
 sky130_fd_sc_hd__buf_4 fanout1831 (.A(net1832),
    .X(net1831));
 sky130_fd_sc_hd__clkbuf_4 fanout1832 (.A(net1833),
    .X(net1832));
 sky130_fd_sc_hd__clkbuf_4 fanout1833 (.A(net1870),
    .X(net1833));
 sky130_fd_sc_hd__buf_4 fanout1834 (.A(net1837),
    .X(net1834));
 sky130_fd_sc_hd__buf_2 fanout1835 (.A(net1837),
    .X(net1835));
 sky130_fd_sc_hd__buf_4 fanout1836 (.A(net1837),
    .X(net1836));
 sky130_fd_sc_hd__buf_4 fanout1837 (.A(net1855),
    .X(net1837));
 sky130_fd_sc_hd__buf_4 fanout1838 (.A(net1840),
    .X(net1838));
 sky130_fd_sc_hd__buf_4 fanout1839 (.A(net1840),
    .X(net1839));
 sky130_fd_sc_hd__buf_2 fanout1840 (.A(net1843),
    .X(net1840));
 sky130_fd_sc_hd__buf_4 fanout1841 (.A(net1842),
    .X(net1841));
 sky130_fd_sc_hd__clkbuf_4 fanout1842 (.A(net1843),
    .X(net1842));
 sky130_fd_sc_hd__clkbuf_8 fanout1843 (.A(net1855),
    .X(net1843));
 sky130_fd_sc_hd__buf_4 fanout1844 (.A(net1846),
    .X(net1844));
 sky130_fd_sc_hd__buf_4 fanout1845 (.A(net1846),
    .X(net1845));
 sky130_fd_sc_hd__buf_4 fanout1846 (.A(net1855),
    .X(net1846));
 sky130_fd_sc_hd__buf_4 fanout1847 (.A(net1849),
    .X(net1847));
 sky130_fd_sc_hd__buf_4 fanout1848 (.A(net1849),
    .X(net1848));
 sky130_fd_sc_hd__buf_4 fanout1849 (.A(net1855),
    .X(net1849));
 sky130_fd_sc_hd__buf_4 fanout1850 (.A(net1853),
    .X(net1850));
 sky130_fd_sc_hd__clkbuf_2 fanout1851 (.A(net1853),
    .X(net1851));
 sky130_fd_sc_hd__clkbuf_4 fanout1852 (.A(net1853),
    .X(net1852));
 sky130_fd_sc_hd__buf_2 fanout1853 (.A(net1854),
    .X(net1853));
 sky130_fd_sc_hd__buf_4 fanout1854 (.A(net1855),
    .X(net1854));
 sky130_fd_sc_hd__buf_6 fanout1855 (.A(net1870),
    .X(net1855));
 sky130_fd_sc_hd__buf_4 fanout1856 (.A(net1863),
    .X(net1856));
 sky130_fd_sc_hd__buf_4 fanout1857 (.A(net1863),
    .X(net1857));
 sky130_fd_sc_hd__buf_4 fanout1858 (.A(net1863),
    .X(net1858));
 sky130_fd_sc_hd__buf_4 fanout1859 (.A(net1863),
    .X(net1859));
 sky130_fd_sc_hd__clkbuf_2 fanout1860 (.A(net1863),
    .X(net1860));
 sky130_fd_sc_hd__buf_4 fanout1861 (.A(net1862),
    .X(net1861));
 sky130_fd_sc_hd__clkbuf_4 fanout1862 (.A(net1863),
    .X(net1862));
 sky130_fd_sc_hd__buf_4 fanout1863 (.A(net1870),
    .X(net1863));
 sky130_fd_sc_hd__buf_4 fanout1864 (.A(net1865),
    .X(net1864));
 sky130_fd_sc_hd__buf_4 fanout1865 (.A(net1869),
    .X(net1865));
 sky130_fd_sc_hd__buf_4 fanout1866 (.A(net1867),
    .X(net1866));
 sky130_fd_sc_hd__buf_2 fanout1867 (.A(net1868),
    .X(net1867));
 sky130_fd_sc_hd__clkbuf_4 fanout1868 (.A(net1869),
    .X(net1868));
 sky130_fd_sc_hd__clkbuf_4 fanout1869 (.A(net1870),
    .X(net1869));
 sky130_fd_sc_hd__buf_12 fanout1870 (.A(_03851_),
    .X(net1870));
 sky130_fd_sc_hd__clkbuf_8 fanout1871 (.A(net1873),
    .X(net1871));
 sky130_fd_sc_hd__buf_4 fanout1872 (.A(net1873),
    .X(net1872));
 sky130_fd_sc_hd__buf_8 fanout1873 (.A(net1874),
    .X(net1873));
 sky130_fd_sc_hd__buf_8 fanout1874 (.A(net1906),
    .X(net1874));
 sky130_fd_sc_hd__buf_6 fanout1875 (.A(net1876),
    .X(net1875));
 sky130_fd_sc_hd__buf_4 fanout1876 (.A(net1879),
    .X(net1876));
 sky130_fd_sc_hd__buf_6 fanout1877 (.A(net1879),
    .X(net1877));
 sky130_fd_sc_hd__clkbuf_4 fanout1878 (.A(net1879),
    .X(net1878));
 sky130_fd_sc_hd__buf_12 fanout1879 (.A(net1906),
    .X(net1879));
 sky130_fd_sc_hd__clkbuf_8 fanout1880 (.A(net1881),
    .X(net1880));
 sky130_fd_sc_hd__buf_6 fanout1881 (.A(net1905),
    .X(net1881));
 sky130_fd_sc_hd__buf_4 fanout1882 (.A(net1883),
    .X(net1882));
 sky130_fd_sc_hd__buf_4 fanout1883 (.A(net1905),
    .X(net1883));
 sky130_fd_sc_hd__buf_2 fanout1884 (.A(net1905),
    .X(net1884));
 sky130_fd_sc_hd__buf_4 fanout1885 (.A(net1905),
    .X(net1885));
 sky130_fd_sc_hd__buf_6 fanout1886 (.A(net1905),
    .X(net1886));
 sky130_fd_sc_hd__buf_4 fanout1887 (.A(net1888),
    .X(net1887));
 sky130_fd_sc_hd__buf_4 fanout1888 (.A(net1904),
    .X(net1888));
 sky130_fd_sc_hd__buf_4 fanout1889 (.A(net1890),
    .X(net1889));
 sky130_fd_sc_hd__buf_2 fanout1890 (.A(net1891),
    .X(net1890));
 sky130_fd_sc_hd__buf_2 fanout1891 (.A(net1904),
    .X(net1891));
 sky130_fd_sc_hd__buf_4 fanout1892 (.A(net1893),
    .X(net1892));
 sky130_fd_sc_hd__buf_4 fanout1893 (.A(net1897),
    .X(net1893));
 sky130_fd_sc_hd__buf_4 fanout1894 (.A(net1896),
    .X(net1894));
 sky130_fd_sc_hd__buf_4 fanout1895 (.A(net1896),
    .X(net1895));
 sky130_fd_sc_hd__clkbuf_4 fanout1896 (.A(net1897),
    .X(net1896));
 sky130_fd_sc_hd__clkbuf_4 fanout1897 (.A(net1904),
    .X(net1897));
 sky130_fd_sc_hd__buf_4 fanout1898 (.A(net1901),
    .X(net1898));
 sky130_fd_sc_hd__buf_4 fanout1899 (.A(net1901),
    .X(net1899));
 sky130_fd_sc_hd__buf_2 fanout1900 (.A(net1901),
    .X(net1900));
 sky130_fd_sc_hd__clkbuf_4 fanout1901 (.A(net1903),
    .X(net1901));
 sky130_fd_sc_hd__buf_6 fanout1902 (.A(net1903),
    .X(net1902));
 sky130_fd_sc_hd__clkbuf_4 fanout1903 (.A(net1904),
    .X(net1903));
 sky130_fd_sc_hd__clkbuf_8 fanout1904 (.A(net1905),
    .X(net1904));
 sky130_fd_sc_hd__buf_8 fanout1905 (.A(net1906),
    .X(net1905));
 sky130_fd_sc_hd__buf_12 fanout1906 (.A(net284),
    .X(net1906));
 sky130_fd_sc_hd__clkbuf_4 fanout1907 (.A(net1908),
    .X(net1907));
 sky130_fd_sc_hd__clkbuf_2 fanout1908 (.A(net1910),
    .X(net1908));
 sky130_fd_sc_hd__buf_4 fanout1909 (.A(net1910),
    .X(net1909));
 sky130_fd_sc_hd__buf_4 fanout1910 (.A(net205),
    .X(net1910));
 sky130_fd_sc_hd__buf_12 fanout488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__buf_12 fanout489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__buf_12 fanout490 (.A(net492),
    .X(net490));
 sky130_fd_sc_hd__buf_4 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_16 fanout492 (.A(_01896_),
    .X(net492));
 sky130_fd_sc_hd__buf_4 fanout493 (.A(_01896_),
    .X(net493));
 sky130_fd_sc_hd__buf_6 fanout494 (.A(_01896_),
    .X(net494));
 sky130_fd_sc_hd__buf_6 fanout495 (.A(net499),
    .X(net495));
 sky130_fd_sc_hd__buf_6 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_4 fanout497 (.A(net499),
    .X(net497));
 sky130_fd_sc_hd__buf_6 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_4 fanout499 (.A(_06829_),
    .X(net499));
 sky130_fd_sc_hd__buf_8 fanout500 (.A(_06692_),
    .X(net500));
 sky130_fd_sc_hd__buf_6 fanout501 (.A(net503),
    .X(net501));
 sky130_fd_sc_hd__buf_4 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__buf_6 fanout503 (.A(net504),
    .X(net503));
 sky130_fd_sc_hd__buf_6 fanout504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__buf_8 fanout505 (.A(_06692_),
    .X(net505));
 sky130_fd_sc_hd__buf_4 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_8 fanout507 (.A(net513),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_2 fanout508 (.A(net513),
    .X(net508));
 sky130_fd_sc_hd__buf_6 fanout509 (.A(net513),
    .X(net509));
 sky130_fd_sc_hd__buf_4 fanout510 (.A(net511),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_4 fanout511 (.A(net513),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_8 fanout512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__buf_6 fanout513 (.A(_03631_),
    .X(net513));
 sky130_fd_sc_hd__buf_4 fanout514 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_8 fanout515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__buf_6 fanout516 (.A(_03527_),
    .X(net516));
 sky130_fd_sc_hd__buf_4 fanout517 (.A(net520),
    .X(net517));
 sky130_fd_sc_hd__buf_4 fanout518 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_8 fanout519 (.A(net520),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_4 fanout520 (.A(_03527_),
    .X(net520));
 sky130_fd_sc_hd__buf_6 fanout521 (.A(net522),
    .X(net521));
 sky130_fd_sc_hd__buf_4 fanout522 (.A(_02263_),
    .X(net522));
 sky130_fd_sc_hd__buf_6 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_6 fanout524 (.A(_02263_),
    .X(net524));
 sky130_fd_sc_hd__buf_4 fanout525 (.A(net531),
    .X(net525));
 sky130_fd_sc_hd__buf_4 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_8 fanout527 (.A(_06710_),
    .X(net527));
 sky130_fd_sc_hd__buf_4 fanout528 (.A(net530),
    .X(net528));
 sky130_fd_sc_hd__buf_2 fanout529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__buf_4 fanout530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__buf_8 fanout531 (.A(_06710_),
    .X(net531));
 sky130_fd_sc_hd__buf_8 fanout532 (.A(_06652_),
    .X(net532));
 sky130_fd_sc_hd__buf_4 fanout533 (.A(net536),
    .X(net533));
 sky130_fd_sc_hd__buf_6 fanout534 (.A(net536),
    .X(net534));
 sky130_fd_sc_hd__buf_2 fanout535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_6 fanout536 (.A(_03459_),
    .X(net536));
 sky130_fd_sc_hd__buf_6 fanout537 (.A(net540),
    .X(net537));
 sky130_fd_sc_hd__buf_6 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_4 fanout539 (.A(net540),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_8 fanout540 (.A(_02262_),
    .X(net540));
 sky130_fd_sc_hd__buf_4 fanout541 (.A(net543),
    .X(net541));
 sky130_fd_sc_hd__buf_4 fanout542 (.A(net543),
    .X(net542));
 sky130_fd_sc_hd__buf_6 fanout543 (.A(net548),
    .X(net543));
 sky130_fd_sc_hd__buf_4 fanout544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_8 fanout545 (.A(net548),
    .X(net545));
 sky130_fd_sc_hd__buf_4 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__buf_6 fanout547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__buf_4 fanout548 (.A(_02259_),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_8 fanout549 (.A(net550),
    .X(net549));
 sky130_fd_sc_hd__buf_6 fanout550 (.A(net552),
    .X(net550));
 sky130_fd_sc_hd__buf_8 fanout551 (.A(net552),
    .X(net551));
 sky130_fd_sc_hd__buf_8 fanout552 (.A(_02258_),
    .X(net552));
 sky130_fd_sc_hd__buf_4 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__buf_6 fanout554 (.A(_02258_),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_8 fanout555 (.A(_02258_),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_4 fanout556 (.A(_02258_),
    .X(net556));
 sky130_fd_sc_hd__buf_4 fanout557 (.A(net558),
    .X(net557));
 sky130_fd_sc_hd__buf_6 fanout558 (.A(_02666_),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_8 fanout559 (.A(net561),
    .X(net559));
 sky130_fd_sc_hd__buf_2 fanout560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__buf_4 fanout561 (.A(_02248_),
    .X(net561));
 sky130_fd_sc_hd__buf_6 fanout562 (.A(net564),
    .X(net562));
 sky130_fd_sc_hd__buf_2 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_8 fanout564 (.A(_02248_),
    .X(net564));
 sky130_fd_sc_hd__buf_4 fanout565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__buf_6 fanout566 (.A(_02268_),
    .X(net566));
 sky130_fd_sc_hd__buf_8 fanout567 (.A(_02260_),
    .X(net567));
 sky130_fd_sc_hd__buf_8 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__buf_12 fanout569 (.A(_02249_),
    .X(net569));
 sky130_fd_sc_hd__buf_8 fanout570 (.A(_02241_),
    .X(net570));
 sky130_fd_sc_hd__buf_6 fanout571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__buf_6 fanout572 (.A(_02241_),
    .X(net572));
 sky130_fd_sc_hd__buf_4 fanout573 (.A(net574),
    .X(net573));
 sky130_fd_sc_hd__buf_4 fanout574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_8 fanout575 (.A(_03068_),
    .X(net575));
 sky130_fd_sc_hd__buf_4 fanout576 (.A(net578),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_2 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__buf_2 fanout578 (.A(_07072_),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_4 fanout579 (.A(net580),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_4 fanout580 (.A(_07072_),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_4 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 fanout582 (.A(_07072_),
    .X(net582));
 sky130_fd_sc_hd__buf_4 fanout583 (.A(_07072_),
    .X(net583));
 sky130_fd_sc_hd__buf_4 fanout584 (.A(_06856_),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_4 fanout585 (.A(_06856_),
    .X(net585));
 sky130_fd_sc_hd__buf_4 fanout586 (.A(net587),
    .X(net586));
 sky130_fd_sc_hd__buf_4 fanout587 (.A(_06856_),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_4 fanout588 (.A(net591),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_4 fanout589 (.A(net591),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_2 fanout590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__buf_4 fanout591 (.A(_06855_),
    .X(net591));
 sky130_fd_sc_hd__buf_4 fanout592 (.A(net594),
    .X(net592));
 sky130_fd_sc_hd__buf_4 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_4 fanout594 (.A(net595),
    .X(net594));
 sky130_fd_sc_hd__buf_4 fanout595 (.A(net598),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_16 fanout596 (.A(net598),
    .X(net596));
 sky130_fd_sc_hd__buf_2 fanout597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_16 fanout598 (.A(_06685_),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_4 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__buf_4 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__buf_8 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_8 fanout602 (.A(_06684_),
    .X(net602));
 sky130_fd_sc_hd__buf_4 fanout603 (.A(net606),
    .X(net603));
 sky130_fd_sc_hd__buf_6 fanout604 (.A(net606),
    .X(net604));
 sky130_fd_sc_hd__buf_2 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__buf_4 fanout606 (.A(_02216_),
    .X(net606));
 sky130_fd_sc_hd__buf_8 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__buf_8 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__buf_6 fanout609 (.A(_07273_),
    .X(net609));
 sky130_fd_sc_hd__buf_12 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__buf_8 fanout611 (.A(net612),
    .X(net611));
 sky130_fd_sc_hd__buf_8 fanout612 (.A(net613),
    .X(net612));
 sky130_fd_sc_hd__buf_8 fanout613 (.A(_06642_),
    .X(net613));
 sky130_fd_sc_hd__buf_4 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__buf_4 fanout615 (.A(net617),
    .X(net615));
 sky130_fd_sc_hd__buf_6 fanout616 (.A(net617),
    .X(net616));
 sky130_fd_sc_hd__buf_4 fanout617 (.A(_03767_),
    .X(net617));
 sky130_fd_sc_hd__buf_4 fanout618 (.A(net619),
    .X(net618));
 sky130_fd_sc_hd__buf_6 fanout619 (.A(net621),
    .X(net619));
 sky130_fd_sc_hd__buf_6 fanout620 (.A(net621),
    .X(net620));
 sky130_fd_sc_hd__buf_6 fanout621 (.A(_03458_),
    .X(net621));
 sky130_fd_sc_hd__buf_6 fanout622 (.A(net623),
    .X(net622));
 sky130_fd_sc_hd__buf_6 fanout623 (.A(_03384_),
    .X(net623));
 sky130_fd_sc_hd__buf_4 fanout624 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__buf_4 fanout625 (.A(_03384_),
    .X(net625));
 sky130_fd_sc_hd__buf_4 fanout626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_4 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_8 fanout628 (.A(_03279_),
    .X(net628));
 sky130_fd_sc_hd__buf_6 fanout629 (.A(_03279_),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_4 fanout630 (.A(_03279_),
    .X(net630));
 sky130_fd_sc_hd__buf_4 fanout631 (.A(_07446_),
    .X(net631));
 sky130_fd_sc_hd__buf_2 fanout632 (.A(_07446_),
    .X(net632));
 sky130_fd_sc_hd__buf_12 fanout633 (.A(_06641_),
    .X(net633));
 sky130_fd_sc_hd__buf_8 fanout634 (.A(net635),
    .X(net634));
 sky130_fd_sc_hd__buf_6 fanout635 (.A(_06640_),
    .X(net635));
 sky130_fd_sc_hd__buf_4 fanout636 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__buf_4 fanout637 (.A(_03765_),
    .X(net637));
 sky130_fd_sc_hd__buf_8 fanout638 (.A(_03592_),
    .X(net638));
 sky130_fd_sc_hd__buf_6 fanout639 (.A(_03592_),
    .X(net639));
 sky130_fd_sc_hd__buf_6 fanout640 (.A(net641),
    .X(net640));
 sky130_fd_sc_hd__buf_4 fanout641 (.A(_03592_),
    .X(net641));
 sky130_fd_sc_hd__buf_6 fanout642 (.A(net643),
    .X(net642));
 sky130_fd_sc_hd__buf_6 fanout643 (.A(_03422_),
    .X(net643));
 sky130_fd_sc_hd__buf_4 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__buf_4 fanout645 (.A(_03422_),
    .X(net645));
 sky130_fd_sc_hd__buf_4 fanout646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__buf_4 fanout647 (.A(_03421_),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_4 fanout648 (.A(net649),
    .X(net648));
 sky130_fd_sc_hd__buf_2 fanout649 (.A(_03421_),
    .X(net649));
 sky130_fd_sc_hd__buf_4 fanout650 (.A(net651),
    .X(net650));
 sky130_fd_sc_hd__buf_4 fanout651 (.A(_03386_),
    .X(net651));
 sky130_fd_sc_hd__buf_4 fanout652 (.A(net653),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_4 fanout653 (.A(_03386_),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_4 fanout654 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__buf_4 fanout655 (.A(net657),
    .X(net655));
 sky130_fd_sc_hd__buf_6 fanout656 (.A(net657),
    .X(net656));
 sky130_fd_sc_hd__buf_4 fanout657 (.A(_07282_),
    .X(net657));
 sky130_fd_sc_hd__buf_4 fanout658 (.A(net659),
    .X(net658));
 sky130_fd_sc_hd__buf_4 fanout659 (.A(net660),
    .X(net659));
 sky130_fd_sc_hd__buf_6 fanout660 (.A(_07271_),
    .X(net660));
 sky130_fd_sc_hd__buf_4 fanout661 (.A(net662),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_8 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__clkbuf_8 fanout663 (.A(_07264_),
    .X(net663));
 sky130_fd_sc_hd__buf_4 fanout664 (.A(net665),
    .X(net664));
 sky130_fd_sc_hd__buf_4 fanout665 (.A(net666),
    .X(net665));
 sky130_fd_sc_hd__buf_6 fanout666 (.A(_07257_),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_16 fanout667 (.A(net669),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_8 fanout668 (.A(net669),
    .X(net668));
 sky130_fd_sc_hd__buf_12 fanout669 (.A(_06638_),
    .X(net669));
 sky130_fd_sc_hd__buf_8 fanout670 (.A(net671),
    .X(net670));
 sky130_fd_sc_hd__buf_4 fanout671 (.A(_06637_),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_16 fanout672 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__buf_4 fanout673 (.A(net675),
    .X(net673));
 sky130_fd_sc_hd__buf_8 fanout674 (.A(net675),
    .X(net674));
 sky130_fd_sc_hd__buf_4 fanout675 (.A(_01923_),
    .X(net675));
 sky130_fd_sc_hd__buf_6 fanout676 (.A(net677),
    .X(net676));
 sky130_fd_sc_hd__buf_6 fanout677 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__buf_6 fanout678 (.A(_07268_),
    .X(net678));
 sky130_fd_sc_hd__buf_8 fanout679 (.A(net680),
    .X(net679));
 sky130_fd_sc_hd__buf_8 fanout680 (.A(net681),
    .X(net680));
 sky130_fd_sc_hd__buf_6 fanout681 (.A(_07267_),
    .X(net681));
 sky130_fd_sc_hd__buf_6 fanout682 (.A(net683),
    .X(net682));
 sky130_fd_sc_hd__buf_6 fanout683 (.A(net684),
    .X(net683));
 sky130_fd_sc_hd__buf_6 fanout684 (.A(_07266_),
    .X(net684));
 sky130_fd_sc_hd__buf_4 fanout685 (.A(net686),
    .X(net685));
 sky130_fd_sc_hd__buf_4 fanout686 (.A(net687),
    .X(net686));
 sky130_fd_sc_hd__buf_6 fanout687 (.A(_07261_),
    .X(net687));
 sky130_fd_sc_hd__buf_4 fanout688 (.A(net689),
    .X(net688));
 sky130_fd_sc_hd__buf_4 fanout689 (.A(net690),
    .X(net689));
 sky130_fd_sc_hd__buf_6 fanout690 (.A(_07260_),
    .X(net690));
 sky130_fd_sc_hd__buf_4 fanout691 (.A(net692),
    .X(net691));
 sky130_fd_sc_hd__buf_4 fanout692 (.A(net693),
    .X(net692));
 sky130_fd_sc_hd__buf_6 fanout693 (.A(_07259_),
    .X(net693));
 sky130_fd_sc_hd__buf_6 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__buf_4 fanout695 (.A(net696),
    .X(net695));
 sky130_fd_sc_hd__buf_6 fanout696 (.A(_07258_),
    .X(net696));
 sky130_fd_sc_hd__buf_4 fanout697 (.A(_07247_),
    .X(net697));
 sky130_fd_sc_hd__buf_2 fanout698 (.A(_07247_),
    .X(net698));
 sky130_fd_sc_hd__buf_4 fanout699 (.A(_07247_),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_4 fanout700 (.A(_07247_),
    .X(net700));
 sky130_fd_sc_hd__buf_4 fanout701 (.A(_07246_),
    .X(net701));
 sky130_fd_sc_hd__buf_2 fanout702 (.A(_07246_),
    .X(net702));
 sky130_fd_sc_hd__buf_4 fanout703 (.A(_07246_),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_4 fanout704 (.A(_07246_),
    .X(net704));
 sky130_fd_sc_hd__buf_6 fanout705 (.A(_07245_),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_4 fanout706 (.A(_07245_),
    .X(net706));
 sky130_fd_sc_hd__buf_6 fanout707 (.A(_07245_),
    .X(net707));
 sky130_fd_sc_hd__buf_2 fanout708 (.A(_07245_),
    .X(net708));
 sky130_fd_sc_hd__buf_8 fanout709 (.A(net712),
    .X(net709));
 sky130_fd_sc_hd__buf_4 fanout710 (.A(net712),
    .X(net710));
 sky130_fd_sc_hd__buf_6 fanout711 (.A(net712),
    .X(net711));
 sky130_fd_sc_hd__buf_4 fanout712 (.A(_07244_),
    .X(net712));
 sky130_fd_sc_hd__buf_4 fanout713 (.A(net716),
    .X(net713));
 sky130_fd_sc_hd__buf_4 fanout714 (.A(net716),
    .X(net714));
 sky130_fd_sc_hd__buf_4 fanout715 (.A(net716),
    .X(net715));
 sky130_fd_sc_hd__buf_4 fanout716 (.A(_07243_),
    .X(net716));
 sky130_fd_sc_hd__buf_8 fanout717 (.A(net719),
    .X(net717));
 sky130_fd_sc_hd__buf_4 fanout718 (.A(net719),
    .X(net718));
 sky130_fd_sc_hd__buf_8 fanout719 (.A(_07234_),
    .X(net719));
 sky130_fd_sc_hd__buf_4 fanout720 (.A(_07199_),
    .X(net720));
 sky130_fd_sc_hd__buf_4 fanout721 (.A(_07199_),
    .X(net721));
 sky130_fd_sc_hd__buf_6 fanout722 (.A(_07199_),
    .X(net722));
 sky130_fd_sc_hd__buf_2 fanout723 (.A(_07199_),
    .X(net723));
 sky130_fd_sc_hd__buf_4 fanout724 (.A(_07197_),
    .X(net724));
 sky130_fd_sc_hd__buf_4 fanout725 (.A(_07197_),
    .X(net725));
 sky130_fd_sc_hd__buf_6 fanout726 (.A(_07197_),
    .X(net726));
 sky130_fd_sc_hd__buf_2 fanout727 (.A(_07197_),
    .X(net727));
 sky130_fd_sc_hd__buf_4 fanout728 (.A(net730),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_4 fanout729 (.A(net730),
    .X(net729));
 sky130_fd_sc_hd__buf_2 fanout730 (.A(_06439_),
    .X(net730));
 sky130_fd_sc_hd__buf_4 fanout731 (.A(_06439_),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_4 fanout732 (.A(net734),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_4 fanout733 (.A(net734),
    .X(net733));
 sky130_fd_sc_hd__buf_2 fanout734 (.A(_06363_),
    .X(net734));
 sky130_fd_sc_hd__buf_4 fanout735 (.A(_06363_),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_4 fanout736 (.A(net737),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_4 fanout737 (.A(net739),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_4 fanout738 (.A(net739),
    .X(net738));
 sky130_fd_sc_hd__buf_2 fanout739 (.A(_06287_),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_4 fanout740 (.A(net741),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_4 fanout741 (.A(net743),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_4 fanout742 (.A(net743),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_8 fanout743 (.A(_06211_),
    .X(net743));
 sky130_fd_sc_hd__buf_4 fanout744 (.A(net745),
    .X(net744));
 sky130_fd_sc_hd__buf_4 fanout745 (.A(_04935_),
    .X(net745));
 sky130_fd_sc_hd__buf_4 fanout746 (.A(net747),
    .X(net746));
 sky130_fd_sc_hd__buf_4 fanout747 (.A(net748),
    .X(net747));
 sky130_fd_sc_hd__buf_6 fanout748 (.A(_04767_),
    .X(net748));
 sky130_fd_sc_hd__buf_4 fanout749 (.A(net751),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_4 fanout750 (.A(net751),
    .X(net750));
 sky130_fd_sc_hd__buf_4 fanout751 (.A(_04766_),
    .X(net751));
 sky130_fd_sc_hd__buf_4 fanout752 (.A(net754),
    .X(net752));
 sky130_fd_sc_hd__buf_6 fanout753 (.A(net754),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_4 fanout754 (.A(_04687_),
    .X(net754));
 sky130_fd_sc_hd__buf_6 fanout755 (.A(net756),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_4 fanout756 (.A(_04686_),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_4 fanout757 (.A(net758),
    .X(net757));
 sky130_fd_sc_hd__buf_6 fanout758 (.A(_04148_),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_4 fanout759 (.A(net760),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_4 fanout760 (.A(_04148_),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_4 fanout761 (.A(net762),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_4 fanout762 (.A(net763),
    .X(net762));
 sky130_fd_sc_hd__buf_2 fanout763 (.A(_04042_),
    .X(net763));
 sky130_fd_sc_hd__buf_4 fanout764 (.A(_04042_),
    .X(net764));
 sky130_fd_sc_hd__buf_12 fanout765 (.A(net768),
    .X(net765));
 sky130_fd_sc_hd__buf_12 fanout766 (.A(net768),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_16 fanout767 (.A(net768),
    .X(net767));
 sky130_fd_sc_hd__buf_12 fanout768 (.A(_03805_),
    .X(net768));
 sky130_fd_sc_hd__buf_12 fanout769 (.A(_03804_),
    .X(net769));
 sky130_fd_sc_hd__buf_6 fanout770 (.A(_03804_),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_16 fanout771 (.A(net772),
    .X(net771));
 sky130_fd_sc_hd__buf_12 fanout772 (.A(_03804_),
    .X(net772));
 sky130_fd_sc_hd__buf_12 fanout773 (.A(_03803_),
    .X(net773));
 sky130_fd_sc_hd__buf_6 fanout774 (.A(_03803_),
    .X(net774));
 sky130_fd_sc_hd__buf_12 fanout775 (.A(net776),
    .X(net775));
 sky130_fd_sc_hd__buf_12 fanout776 (.A(_03803_),
    .X(net776));
 sky130_fd_sc_hd__buf_12 fanout777 (.A(net780),
    .X(net777));
 sky130_fd_sc_hd__buf_12 fanout778 (.A(net779),
    .X(net778));
 sky130_fd_sc_hd__buf_12 fanout779 (.A(net780),
    .X(net779));
 sky130_fd_sc_hd__buf_8 fanout780 (.A(_03128_),
    .X(net780));
 sky130_fd_sc_hd__buf_12 fanout781 (.A(net784),
    .X(net781));
 sky130_fd_sc_hd__buf_12 fanout782 (.A(net783),
    .X(net782));
 sky130_fd_sc_hd__buf_12 fanout783 (.A(net784),
    .X(net783));
 sky130_fd_sc_hd__buf_8 fanout784 (.A(_03127_),
    .X(net784));
 sky130_fd_sc_hd__buf_12 fanout785 (.A(_03126_),
    .X(net785));
 sky130_fd_sc_hd__buf_6 fanout786 (.A(_03126_),
    .X(net786));
 sky130_fd_sc_hd__buf_12 fanout787 (.A(net788),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_16 fanout788 (.A(_03126_),
    .X(net788));
 sky130_fd_sc_hd__buf_12 fanout789 (.A(_03125_),
    .X(net789));
 sky130_fd_sc_hd__buf_6 fanout790 (.A(_03125_),
    .X(net790));
 sky130_fd_sc_hd__buf_12 fanout791 (.A(net792),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_16 fanout792 (.A(_03125_),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_16 fanout793 (.A(net794),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_16 fanout794 (.A(_03119_),
    .X(net794));
 sky130_fd_sc_hd__buf_12 fanout795 (.A(net796),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_16 fanout796 (.A(_03119_),
    .X(net796));
 sky130_fd_sc_hd__buf_12 fanout797 (.A(net800),
    .X(net797));
 sky130_fd_sc_hd__buf_12 fanout798 (.A(net800),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_16 fanout799 (.A(net800),
    .X(net799));
 sky130_fd_sc_hd__buf_12 fanout800 (.A(_03118_),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_16 fanout801 (.A(net804),
    .X(net801));
 sky130_fd_sc_hd__buf_12 fanout802 (.A(net803),
    .X(net802));
 sky130_fd_sc_hd__buf_12 fanout803 (.A(net804),
    .X(net803));
 sky130_fd_sc_hd__buf_12 fanout804 (.A(_03114_),
    .X(net804));
 sky130_fd_sc_hd__buf_12 fanout805 (.A(net808),
    .X(net805));
 sky130_fd_sc_hd__buf_12 fanout806 (.A(net808),
    .X(net806));
 sky130_fd_sc_hd__buf_8 fanout807 (.A(net808),
    .X(net807));
 sky130_fd_sc_hd__buf_12 fanout808 (.A(_02907_),
    .X(net808));
 sky130_fd_sc_hd__buf_12 fanout809 (.A(_08769_),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_8 fanout810 (.A(_08769_),
    .X(net810));
 sky130_fd_sc_hd__buf_12 fanout811 (.A(net812),
    .X(net811));
 sky130_fd_sc_hd__buf_12 fanout812 (.A(_08769_),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_16 fanout813 (.A(net814),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_16 fanout814 (.A(_08767_),
    .X(net814));
 sky130_fd_sc_hd__buf_12 fanout815 (.A(net816),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_16 fanout816 (.A(_08767_),
    .X(net816));
 sky130_fd_sc_hd__buf_12 fanout817 (.A(net820),
    .X(net817));
 sky130_fd_sc_hd__buf_12 fanout818 (.A(net820),
    .X(net818));
 sky130_fd_sc_hd__buf_8 fanout819 (.A(net820),
    .X(net819));
 sky130_fd_sc_hd__buf_12 fanout820 (.A(_08764_),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_16 fanout821 (.A(net824),
    .X(net821));
 sky130_fd_sc_hd__buf_12 fanout822 (.A(net823),
    .X(net822));
 sky130_fd_sc_hd__buf_12 fanout823 (.A(net824),
    .X(net823));
 sky130_fd_sc_hd__buf_12 fanout824 (.A(_08762_),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_8 fanout825 (.A(_07464_),
    .X(net825));
 sky130_fd_sc_hd__buf_12 fanout826 (.A(_06854_),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_8 fanout827 (.A(_06854_),
    .X(net827));
 sky130_fd_sc_hd__buf_12 fanout828 (.A(net829),
    .X(net828));
 sky130_fd_sc_hd__buf_12 fanout829 (.A(_06854_),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_4 fanout830 (.A(net833),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_4 fanout831 (.A(net832),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_4 fanout832 (.A(net833),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_2 fanout833 (.A(_06132_),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_4 fanout834 (.A(net835),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_4 fanout835 (.A(net837),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_2 fanout836 (.A(net837),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_4 fanout837 (.A(_06055_),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_4 fanout838 (.A(net840),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 fanout839 (.A(net840),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_4 fanout840 (.A(_05977_),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_8 fanout841 (.A(_05977_),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_4 fanout842 (.A(net843),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_4 fanout843 (.A(net844),
    .X(net843));
 sky130_fd_sc_hd__buf_4 fanout844 (.A(net845),
    .X(net844));
 sky130_fd_sc_hd__buf_4 fanout845 (.A(_05901_),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_4 fanout846 (.A(net847),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_4 fanout847 (.A(net849),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_4 fanout848 (.A(net849),
    .X(net848));
 sky130_fd_sc_hd__buf_4 fanout849 (.A(_05825_),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_4 fanout850 (.A(net854),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_2 fanout851 (.A(net854),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_4 fanout852 (.A(net854),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_2 fanout853 (.A(net854),
    .X(net853));
 sky130_fd_sc_hd__buf_6 fanout854 (.A(_05748_),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_4 fanout855 (.A(net859),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_2 fanout856 (.A(net859),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_4 fanout857 (.A(net859),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_2 fanout858 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__buf_4 fanout859 (.A(_05670_),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_4 fanout860 (.A(net861),
    .X(net860));
 sky130_fd_sc_hd__buf_4 fanout861 (.A(_05597_),
    .X(net861));
 sky130_fd_sc_hd__buf_4 fanout862 (.A(_05597_),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_2 fanout863 (.A(_05597_),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_4 fanout864 (.A(net868),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_2 fanout865 (.A(net868),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_4 fanout866 (.A(net868),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_2 fanout867 (.A(net868),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_16 fanout868 (.A(_05300_),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_4 fanout869 (.A(net870),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_4 fanout870 (.A(net872),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_4 fanout871 (.A(net872),
    .X(net871));
 sky130_fd_sc_hd__buf_4 fanout872 (.A(_05226_),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_4 fanout873 (.A(_05154_),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_4 fanout874 (.A(net876),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_2 fanout875 (.A(net876),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_4 fanout876 (.A(_05154_),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_4 fanout877 (.A(net880),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_4 fanout878 (.A(net879),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_4 fanout879 (.A(net880),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_2 fanout880 (.A(_05076_),
    .X(net880));
 sky130_fd_sc_hd__buf_4 fanout881 (.A(net882),
    .X(net881));
 sky130_fd_sc_hd__buf_4 fanout882 (.A(net883),
    .X(net882));
 sky130_fd_sc_hd__buf_4 fanout883 (.A(net884),
    .X(net883));
 sky130_fd_sc_hd__buf_4 fanout884 (.A(net885),
    .X(net884));
 sky130_fd_sc_hd__buf_4 fanout885 (.A(_05016_),
    .X(net885));
 sky130_fd_sc_hd__buf_6 fanout886 (.A(net887),
    .X(net886));
 sky130_fd_sc_hd__buf_4 fanout887 (.A(net888),
    .X(net887));
 sky130_fd_sc_hd__buf_4 fanout888 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__buf_8 fanout889 (.A(_04934_),
    .X(net889));
 sky130_fd_sc_hd__buf_4 fanout890 (.A(net892),
    .X(net890));
 sky130_fd_sc_hd__buf_2 fanout891 (.A(net892),
    .X(net891));
 sky130_fd_sc_hd__clkbuf_4 fanout892 (.A(_04853_),
    .X(net892));
 sky130_fd_sc_hd__buf_4 fanout893 (.A(net894),
    .X(net893));
 sky130_fd_sc_hd__buf_2 fanout894 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_4 fanout895 (.A(_04852_),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_4 fanout896 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_2 fanout897 (.A(_04322_),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_4 fanout898 (.A(net899),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_4 fanout899 (.A(_04322_),
    .X(net899));
 sky130_fd_sc_hd__clkbuf_4 fanout900 (.A(net903),
    .X(net900));
 sky130_fd_sc_hd__buf_2 fanout901 (.A(net903),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_4 fanout902 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__buf_6 fanout903 (.A(_04236_),
    .X(net903));
 sky130_fd_sc_hd__buf_12 fanout904 (.A(net907),
    .X(net904));
 sky130_fd_sc_hd__buf_12 fanout905 (.A(net906),
    .X(net905));
 sky130_fd_sc_hd__buf_12 fanout906 (.A(net907),
    .X(net906));
 sky130_fd_sc_hd__buf_8 fanout907 (.A(_03123_),
    .X(net907));
 sky130_fd_sc_hd__buf_12 fanout908 (.A(net911),
    .X(net908));
 sky130_fd_sc_hd__buf_12 fanout909 (.A(net910),
    .X(net909));
 sky130_fd_sc_hd__buf_12 fanout910 (.A(net911),
    .X(net910));
 sky130_fd_sc_hd__buf_12 fanout911 (.A(_03122_),
    .X(net911));
 sky130_fd_sc_hd__buf_8 fanout912 (.A(net913),
    .X(net912));
 sky130_fd_sc_hd__buf_12 fanout913 (.A(_03120_),
    .X(net913));
 sky130_fd_sc_hd__buf_12 fanout914 (.A(net915),
    .X(net914));
 sky130_fd_sc_hd__buf_8 fanout915 (.A(_03120_),
    .X(net915));
 sky130_fd_sc_hd__buf_12 fanout916 (.A(net919),
    .X(net916));
 sky130_fd_sc_hd__buf_12 fanout917 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__buf_12 fanout918 (.A(net919),
    .X(net918));
 sky130_fd_sc_hd__buf_8 fanout919 (.A(_03117_),
    .X(net919));
 sky130_fd_sc_hd__buf_12 fanout920 (.A(net923),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_16 fanout921 (.A(net922),
    .X(net921));
 sky130_fd_sc_hd__buf_12 fanout922 (.A(net923),
    .X(net922));
 sky130_fd_sc_hd__buf_8 fanout923 (.A(_03116_),
    .X(net923));
 sky130_fd_sc_hd__buf_12 fanout924 (.A(net927),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_16 fanout925 (.A(net926),
    .X(net925));
 sky130_fd_sc_hd__buf_12 fanout926 (.A(net927),
    .X(net926));
 sky130_fd_sc_hd__buf_12 fanout927 (.A(_03115_),
    .X(net927));
 sky130_fd_sc_hd__buf_4 fanout928 (.A(net929),
    .X(net928));
 sky130_fd_sc_hd__buf_2 fanout929 (.A(net930),
    .X(net929));
 sky130_fd_sc_hd__buf_2 fanout930 (.A(_02219_),
    .X(net930));
 sky130_fd_sc_hd__buf_6 fanout931 (.A(_02219_),
    .X(net931));
 sky130_fd_sc_hd__buf_2 fanout932 (.A(_02219_),
    .X(net932));
 sky130_fd_sc_hd__buf_4 fanout933 (.A(net935),
    .X(net933));
 sky130_fd_sc_hd__buf_4 fanout934 (.A(net935),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_4 fanout935 (.A(_01908_),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_4 fanout936 (.A(net938),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_2 fanout937 (.A(net938),
    .X(net937));
 sky130_fd_sc_hd__buf_4 fanout938 (.A(_01902_),
    .X(net938));
 sky130_fd_sc_hd__buf_4 fanout939 (.A(net941),
    .X(net939));
 sky130_fd_sc_hd__buf_4 fanout940 (.A(net941),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_4 fanout941 (.A(_01901_),
    .X(net941));
 sky130_fd_sc_hd__buf_4 fanout942 (.A(net944),
    .X(net942));
 sky130_fd_sc_hd__buf_4 fanout943 (.A(net944),
    .X(net943));
 sky130_fd_sc_hd__buf_4 fanout944 (.A(_01900_),
    .X(net944));
 sky130_fd_sc_hd__buf_4 fanout945 (.A(_01899_),
    .X(net945));
 sky130_fd_sc_hd__buf_2 fanout946 (.A(_01899_),
    .X(net946));
 sky130_fd_sc_hd__buf_4 fanout947 (.A(_01899_),
    .X(net947));
 sky130_fd_sc_hd__buf_2 fanout948 (.A(_01899_),
    .X(net948));
 sky130_fd_sc_hd__buf_12 fanout949 (.A(net952),
    .X(net949));
 sky130_fd_sc_hd__buf_12 fanout950 (.A(net951),
    .X(net950));
 sky130_fd_sc_hd__buf_12 fanout951 (.A(net952),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_16 fanout952 (.A(_01893_),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_16 fanout953 (.A(_08814_),
    .X(net953));
 sky130_fd_sc_hd__buf_4 fanout954 (.A(_08814_),
    .X(net954));
 sky130_fd_sc_hd__buf_12 fanout955 (.A(net956),
    .X(net955));
 sky130_fd_sc_hd__buf_12 fanout956 (.A(_08814_),
    .X(net956));
 sky130_fd_sc_hd__buf_12 fanout957 (.A(net960),
    .X(net957));
 sky130_fd_sc_hd__buf_12 fanout958 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__buf_12 fanout959 (.A(net960),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_16 fanout960 (.A(_08771_),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_16 fanout961 (.A(_08682_),
    .X(net961));
 sky130_fd_sc_hd__buf_8 fanout962 (.A(_08682_),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_16 fanout963 (.A(net964),
    .X(net963));
 sky130_fd_sc_hd__buf_8 fanout964 (.A(_08682_),
    .X(net964));
 sky130_fd_sc_hd__buf_12 fanout965 (.A(_08681_),
    .X(net965));
 sky130_fd_sc_hd__buf_6 fanout966 (.A(_08681_),
    .X(net966));
 sky130_fd_sc_hd__buf_12 fanout967 (.A(net968),
    .X(net967));
 sky130_fd_sc_hd__buf_12 fanout968 (.A(_08681_),
    .X(net968));
 sky130_fd_sc_hd__buf_12 fanout969 (.A(_08679_),
    .X(net969));
 sky130_fd_sc_hd__buf_6 fanout970 (.A(_08679_),
    .X(net970));
 sky130_fd_sc_hd__buf_12 fanout971 (.A(net972),
    .X(net971));
 sky130_fd_sc_hd__buf_12 fanout972 (.A(_08679_),
    .X(net972));
 sky130_fd_sc_hd__buf_6 fanout973 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__buf_6 fanout974 (.A(net977),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_16 fanout975 (.A(net977),
    .X(net975));
 sky130_fd_sc_hd__buf_4 fanout976 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__buf_4 fanout977 (.A(_07165_),
    .X(net977));
 sky130_fd_sc_hd__buf_6 fanout978 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__buf_4 fanout979 (.A(_07165_),
    .X(net979));
 sky130_fd_sc_hd__buf_6 fanout980 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_4 fanout981 (.A(_07165_),
    .X(net981));
 sky130_fd_sc_hd__buf_6 fanout982 (.A(net983),
    .X(net982));
 sky130_fd_sc_hd__buf_8 fanout983 (.A(net985),
    .X(net983));
 sky130_fd_sc_hd__buf_4 fanout984 (.A(net985),
    .X(net984));
 sky130_fd_sc_hd__buf_6 fanout985 (.A(_07152_),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_8 fanout986 (.A(net988),
    .X(net986));
 sky130_fd_sc_hd__buf_2 fanout987 (.A(net988),
    .X(net987));
 sky130_fd_sc_hd__buf_6 fanout988 (.A(_07151_),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_8 fanout990 (.A(_06635_),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_4 fanout991 (.A(_06635_),
    .X(net991));
 sky130_fd_sc_hd__buf_4 fanout992 (.A(_05519_),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_2 fanout993 (.A(_05519_),
    .X(net993));
 sky130_fd_sc_hd__clkbuf_4 fanout994 (.A(_05519_),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_4 fanout995 (.A(_05519_),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_4 fanout996 (.A(net997),
    .X(net996));
 sky130_fd_sc_hd__buf_2 fanout997 (.A(_05447_),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_4 fanout998 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__buf_4 fanout999 (.A(_05447_),
    .X(net999));
 sky130_fd_sc_hd__buf_8 input1 (.A(coreIndex[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(core_wb_data_i[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(dout0[61]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(dout0[62]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(dout0[63]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(dout0[6]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(dout0[7]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(dout0[8]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(dout0[9]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(dout1[0]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(dout1[10]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(dout1[11]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(core_wb_data_i[10]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(dout1[12]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(dout1[13]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 input112 (.A(dout1[14]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 input113 (.A(dout1[15]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(dout1[16]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(dout1[17]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(dout1[18]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(dout1[19]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(dout1[1]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(dout1[20]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(core_wb_data_i[11]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(dout1[21]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(dout1[22]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(dout1[23]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(dout1[24]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(dout1[25]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(dout1[26]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(dout1[27]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(dout1[28]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(dout1[29]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(dout1[2]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(core_wb_data_i[12]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(dout1[30]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(dout1[31]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(dout1[32]),
    .X(net132));
 sky130_fd_sc_hd__buf_2 input133 (.A(dout1[33]),
    .X(net133));
 sky130_fd_sc_hd__buf_2 input134 (.A(dout1[34]),
    .X(net134));
 sky130_fd_sc_hd__buf_2 input135 (.A(dout1[35]),
    .X(net135));
 sky130_fd_sc_hd__buf_2 input136 (.A(dout1[36]),
    .X(net136));
 sky130_fd_sc_hd__buf_2 input137 (.A(dout1[37]),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input138 (.A(dout1[38]),
    .X(net138));
 sky130_fd_sc_hd__buf_2 input139 (.A(dout1[39]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(core_wb_data_i[13]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input140 (.A(dout1[3]),
    .X(net140));
 sky130_fd_sc_hd__buf_2 input141 (.A(dout1[40]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(dout1[41]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(dout1[42]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 input144 (.A(dout1[43]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(dout1[44]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 input146 (.A(dout1[45]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(dout1[46]),
    .X(net147));
 sky130_fd_sc_hd__buf_2 input148 (.A(dout1[47]),
    .X(net148));
 sky130_fd_sc_hd__buf_2 input149 (.A(dout1[48]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(core_wb_data_i[14]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input150 (.A(dout1[49]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 input151 (.A(dout1[4]),
    .X(net151));
 sky130_fd_sc_hd__buf_2 input152 (.A(dout1[50]),
    .X(net152));
 sky130_fd_sc_hd__buf_2 input153 (.A(dout1[51]),
    .X(net153));
 sky130_fd_sc_hd__buf_2 input154 (.A(dout1[52]),
    .X(net154));
 sky130_fd_sc_hd__buf_2 input155 (.A(dout1[53]),
    .X(net155));
 sky130_fd_sc_hd__buf_2 input156 (.A(dout1[54]),
    .X(net156));
 sky130_fd_sc_hd__buf_2 input157 (.A(dout1[55]),
    .X(net157));
 sky130_fd_sc_hd__buf_2 input158 (.A(dout1[56]),
    .X(net158));
 sky130_fd_sc_hd__buf_2 input159 (.A(dout1[57]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(core_wb_data_i[15]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input160 (.A(dout1[58]),
    .X(net160));
 sky130_fd_sc_hd__buf_2 input161 (.A(dout1[59]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 input162 (.A(dout1[5]),
    .X(net162));
 sky130_fd_sc_hd__buf_2 input163 (.A(dout1[60]),
    .X(net163));
 sky130_fd_sc_hd__buf_2 input164 (.A(dout1[61]),
    .X(net164));
 sky130_fd_sc_hd__buf_2 input165 (.A(dout1[62]),
    .X(net165));
 sky130_fd_sc_hd__buf_2 input166 (.A(dout1[63]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 input167 (.A(dout1[6]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 input168 (.A(dout1[7]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 input169 (.A(dout1[8]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(core_wb_data_i[16]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input170 (.A(dout1[9]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 input171 (.A(irq[0]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(irq[10]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 input173 (.A(irq[11]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 input174 (.A(irq[12]),
    .X(net174));
 sky130_fd_sc_hd__buf_2 input175 (.A(irq[13]),
    .X(net175));
 sky130_fd_sc_hd__buf_4 input176 (.A(irq[14]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 input177 (.A(irq[15]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 input178 (.A(irq[1]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 input179 (.A(irq[2]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(core_wb_data_i[17]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(irq[3]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 input181 (.A(irq[4]),
    .X(net181));
 sky130_fd_sc_hd__buf_2 input182 (.A(irq[5]),
    .X(net182));
 sky130_fd_sc_hd__buf_2 input183 (.A(irq[6]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 input184 (.A(irq[7]),
    .X(net184));
 sky130_fd_sc_hd__buf_2 input185 (.A(irq[8]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(irq[9]),
    .X(net186));
 sky130_fd_sc_hd__buf_4 input187 (.A(jtag_tck),
    .X(net187));
 sky130_fd_sc_hd__buf_12 input188 (.A(jtag_tdi),
    .X(net188));
 sky130_fd_sc_hd__buf_6 input189 (.A(jtag_tms),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(core_wb_data_i[18]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(localMemory_wb_adr_i[0]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 input191 (.A(localMemory_wb_adr_i[10]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 input192 (.A(localMemory_wb_adr_i[11]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_2 input193 (.A(localMemory_wb_adr_i[12]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 input194 (.A(localMemory_wb_adr_i[13]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input195 (.A(localMemory_wb_adr_i[14]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 input196 (.A(localMemory_wb_adr_i[15]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 input197 (.A(localMemory_wb_adr_i[16]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(localMemory_wb_adr_i[17]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 input199 (.A(localMemory_wb_adr_i[18]),
    .X(net199));
 sky130_fd_sc_hd__buf_8 input2 (.A(coreIndex[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(core_wb_data_i[19]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input200 (.A(localMemory_wb_adr_i[19]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 input201 (.A(localMemory_wb_adr_i[1]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 input202 (.A(localMemory_wb_adr_i[20]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 input203 (.A(localMemory_wb_adr_i[21]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 input204 (.A(localMemory_wb_adr_i[22]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_8 input205 (.A(localMemory_wb_adr_i[23]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 input206 (.A(localMemory_wb_adr_i[2]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 input207 (.A(localMemory_wb_adr_i[3]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 input208 (.A(localMemory_wb_adr_i[4]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 input209 (.A(localMemory_wb_adr_i[5]),
    .X(net209));
 sky130_fd_sc_hd__buf_2 input21 (.A(core_wb_data_i[1]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input210 (.A(localMemory_wb_adr_i[6]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 input211 (.A(localMemory_wb_adr_i[7]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 input212 (.A(localMemory_wb_adr_i[8]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(localMemory_wb_adr_i[9]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 input214 (.A(localMemory_wb_cyc_i),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_16 input215 (.A(localMemory_wb_data_i[0]),
    .X(net215));
 sky130_fd_sc_hd__buf_8 input216 (.A(localMemory_wb_data_i[10]),
    .X(net216));
 sky130_fd_sc_hd__buf_8 input217 (.A(localMemory_wb_data_i[11]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_16 input218 (.A(localMemory_wb_data_i[12]),
    .X(net218));
 sky130_fd_sc_hd__buf_8 input219 (.A(localMemory_wb_data_i[13]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(core_wb_data_i[20]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_16 input220 (.A(localMemory_wb_data_i[14]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_16 input221 (.A(localMemory_wb_data_i[15]),
    .X(net221));
 sky130_fd_sc_hd__buf_8 input222 (.A(localMemory_wb_data_i[16]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_16 input223 (.A(localMemory_wb_data_i[17]),
    .X(net223));
 sky130_fd_sc_hd__buf_8 input224 (.A(localMemory_wb_data_i[18]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_16 input225 (.A(localMemory_wb_data_i[19]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_16 input226 (.A(localMemory_wb_data_i[1]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_16 input227 (.A(localMemory_wb_data_i[20]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_16 input228 (.A(localMemory_wb_data_i[21]),
    .X(net228));
 sky130_fd_sc_hd__buf_12 input229 (.A(localMemory_wb_data_i[22]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(core_wb_data_i[21]),
    .X(net23));
 sky130_fd_sc_hd__buf_12 input230 (.A(localMemory_wb_data_i[23]),
    .X(net230));
 sky130_fd_sc_hd__buf_12 input231 (.A(localMemory_wb_data_i[24]),
    .X(net231));
 sky130_fd_sc_hd__buf_12 input232 (.A(localMemory_wb_data_i[25]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_16 input233 (.A(localMemory_wb_data_i[26]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_16 input234 (.A(localMemory_wb_data_i[27]),
    .X(net234));
 sky130_fd_sc_hd__buf_12 input235 (.A(localMemory_wb_data_i[28]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_16 input236 (.A(localMemory_wb_data_i[29]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_16 input237 (.A(localMemory_wb_data_i[2]),
    .X(net237));
 sky130_fd_sc_hd__buf_12 input238 (.A(localMemory_wb_data_i[30]),
    .X(net238));
 sky130_fd_sc_hd__buf_12 input239 (.A(localMemory_wb_data_i[31]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(core_wb_data_i[22]),
    .X(net24));
 sky130_fd_sc_hd__buf_8 input240 (.A(localMemory_wb_data_i[3]),
    .X(net240));
 sky130_fd_sc_hd__buf_8 input241 (.A(localMemory_wb_data_i[4]),
    .X(net241));
 sky130_fd_sc_hd__buf_8 input242 (.A(localMemory_wb_data_i[5]),
    .X(net242));
 sky130_fd_sc_hd__buf_8 input243 (.A(localMemory_wb_data_i[6]),
    .X(net243));
 sky130_fd_sc_hd__buf_8 input244 (.A(localMemory_wb_data_i[7]),
    .X(net244));
 sky130_fd_sc_hd__buf_8 input245 (.A(localMemory_wb_data_i[8]),
    .X(net245));
 sky130_fd_sc_hd__buf_8 input246 (.A(localMemory_wb_data_i[9]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 input247 (.A(localMemory_wb_sel_i[0]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 input248 (.A(localMemory_wb_sel_i[1]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 input249 (.A(localMemory_wb_sel_i[2]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(core_wb_data_i[23]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input250 (.A(localMemory_wb_sel_i[3]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 input251 (.A(localMemory_wb_stb_i),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_2 input252 (.A(localMemory_wb_we_i),
    .X(net252));
 sky130_fd_sc_hd__buf_4 input253 (.A(manufacturerID[0]),
    .X(net253));
 sky130_fd_sc_hd__buf_4 input254 (.A(manufacturerID[10]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_4 input255 (.A(manufacturerID[1]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 input256 (.A(manufacturerID[2]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 input257 (.A(manufacturerID[3]),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_4 input258 (.A(manufacturerID[4]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 input259 (.A(manufacturerID[5]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(core_wb_data_i[24]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input260 (.A(manufacturerID[6]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 input261 (.A(manufacturerID[7]),
    .X(net261));
 sky130_fd_sc_hd__buf_4 input262 (.A(manufacturerID[8]),
    .X(net262));
 sky130_fd_sc_hd__buf_4 input263 (.A(manufacturerID[9]),
    .X(net263));
 sky130_fd_sc_hd__buf_2 input264 (.A(partID[0]),
    .X(net264));
 sky130_fd_sc_hd__buf_2 input265 (.A(partID[10]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_2 input266 (.A(partID[11]),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 input267 (.A(partID[12]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 input268 (.A(partID[13]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 input269 (.A(partID[14]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(core_wb_data_i[25]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input270 (.A(partID[15]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 input271 (.A(partID[1]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 input272 (.A(partID[2]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 input273 (.A(partID[3]),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_2 input274 (.A(partID[4]),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_2 input275 (.A(partID[5]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 input276 (.A(partID[6]),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 input277 (.A(partID[7]),
    .X(net277));
 sky130_fd_sc_hd__buf_2 input278 (.A(partID[8]),
    .X(net278));
 sky130_fd_sc_hd__buf_2 input279 (.A(partID[9]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(core_wb_data_i[26]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input280 (.A(versionID[0]),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_2 input281 (.A(versionID[1]),
    .X(net281));
 sky130_fd_sc_hd__buf_2 input282 (.A(versionID[2]),
    .X(net282));
 sky130_fd_sc_hd__buf_2 input283 (.A(versionID[3]),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_2 input284 (.A(wb_rst_i),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(core_wb_data_i[27]),
    .X(net29));
 sky130_fd_sc_hd__buf_8 input3 (.A(coreIndex[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(core_wb_data_i[28]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(core_wb_data_i[29]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(core_wb_data_i[2]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(core_wb_data_i[30]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(core_wb_data_i[31]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(core_wb_data_i[3]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(core_wb_data_i[4]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(core_wb_data_i[5]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(core_wb_data_i[6]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(core_wb_data_i[7]),
    .X(net39));
 sky130_fd_sc_hd__buf_6 input4 (.A(coreIndex[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input40 (.A(core_wb_data_i[8]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(core_wb_data_i[9]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(core_wb_error_i),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(dout0[0]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(dout0[10]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(dout0[11]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(dout0[12]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(dout0[13]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(dout0[14]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(dout0[15]),
    .X(net49));
 sky130_fd_sc_hd__buf_6 input5 (.A(coreIndex[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(dout0[16]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(dout0[17]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(dout0[18]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(dout0[19]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(dout0[1]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(dout0[20]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(dout0[21]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(dout0[22]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(dout0[23]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(dout0[24]),
    .X(net59));
 sky130_fd_sc_hd__buf_6 input6 (.A(coreIndex[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(dout0[25]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(dout0[26]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(dout0[27]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(dout0[28]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(dout0[29]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(dout0[2]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(dout0[30]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(dout0[31]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(dout0[32]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(dout0[33]),
    .X(net69));
 sky130_fd_sc_hd__buf_6 input7 (.A(coreIndex[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(dout0[34]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(dout0[35]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(dout0[36]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(dout0[37]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(dout0[38]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(dout0[39]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input76 (.A(dout0[3]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(dout0[40]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(dout0[41]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(dout0[42]),
    .X(net79));
 sky130_fd_sc_hd__buf_6 input8 (.A(coreIndex[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(dout0[43]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(dout0[44]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(dout0[45]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(dout0[46]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(dout0[47]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(dout0[48]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(dout0[49]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(dout0[4]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(dout0[50]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(dout0[51]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(core_wb_ack_i),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(dout0[52]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 input91 (.A(dout0[53]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(dout0[54]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(dout0[55]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(dout0[56]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(dout0[57]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(dout0[58]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(dout0[59]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(dout0[5]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(dout0[60]),
    .X(net99));
 sky130_fd_sc_hd__buf_4 output285 (.A(net285),
    .X(addr0[0]));
 sky130_fd_sc_hd__buf_4 output286 (.A(net286),
    .X(addr0[1]));
 sky130_fd_sc_hd__buf_4 output287 (.A(net287),
    .X(addr0[2]));
 sky130_fd_sc_hd__buf_4 output288 (.A(net288),
    .X(addr0[3]));
 sky130_fd_sc_hd__buf_4 output289 (.A(net289),
    .X(addr0[4]));
 sky130_fd_sc_hd__buf_4 output290 (.A(net290),
    .X(addr0[5]));
 sky130_fd_sc_hd__buf_4 output291 (.A(net291),
    .X(addr0[6]));
 sky130_fd_sc_hd__buf_4 output292 (.A(net292),
    .X(addr0[7]));
 sky130_fd_sc_hd__buf_4 output293 (.A(net293),
    .X(addr0[8]));
 sky130_fd_sc_hd__buf_4 output294 (.A(net294),
    .X(addr1[0]));
 sky130_fd_sc_hd__buf_4 output295 (.A(net295),
    .X(addr1[1]));
 sky130_fd_sc_hd__buf_4 output296 (.A(net296),
    .X(addr1[2]));
 sky130_fd_sc_hd__buf_4 output297 (.A(net297),
    .X(addr1[3]));
 sky130_fd_sc_hd__buf_4 output298 (.A(net298),
    .X(addr1[4]));
 sky130_fd_sc_hd__buf_4 output299 (.A(net299),
    .X(addr1[5]));
 sky130_fd_sc_hd__buf_4 output300 (.A(net300),
    .X(addr1[6]));
 sky130_fd_sc_hd__buf_4 output301 (.A(net301),
    .X(addr1[7]));
 sky130_fd_sc_hd__buf_4 output302 (.A(net302),
    .X(addr1[8]));
 sky130_fd_sc_hd__clkbuf_2 output303 (.A(net303),
    .X(clk0));
 sky130_fd_sc_hd__clkbuf_2 output304 (.A(net304),
    .X(clk1));
 sky130_fd_sc_hd__buf_4 output305 (.A(net305),
    .X(core_wb_adr_o[0]));
 sky130_fd_sc_hd__buf_4 output306 (.A(net306),
    .X(core_wb_adr_o[10]));
 sky130_fd_sc_hd__buf_4 output307 (.A(net307),
    .X(core_wb_adr_o[11]));
 sky130_fd_sc_hd__buf_4 output308 (.A(net308),
    .X(core_wb_adr_o[12]));
 sky130_fd_sc_hd__buf_4 output309 (.A(net309),
    .X(core_wb_adr_o[13]));
 sky130_fd_sc_hd__buf_4 output310 (.A(net310),
    .X(core_wb_adr_o[14]));
 sky130_fd_sc_hd__buf_4 output311 (.A(net311),
    .X(core_wb_adr_o[15]));
 sky130_fd_sc_hd__buf_4 output312 (.A(net312),
    .X(core_wb_adr_o[16]));
 sky130_fd_sc_hd__buf_4 output313 (.A(net313),
    .X(core_wb_adr_o[17]));
 sky130_fd_sc_hd__buf_4 output314 (.A(net314),
    .X(core_wb_adr_o[18]));
 sky130_fd_sc_hd__buf_4 output315 (.A(net315),
    .X(core_wb_adr_o[19]));
 sky130_fd_sc_hd__buf_4 output316 (.A(net316),
    .X(core_wb_adr_o[1]));
 sky130_fd_sc_hd__buf_4 output317 (.A(net317),
    .X(core_wb_adr_o[20]));
 sky130_fd_sc_hd__buf_4 output318 (.A(net318),
    .X(core_wb_adr_o[21]));
 sky130_fd_sc_hd__buf_4 output319 (.A(net319),
    .X(core_wb_adr_o[22]));
 sky130_fd_sc_hd__buf_4 output320 (.A(net320),
    .X(core_wb_adr_o[23]));
 sky130_fd_sc_hd__buf_4 output321 (.A(net321),
    .X(core_wb_adr_o[24]));
 sky130_fd_sc_hd__buf_4 output322 (.A(net322),
    .X(core_wb_adr_o[25]));
 sky130_fd_sc_hd__buf_4 output323 (.A(net323),
    .X(core_wb_adr_o[26]));
 sky130_fd_sc_hd__buf_4 output324 (.A(net324),
    .X(core_wb_adr_o[27]));
 sky130_fd_sc_hd__buf_4 output325 (.A(net325),
    .X(core_wb_adr_o[2]));
 sky130_fd_sc_hd__buf_4 output326 (.A(net326),
    .X(core_wb_adr_o[3]));
 sky130_fd_sc_hd__buf_4 output327 (.A(net327),
    .X(core_wb_adr_o[4]));
 sky130_fd_sc_hd__buf_4 output328 (.A(net328),
    .X(core_wb_adr_o[5]));
 sky130_fd_sc_hd__buf_4 output329 (.A(net329),
    .X(core_wb_adr_o[6]));
 sky130_fd_sc_hd__buf_4 output330 (.A(net330),
    .X(core_wb_adr_o[7]));
 sky130_fd_sc_hd__buf_4 output331 (.A(net331),
    .X(core_wb_adr_o[8]));
 sky130_fd_sc_hd__buf_4 output332 (.A(net332),
    .X(core_wb_adr_o[9]));
 sky130_fd_sc_hd__buf_4 output333 (.A(net333),
    .X(core_wb_cyc_o));
 sky130_fd_sc_hd__buf_4 output334 (.A(net334),
    .X(core_wb_data_o[0]));
 sky130_fd_sc_hd__buf_4 output335 (.A(net335),
    .X(core_wb_data_o[10]));
 sky130_fd_sc_hd__buf_4 output336 (.A(net336),
    .X(core_wb_data_o[11]));
 sky130_fd_sc_hd__buf_4 output337 (.A(net337),
    .X(core_wb_data_o[12]));
 sky130_fd_sc_hd__buf_4 output338 (.A(net338),
    .X(core_wb_data_o[13]));
 sky130_fd_sc_hd__buf_4 output339 (.A(net339),
    .X(core_wb_data_o[14]));
 sky130_fd_sc_hd__buf_4 output340 (.A(net340),
    .X(core_wb_data_o[15]));
 sky130_fd_sc_hd__buf_4 output341 (.A(net341),
    .X(core_wb_data_o[16]));
 sky130_fd_sc_hd__buf_4 output342 (.A(net342),
    .X(core_wb_data_o[17]));
 sky130_fd_sc_hd__buf_4 output343 (.A(net343),
    .X(core_wb_data_o[18]));
 sky130_fd_sc_hd__buf_4 output344 (.A(net344),
    .X(core_wb_data_o[19]));
 sky130_fd_sc_hd__buf_4 output345 (.A(net345),
    .X(core_wb_data_o[1]));
 sky130_fd_sc_hd__buf_4 output346 (.A(net346),
    .X(core_wb_data_o[20]));
 sky130_fd_sc_hd__buf_4 output347 (.A(net347),
    .X(core_wb_data_o[21]));
 sky130_fd_sc_hd__buf_4 output348 (.A(net348),
    .X(core_wb_data_o[22]));
 sky130_fd_sc_hd__buf_4 output349 (.A(net349),
    .X(core_wb_data_o[23]));
 sky130_fd_sc_hd__buf_4 output350 (.A(net350),
    .X(core_wb_data_o[24]));
 sky130_fd_sc_hd__buf_4 output351 (.A(net351),
    .X(core_wb_data_o[25]));
 sky130_fd_sc_hd__buf_4 output352 (.A(net352),
    .X(core_wb_data_o[26]));
 sky130_fd_sc_hd__buf_4 output353 (.A(net353),
    .X(core_wb_data_o[27]));
 sky130_fd_sc_hd__buf_4 output354 (.A(net354),
    .X(core_wb_data_o[28]));
 sky130_fd_sc_hd__buf_4 output355 (.A(net355),
    .X(core_wb_data_o[29]));
 sky130_fd_sc_hd__buf_4 output356 (.A(net356),
    .X(core_wb_data_o[2]));
 sky130_fd_sc_hd__buf_4 output357 (.A(net357),
    .X(core_wb_data_o[30]));
 sky130_fd_sc_hd__buf_4 output358 (.A(net358),
    .X(core_wb_data_o[31]));
 sky130_fd_sc_hd__buf_4 output359 (.A(net359),
    .X(core_wb_data_o[3]));
 sky130_fd_sc_hd__buf_4 output360 (.A(net360),
    .X(core_wb_data_o[4]));
 sky130_fd_sc_hd__buf_4 output361 (.A(net361),
    .X(core_wb_data_o[5]));
 sky130_fd_sc_hd__buf_4 output362 (.A(net362),
    .X(core_wb_data_o[6]));
 sky130_fd_sc_hd__buf_4 output363 (.A(net363),
    .X(core_wb_data_o[7]));
 sky130_fd_sc_hd__buf_4 output364 (.A(net364),
    .X(core_wb_data_o[8]));
 sky130_fd_sc_hd__buf_4 output365 (.A(net365),
    .X(core_wb_data_o[9]));
 sky130_fd_sc_hd__buf_4 output366 (.A(net366),
    .X(core_wb_sel_o[0]));
 sky130_fd_sc_hd__buf_4 output367 (.A(net367),
    .X(core_wb_sel_o[1]));
 sky130_fd_sc_hd__buf_4 output368 (.A(net368),
    .X(core_wb_sel_o[2]));
 sky130_fd_sc_hd__buf_4 output369 (.A(net369),
    .X(core_wb_sel_o[3]));
 sky130_fd_sc_hd__buf_4 output370 (.A(net370),
    .X(core_wb_stb_o));
 sky130_fd_sc_hd__buf_4 output371 (.A(net371),
    .X(core_wb_we_o));
 sky130_fd_sc_hd__buf_4 output372 (.A(net372),
    .X(csb0[0]));
 sky130_fd_sc_hd__buf_4 output373 (.A(net373),
    .X(csb0[1]));
 sky130_fd_sc_hd__buf_4 output374 (.A(net374),
    .X(csb1[0]));
 sky130_fd_sc_hd__buf_4 output375 (.A(net375),
    .X(csb1[1]));
 sky130_fd_sc_hd__buf_4 output376 (.A(net376),
    .X(din0[0]));
 sky130_fd_sc_hd__buf_4 output377 (.A(net377),
    .X(din0[10]));
 sky130_fd_sc_hd__buf_4 output378 (.A(net378),
    .X(din0[11]));
 sky130_fd_sc_hd__buf_4 output379 (.A(net379),
    .X(din0[12]));
 sky130_fd_sc_hd__buf_4 output380 (.A(net380),
    .X(din0[13]));
 sky130_fd_sc_hd__buf_4 output381 (.A(net381),
    .X(din0[14]));
 sky130_fd_sc_hd__buf_4 output382 (.A(net382),
    .X(din0[15]));
 sky130_fd_sc_hd__buf_4 output383 (.A(net383),
    .X(din0[16]));
 sky130_fd_sc_hd__buf_4 output384 (.A(net384),
    .X(din0[17]));
 sky130_fd_sc_hd__buf_4 output385 (.A(net385),
    .X(din0[18]));
 sky130_fd_sc_hd__buf_4 output386 (.A(net386),
    .X(din0[19]));
 sky130_fd_sc_hd__buf_4 output387 (.A(net387),
    .X(din0[1]));
 sky130_fd_sc_hd__buf_4 output388 (.A(net388),
    .X(din0[20]));
 sky130_fd_sc_hd__buf_4 output389 (.A(net389),
    .X(din0[21]));
 sky130_fd_sc_hd__buf_4 output390 (.A(net390),
    .X(din0[22]));
 sky130_fd_sc_hd__buf_4 output391 (.A(net391),
    .X(din0[23]));
 sky130_fd_sc_hd__buf_4 output392 (.A(net392),
    .X(din0[24]));
 sky130_fd_sc_hd__buf_4 output393 (.A(net393),
    .X(din0[25]));
 sky130_fd_sc_hd__buf_4 output394 (.A(net394),
    .X(din0[26]));
 sky130_fd_sc_hd__buf_4 output395 (.A(net395),
    .X(din0[27]));
 sky130_fd_sc_hd__buf_4 output396 (.A(net396),
    .X(din0[28]));
 sky130_fd_sc_hd__buf_4 output397 (.A(net397),
    .X(din0[29]));
 sky130_fd_sc_hd__buf_4 output398 (.A(net398),
    .X(din0[2]));
 sky130_fd_sc_hd__buf_4 output399 (.A(net399),
    .X(din0[30]));
 sky130_fd_sc_hd__buf_4 output400 (.A(net400),
    .X(din0[31]));
 sky130_fd_sc_hd__buf_4 output401 (.A(net401),
    .X(din0[3]));
 sky130_fd_sc_hd__buf_4 output402 (.A(net402),
    .X(din0[4]));
 sky130_fd_sc_hd__buf_4 output403 (.A(net403),
    .X(din0[5]));
 sky130_fd_sc_hd__buf_4 output404 (.A(net404),
    .X(din0[6]));
 sky130_fd_sc_hd__buf_4 output405 (.A(net405),
    .X(din0[7]));
 sky130_fd_sc_hd__buf_4 output406 (.A(net406),
    .X(din0[8]));
 sky130_fd_sc_hd__buf_4 output407 (.A(net407),
    .X(din0[9]));
 sky130_fd_sc_hd__buf_4 output408 (.A(net408),
    .X(jtag_tdo));
 sky130_fd_sc_hd__buf_4 output409 (.A(net409),
    .X(localMemory_wb_ack_o));
 sky130_fd_sc_hd__buf_4 output410 (.A(net410),
    .X(localMemory_wb_data_o[0]));
 sky130_fd_sc_hd__buf_4 output411 (.A(net411),
    .X(localMemory_wb_data_o[10]));
 sky130_fd_sc_hd__buf_4 output412 (.A(net412),
    .X(localMemory_wb_data_o[11]));
 sky130_fd_sc_hd__buf_4 output413 (.A(net413),
    .X(localMemory_wb_data_o[12]));
 sky130_fd_sc_hd__buf_4 output414 (.A(net414),
    .X(localMemory_wb_data_o[13]));
 sky130_fd_sc_hd__buf_4 output415 (.A(net415),
    .X(localMemory_wb_data_o[14]));
 sky130_fd_sc_hd__buf_4 output416 (.A(net416),
    .X(localMemory_wb_data_o[15]));
 sky130_fd_sc_hd__buf_4 output417 (.A(net417),
    .X(localMemory_wb_data_o[16]));
 sky130_fd_sc_hd__buf_4 output418 (.A(net418),
    .X(localMemory_wb_data_o[17]));
 sky130_fd_sc_hd__buf_4 output419 (.A(net419),
    .X(localMemory_wb_data_o[18]));
 sky130_fd_sc_hd__buf_4 output420 (.A(net420),
    .X(localMemory_wb_data_o[19]));
 sky130_fd_sc_hd__buf_4 output421 (.A(net421),
    .X(localMemory_wb_data_o[1]));
 sky130_fd_sc_hd__buf_4 output422 (.A(net422),
    .X(localMemory_wb_data_o[20]));
 sky130_fd_sc_hd__buf_4 output423 (.A(net423),
    .X(localMemory_wb_data_o[21]));
 sky130_fd_sc_hd__buf_4 output424 (.A(net424),
    .X(localMemory_wb_data_o[22]));
 sky130_fd_sc_hd__buf_4 output425 (.A(net425),
    .X(localMemory_wb_data_o[23]));
 sky130_fd_sc_hd__buf_4 output426 (.A(net426),
    .X(localMemory_wb_data_o[24]));
 sky130_fd_sc_hd__buf_4 output427 (.A(net427),
    .X(localMemory_wb_data_o[25]));
 sky130_fd_sc_hd__buf_4 output428 (.A(net428),
    .X(localMemory_wb_data_o[26]));
 sky130_fd_sc_hd__buf_4 output429 (.A(net429),
    .X(localMemory_wb_data_o[27]));
 sky130_fd_sc_hd__buf_4 output430 (.A(net430),
    .X(localMemory_wb_data_o[28]));
 sky130_fd_sc_hd__buf_4 output431 (.A(net431),
    .X(localMemory_wb_data_o[29]));
 sky130_fd_sc_hd__buf_4 output432 (.A(net432),
    .X(localMemory_wb_data_o[2]));
 sky130_fd_sc_hd__buf_4 output433 (.A(net433),
    .X(localMemory_wb_data_o[30]));
 sky130_fd_sc_hd__buf_4 output434 (.A(net434),
    .X(localMemory_wb_data_o[31]));
 sky130_fd_sc_hd__buf_4 output435 (.A(net435),
    .X(localMemory_wb_data_o[3]));
 sky130_fd_sc_hd__buf_4 output436 (.A(net436),
    .X(localMemory_wb_data_o[4]));
 sky130_fd_sc_hd__buf_4 output437 (.A(net437),
    .X(localMemory_wb_data_o[5]));
 sky130_fd_sc_hd__buf_4 output438 (.A(net438),
    .X(localMemory_wb_data_o[6]));
 sky130_fd_sc_hd__buf_4 output439 (.A(net439),
    .X(localMemory_wb_data_o[7]));
 sky130_fd_sc_hd__buf_4 output440 (.A(net440),
    .X(localMemory_wb_data_o[8]));
 sky130_fd_sc_hd__buf_4 output441 (.A(net441),
    .X(localMemory_wb_data_o[9]));
 sky130_fd_sc_hd__buf_4 output442 (.A(net442),
    .X(localMemory_wb_stall_o));
 sky130_fd_sc_hd__buf_4 output443 (.A(net443),
    .X(probe_env[0]));
 sky130_fd_sc_hd__buf_4 output444 (.A(net444),
    .X(probe_env[1]));
 sky130_fd_sc_hd__buf_4 output445 (.A(net445),
    .X(probe_jtagInstruction[0]));
 sky130_fd_sc_hd__buf_4 output446 (.A(net446),
    .X(probe_jtagInstruction[1]));
 sky130_fd_sc_hd__buf_4 output447 (.A(net447),
    .X(probe_jtagInstruction[2]));
 sky130_fd_sc_hd__buf_4 output448 (.A(net448),
    .X(probe_jtagInstruction[3]));
 sky130_fd_sc_hd__buf_4 output449 (.A(net449),
    .X(probe_jtagInstruction[4]));
 sky130_fd_sc_hd__buf_4 output450 (.A(net450),
    .X(probe_programCounter[0]));
 sky130_fd_sc_hd__buf_4 output451 (.A(net451),
    .X(probe_programCounter[10]));
 sky130_fd_sc_hd__buf_4 output452 (.A(net452),
    .X(probe_programCounter[11]));
 sky130_fd_sc_hd__buf_4 output453 (.A(net453),
    .X(probe_programCounter[12]));
 sky130_fd_sc_hd__buf_4 output454 (.A(net454),
    .X(probe_programCounter[13]));
 sky130_fd_sc_hd__buf_4 output455 (.A(net455),
    .X(probe_programCounter[14]));
 sky130_fd_sc_hd__buf_4 output456 (.A(net456),
    .X(probe_programCounter[15]));
 sky130_fd_sc_hd__buf_4 output457 (.A(net1747),
    .X(probe_programCounter[16]));
 sky130_fd_sc_hd__buf_4 output458 (.A(net458),
    .X(probe_programCounter[17]));
 sky130_fd_sc_hd__buf_4 output459 (.A(net459),
    .X(probe_programCounter[18]));
 sky130_fd_sc_hd__buf_4 output460 (.A(net460),
    .X(probe_programCounter[19]));
 sky130_fd_sc_hd__buf_4 output461 (.A(net461),
    .X(probe_programCounter[1]));
 sky130_fd_sc_hd__buf_4 output462 (.A(net462),
    .X(probe_programCounter[20]));
 sky130_fd_sc_hd__buf_4 output463 (.A(net463),
    .X(probe_programCounter[21]));
 sky130_fd_sc_hd__buf_4 output464 (.A(net464),
    .X(probe_programCounter[22]));
 sky130_fd_sc_hd__buf_4 output465 (.A(net465),
    .X(probe_programCounter[23]));
 sky130_fd_sc_hd__buf_4 output466 (.A(net466),
    .X(probe_programCounter[24]));
 sky130_fd_sc_hd__buf_4 output467 (.A(net467),
    .X(probe_programCounter[25]));
 sky130_fd_sc_hd__buf_4 output468 (.A(net468),
    .X(probe_programCounter[26]));
 sky130_fd_sc_hd__buf_4 output469 (.A(net469),
    .X(probe_programCounter[27]));
 sky130_fd_sc_hd__buf_4 output470 (.A(net470),
    .X(probe_programCounter[28]));
 sky130_fd_sc_hd__buf_4 output471 (.A(net471),
    .X(probe_programCounter[29]));
 sky130_fd_sc_hd__buf_4 output472 (.A(net472),
    .X(probe_programCounter[2]));
 sky130_fd_sc_hd__buf_4 output473 (.A(net473),
    .X(probe_programCounter[30]));
 sky130_fd_sc_hd__buf_4 output474 (.A(net474),
    .X(probe_programCounter[31]));
 sky130_fd_sc_hd__buf_4 output475 (.A(net475),
    .X(probe_programCounter[3]));
 sky130_fd_sc_hd__buf_4 output476 (.A(net1748),
    .X(probe_programCounter[4]));
 sky130_fd_sc_hd__buf_4 output477 (.A(net477),
    .X(probe_programCounter[5]));
 sky130_fd_sc_hd__buf_4 output478 (.A(net478),
    .X(probe_programCounter[6]));
 sky130_fd_sc_hd__buf_4 output479 (.A(net479),
    .X(probe_programCounter[7]));
 sky130_fd_sc_hd__buf_4 output480 (.A(net480),
    .X(probe_programCounter[8]));
 sky130_fd_sc_hd__buf_4 output481 (.A(net481),
    .X(probe_programCounter[9]));
 sky130_fd_sc_hd__buf_4 output482 (.A(net1719),
    .X(probe_state));
 sky130_fd_sc_hd__buf_4 output483 (.A(net483),
    .X(web0));
 sky130_fd_sc_hd__buf_4 output484 (.A(net484),
    .X(wmask0[0]));
 sky130_fd_sc_hd__buf_4 output485 (.A(net485),
    .X(wmask0[1]));
 sky130_fd_sc_hd__buf_4 output486 (.A(net486),
    .X(wmask0[2]));
 sky130_fd_sc_hd__buf_4 output487 (.A(net487),
    .X(wmask0[3]));
 sky130_fd_sc_hd__buf_6 wire1236 (.A(_06701_),
    .X(net1236));
 sky130_fd_sc_hd__buf_6 wire989 (.A(_06738_),
    .X(net989));
 assign localMemory_wb_error_o = net1911;
endmodule

