magic
tech sky130A
magscale 1 2
timestamp 1653408436
<< obsli1 >>
rect 1104 2159 118864 157777
<< obsm1 >>
rect 1026 1368 119126 157956
<< metal2 >>
rect 754 159200 810 160000
rect 2318 159200 2374 160000
rect 3882 159200 3938 160000
rect 5446 159200 5502 160000
rect 7010 159200 7066 160000
rect 8574 159200 8630 160000
rect 10138 159200 10194 160000
rect 11794 159200 11850 160000
rect 13358 159200 13414 160000
rect 14922 159200 14978 160000
rect 16486 159200 16542 160000
rect 18050 159200 18106 160000
rect 19614 159200 19670 160000
rect 21270 159200 21326 160000
rect 22834 159200 22890 160000
rect 24398 159200 24454 160000
rect 25962 159200 26018 160000
rect 27526 159200 27582 160000
rect 29090 159200 29146 160000
rect 30746 159200 30802 160000
rect 32310 159200 32366 160000
rect 33874 159200 33930 160000
rect 35438 159200 35494 160000
rect 37002 159200 37058 160000
rect 38566 159200 38622 160000
rect 40130 159200 40186 160000
rect 41786 159200 41842 160000
rect 43350 159200 43406 160000
rect 44914 159200 44970 160000
rect 46478 159200 46534 160000
rect 48042 159200 48098 160000
rect 49606 159200 49662 160000
rect 51262 159200 51318 160000
rect 52826 159200 52882 160000
rect 54390 159200 54446 160000
rect 55954 159200 56010 160000
rect 57518 159200 57574 160000
rect 59082 159200 59138 160000
rect 60738 159200 60794 160000
rect 62302 159200 62358 160000
rect 63866 159200 63922 160000
rect 65430 159200 65486 160000
rect 66994 159200 67050 160000
rect 68558 159200 68614 160000
rect 70122 159200 70178 160000
rect 71778 159200 71834 160000
rect 73342 159200 73398 160000
rect 74906 159200 74962 160000
rect 76470 159200 76526 160000
rect 78034 159200 78090 160000
rect 79598 159200 79654 160000
rect 81254 159200 81310 160000
rect 82818 159200 82874 160000
rect 84382 159200 84438 160000
rect 85946 159200 86002 160000
rect 87510 159200 87566 160000
rect 89074 159200 89130 160000
rect 90730 159200 90786 160000
rect 92294 159200 92350 160000
rect 93858 159200 93914 160000
rect 95422 159200 95478 160000
rect 96986 159200 97042 160000
rect 98550 159200 98606 160000
rect 100114 159200 100170 160000
rect 101770 159200 101826 160000
rect 103334 159200 103390 160000
rect 104898 159200 104954 160000
rect 106462 159200 106518 160000
rect 108026 159200 108082 160000
rect 109590 159200 109646 160000
rect 111246 159200 111302 160000
rect 112810 159200 112866 160000
rect 114374 159200 114430 160000
rect 115938 159200 115994 160000
rect 117502 159200 117558 160000
rect 119066 159200 119122 160000
rect 1030 0 1086 800
rect 3146 0 3202 800
rect 5262 0 5318 800
rect 7378 0 7434 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 16026 0 16082 800
rect 18142 0 18198 800
rect 20258 0 20314 800
rect 22374 0 22430 800
rect 24582 0 24638 800
rect 26698 0 26754 800
rect 28814 0 28870 800
rect 31022 0 31078 800
rect 33138 0 33194 800
rect 35254 0 35310 800
rect 37370 0 37426 800
rect 39578 0 39634 800
rect 41694 0 41750 800
rect 43810 0 43866 800
rect 46018 0 46074 800
rect 48134 0 48190 800
rect 50250 0 50306 800
rect 52366 0 52422 800
rect 54574 0 54630 800
rect 56690 0 56746 800
rect 58806 0 58862 800
rect 61014 0 61070 800
rect 63130 0 63186 800
rect 65246 0 65302 800
rect 67362 0 67418 800
rect 69570 0 69626 800
rect 71686 0 71742 800
rect 73802 0 73858 800
rect 76010 0 76066 800
rect 78126 0 78182 800
rect 80242 0 80298 800
rect 82358 0 82414 800
rect 84566 0 84622 800
rect 86682 0 86738 800
rect 88798 0 88854 800
rect 91006 0 91062 800
rect 93122 0 93178 800
rect 95238 0 95294 800
rect 97354 0 97410 800
rect 99562 0 99618 800
rect 101678 0 101734 800
rect 103794 0 103850 800
rect 106002 0 106058 800
rect 108118 0 108174 800
rect 110234 0 110290 800
rect 112350 0 112406 800
rect 114558 0 114614 800
rect 116674 0 116730 800
rect 118790 0 118846 800
<< obsm2 >>
rect 1032 159144 2262 159338
rect 2430 159144 3826 159338
rect 3994 159144 5390 159338
rect 5558 159144 6954 159338
rect 7122 159144 8518 159338
rect 8686 159144 10082 159338
rect 10250 159144 11738 159338
rect 11906 159144 13302 159338
rect 13470 159144 14866 159338
rect 15034 159144 16430 159338
rect 16598 159144 17994 159338
rect 18162 159144 19558 159338
rect 19726 159144 21214 159338
rect 21382 159144 22778 159338
rect 22946 159144 24342 159338
rect 24510 159144 25906 159338
rect 26074 159144 27470 159338
rect 27638 159144 29034 159338
rect 29202 159144 30690 159338
rect 30858 159144 32254 159338
rect 32422 159144 33818 159338
rect 33986 159144 35382 159338
rect 35550 159144 36946 159338
rect 37114 159144 38510 159338
rect 38678 159144 40074 159338
rect 40242 159144 41730 159338
rect 41898 159144 43294 159338
rect 43462 159144 44858 159338
rect 45026 159144 46422 159338
rect 46590 159144 47986 159338
rect 48154 159144 49550 159338
rect 49718 159144 51206 159338
rect 51374 159144 52770 159338
rect 52938 159144 54334 159338
rect 54502 159144 55898 159338
rect 56066 159144 57462 159338
rect 57630 159144 59026 159338
rect 59194 159144 60682 159338
rect 60850 159144 62246 159338
rect 62414 159144 63810 159338
rect 63978 159144 65374 159338
rect 65542 159144 66938 159338
rect 67106 159144 68502 159338
rect 68670 159144 70066 159338
rect 70234 159144 71722 159338
rect 71890 159144 73286 159338
rect 73454 159144 74850 159338
rect 75018 159144 76414 159338
rect 76582 159144 77978 159338
rect 78146 159144 79542 159338
rect 79710 159144 81198 159338
rect 81366 159144 82762 159338
rect 82930 159144 84326 159338
rect 84494 159144 85890 159338
rect 86058 159144 87454 159338
rect 87622 159144 89018 159338
rect 89186 159144 90674 159338
rect 90842 159144 92238 159338
rect 92406 159144 93802 159338
rect 93970 159144 95366 159338
rect 95534 159144 96930 159338
rect 97098 159144 98494 159338
rect 98662 159144 100058 159338
rect 100226 159144 101714 159338
rect 101882 159144 103278 159338
rect 103446 159144 104842 159338
rect 105010 159144 106406 159338
rect 106574 159144 107970 159338
rect 108138 159144 109534 159338
rect 109702 159144 111190 159338
rect 111358 159144 112754 159338
rect 112922 159144 114318 159338
rect 114486 159144 115882 159338
rect 116050 159144 117446 159338
rect 117614 159144 119010 159338
rect 1032 856 119120 159144
rect 1142 711 3090 856
rect 3258 711 5206 856
rect 5374 711 7322 856
rect 7490 711 9530 856
rect 9698 711 11646 856
rect 11814 711 13762 856
rect 13930 711 15970 856
rect 16138 711 18086 856
rect 18254 711 20202 856
rect 20370 711 22318 856
rect 22486 711 24526 856
rect 24694 711 26642 856
rect 26810 711 28758 856
rect 28926 711 30966 856
rect 31134 711 33082 856
rect 33250 711 35198 856
rect 35366 711 37314 856
rect 37482 711 39522 856
rect 39690 711 41638 856
rect 41806 711 43754 856
rect 43922 711 45962 856
rect 46130 711 48078 856
rect 48246 711 50194 856
rect 50362 711 52310 856
rect 52478 711 54518 856
rect 54686 711 56634 856
rect 56802 711 58750 856
rect 58918 711 60958 856
rect 61126 711 63074 856
rect 63242 711 65190 856
rect 65358 711 67306 856
rect 67474 711 69514 856
rect 69682 711 71630 856
rect 71798 711 73746 856
rect 73914 711 75954 856
rect 76122 711 78070 856
rect 78238 711 80186 856
rect 80354 711 82302 856
rect 82470 711 84510 856
rect 84678 711 86626 856
rect 86794 711 88742 856
rect 88910 711 90950 856
rect 91118 711 93066 856
rect 93234 711 95182 856
rect 95350 711 97298 856
rect 97466 711 99506 856
rect 99674 711 101622 856
rect 101790 711 103738 856
rect 103906 711 105946 856
rect 106114 711 108062 856
rect 108230 711 110178 856
rect 110346 711 112294 856
rect 112462 711 114502 856
rect 114670 711 116618 856
rect 116786 711 118734 856
rect 118902 711 119120 856
<< metal3 >>
rect 0 158992 800 159112
rect 0 157360 800 157480
rect 0 155728 800 155848
rect 0 154096 800 154216
rect 0 152600 800 152720
rect 0 150968 800 151088
rect 0 149336 800 149456
rect 0 147704 800 147824
rect 119200 146616 120000 146736
rect 0 146208 800 146328
rect 0 144576 800 144696
rect 0 142944 800 143064
rect 0 141312 800 141432
rect 0 139816 800 139936
rect 0 138184 800 138304
rect 0 136552 800 136672
rect 0 134920 800 135040
rect 0 133424 800 133544
rect 0 131792 800 131912
rect 0 130160 800 130280
rect 0 128528 800 128648
rect 0 127032 800 127152
rect 0 125400 800 125520
rect 0 123768 800 123888
rect 0 122136 800 122256
rect 0 120640 800 120760
rect 119200 119960 120000 120080
rect 0 119008 800 119128
rect 0 117376 800 117496
rect 0 115744 800 115864
rect 0 114112 800 114232
rect 0 112616 800 112736
rect 0 110984 800 111104
rect 0 109352 800 109472
rect 0 107720 800 107840
rect 0 106224 800 106344
rect 0 104592 800 104712
rect 0 102960 800 103080
rect 0 101328 800 101448
rect 0 99832 800 99952
rect 0 98200 800 98320
rect 0 96568 800 96688
rect 0 94936 800 95056
rect 0 93440 800 93560
rect 119200 93304 120000 93424
rect 0 91808 800 91928
rect 0 90176 800 90296
rect 0 88544 800 88664
rect 0 87048 800 87168
rect 0 85416 800 85536
rect 0 83784 800 83904
rect 0 82152 800 82272
rect 0 80656 800 80776
rect 0 79024 800 79144
rect 0 77392 800 77512
rect 0 75760 800 75880
rect 0 74128 800 74248
rect 0 72632 800 72752
rect 0 71000 800 71120
rect 0 69368 800 69488
rect 0 67736 800 67856
rect 119200 66648 120000 66768
rect 0 66240 800 66360
rect 0 64608 800 64728
rect 0 62976 800 63096
rect 0 61344 800 61464
rect 0 59848 800 59968
rect 0 58216 800 58336
rect 0 56584 800 56704
rect 0 54952 800 55072
rect 0 53456 800 53576
rect 0 51824 800 51944
rect 0 50192 800 50312
rect 0 48560 800 48680
rect 0 47064 800 47184
rect 0 45432 800 45552
rect 0 43800 800 43920
rect 0 42168 800 42288
rect 0 40672 800 40792
rect 119200 39992 120000 40112
rect 0 39040 800 39160
rect 0 37408 800 37528
rect 0 35776 800 35896
rect 0 34144 800 34264
rect 0 32648 800 32768
rect 0 31016 800 31136
rect 0 29384 800 29504
rect 0 27752 800 27872
rect 0 26256 800 26376
rect 0 24624 800 24744
rect 0 22992 800 23112
rect 0 21360 800 21480
rect 0 19864 800 19984
rect 0 18232 800 18352
rect 0 16600 800 16720
rect 0 14968 800 15088
rect 0 13472 800 13592
rect 119200 13336 120000 13456
rect 0 11840 800 11960
rect 0 10208 800 10328
rect 0 8576 800 8696
rect 0 7080 800 7200
rect 0 5448 800 5568
rect 0 3816 800 3936
rect 0 2184 800 2304
rect 0 688 800 808
<< obsm3 >>
rect 880 158912 119200 159085
rect 800 157560 119200 158912
rect 880 157280 119200 157560
rect 800 155928 119200 157280
rect 880 155648 119200 155928
rect 800 154296 119200 155648
rect 880 154016 119200 154296
rect 800 152800 119200 154016
rect 880 152520 119200 152800
rect 800 151168 119200 152520
rect 880 150888 119200 151168
rect 800 149536 119200 150888
rect 880 149256 119200 149536
rect 800 147904 119200 149256
rect 880 147624 119200 147904
rect 800 146816 119200 147624
rect 800 146536 119120 146816
rect 800 146408 119200 146536
rect 880 146128 119200 146408
rect 800 144776 119200 146128
rect 880 144496 119200 144776
rect 800 143144 119200 144496
rect 880 142864 119200 143144
rect 800 141512 119200 142864
rect 880 141232 119200 141512
rect 800 140016 119200 141232
rect 880 139736 119200 140016
rect 800 138384 119200 139736
rect 880 138104 119200 138384
rect 800 136752 119200 138104
rect 880 136472 119200 136752
rect 800 135120 119200 136472
rect 880 134840 119200 135120
rect 800 133624 119200 134840
rect 880 133344 119200 133624
rect 800 131992 119200 133344
rect 880 131712 119200 131992
rect 800 130360 119200 131712
rect 880 130080 119200 130360
rect 800 128728 119200 130080
rect 880 128448 119200 128728
rect 800 127232 119200 128448
rect 880 126952 119200 127232
rect 800 125600 119200 126952
rect 880 125320 119200 125600
rect 800 123968 119200 125320
rect 880 123688 119200 123968
rect 800 122336 119200 123688
rect 880 122056 119200 122336
rect 800 120840 119200 122056
rect 880 120560 119200 120840
rect 800 120160 119200 120560
rect 800 119880 119120 120160
rect 800 119208 119200 119880
rect 880 118928 119200 119208
rect 800 117576 119200 118928
rect 880 117296 119200 117576
rect 800 115944 119200 117296
rect 880 115664 119200 115944
rect 800 114312 119200 115664
rect 880 114032 119200 114312
rect 800 112816 119200 114032
rect 880 112536 119200 112816
rect 800 111184 119200 112536
rect 880 110904 119200 111184
rect 800 109552 119200 110904
rect 880 109272 119200 109552
rect 800 107920 119200 109272
rect 880 107640 119200 107920
rect 800 106424 119200 107640
rect 880 106144 119200 106424
rect 800 104792 119200 106144
rect 880 104512 119200 104792
rect 800 103160 119200 104512
rect 880 102880 119200 103160
rect 800 101528 119200 102880
rect 880 101248 119200 101528
rect 800 100032 119200 101248
rect 880 99752 119200 100032
rect 800 98400 119200 99752
rect 880 98120 119200 98400
rect 800 96768 119200 98120
rect 880 96488 119200 96768
rect 800 95136 119200 96488
rect 880 94856 119200 95136
rect 800 93640 119200 94856
rect 880 93504 119200 93640
rect 880 93360 119120 93504
rect 800 93224 119120 93360
rect 800 92008 119200 93224
rect 880 91728 119200 92008
rect 800 90376 119200 91728
rect 880 90096 119200 90376
rect 800 88744 119200 90096
rect 880 88464 119200 88744
rect 800 87248 119200 88464
rect 880 86968 119200 87248
rect 800 85616 119200 86968
rect 880 85336 119200 85616
rect 800 83984 119200 85336
rect 880 83704 119200 83984
rect 800 82352 119200 83704
rect 880 82072 119200 82352
rect 800 80856 119200 82072
rect 880 80576 119200 80856
rect 800 79224 119200 80576
rect 880 78944 119200 79224
rect 800 77592 119200 78944
rect 880 77312 119200 77592
rect 800 75960 119200 77312
rect 880 75680 119200 75960
rect 800 74328 119200 75680
rect 880 74048 119200 74328
rect 800 72832 119200 74048
rect 880 72552 119200 72832
rect 800 71200 119200 72552
rect 880 70920 119200 71200
rect 800 69568 119200 70920
rect 880 69288 119200 69568
rect 800 67936 119200 69288
rect 880 67656 119200 67936
rect 800 66848 119200 67656
rect 800 66568 119120 66848
rect 800 66440 119200 66568
rect 880 66160 119200 66440
rect 800 64808 119200 66160
rect 880 64528 119200 64808
rect 800 63176 119200 64528
rect 880 62896 119200 63176
rect 800 61544 119200 62896
rect 880 61264 119200 61544
rect 800 60048 119200 61264
rect 880 59768 119200 60048
rect 800 58416 119200 59768
rect 880 58136 119200 58416
rect 800 56784 119200 58136
rect 880 56504 119200 56784
rect 800 55152 119200 56504
rect 880 54872 119200 55152
rect 800 53656 119200 54872
rect 880 53376 119200 53656
rect 800 52024 119200 53376
rect 880 51744 119200 52024
rect 800 50392 119200 51744
rect 880 50112 119200 50392
rect 800 48760 119200 50112
rect 880 48480 119200 48760
rect 800 47264 119200 48480
rect 880 46984 119200 47264
rect 800 45632 119200 46984
rect 880 45352 119200 45632
rect 800 44000 119200 45352
rect 880 43720 119200 44000
rect 800 42368 119200 43720
rect 880 42088 119200 42368
rect 800 40872 119200 42088
rect 880 40592 119200 40872
rect 800 40192 119200 40592
rect 800 39912 119120 40192
rect 800 39240 119200 39912
rect 880 38960 119200 39240
rect 800 37608 119200 38960
rect 880 37328 119200 37608
rect 800 35976 119200 37328
rect 880 35696 119200 35976
rect 800 34344 119200 35696
rect 880 34064 119200 34344
rect 800 32848 119200 34064
rect 880 32568 119200 32848
rect 800 31216 119200 32568
rect 880 30936 119200 31216
rect 800 29584 119200 30936
rect 880 29304 119200 29584
rect 800 27952 119200 29304
rect 880 27672 119200 27952
rect 800 26456 119200 27672
rect 880 26176 119200 26456
rect 800 24824 119200 26176
rect 880 24544 119200 24824
rect 800 23192 119200 24544
rect 880 22912 119200 23192
rect 800 21560 119200 22912
rect 880 21280 119200 21560
rect 800 20064 119200 21280
rect 880 19784 119200 20064
rect 800 18432 119200 19784
rect 880 18152 119200 18432
rect 800 16800 119200 18152
rect 880 16520 119200 16800
rect 800 15168 119200 16520
rect 880 14888 119200 15168
rect 800 13672 119200 14888
rect 880 13536 119200 13672
rect 880 13392 119120 13536
rect 800 13256 119120 13392
rect 800 12040 119200 13256
rect 880 11760 119200 12040
rect 800 10408 119200 11760
rect 880 10128 119200 10408
rect 800 8776 119200 10128
rect 880 8496 119200 8776
rect 800 7280 119200 8496
rect 880 7000 119200 7280
rect 800 5648 119200 7000
rect 880 5368 119200 5648
rect 800 4016 119200 5368
rect 880 3736 119200 4016
rect 800 2384 119200 3736
rect 880 2104 119200 2384
rect 800 888 119200 2104
rect 880 715 119200 888
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
<< obsm4 >>
rect 3371 3979 4128 156093
rect 4608 3979 19488 156093
rect 19968 3979 34848 156093
rect 35328 3979 50208 156093
rect 50688 3979 65568 156093
rect 66048 3979 80928 156093
rect 81408 3979 96288 156093
rect 96768 3979 111648 156093
rect 112128 3979 116229 156093
<< labels >>
rlabel metal2 s 86682 0 86738 800 6 flash_csb
port 1 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 flash_io0_read
port 2 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 flash_io0_we
port 3 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 flash_io0_write
port 4 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 flash_io1_read
port 5 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 flash_io1_we
port 6 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 flash_io1_write
port 7 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 flash_sck
port 8 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 internal_uart_rx
port 9 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 internal_uart_tx
port 10 nsew signal output
rlabel metal2 s 754 159200 810 160000 6 io_in[0]
port 11 nsew signal input
rlabel metal2 s 16486 159200 16542 160000 6 io_in[10]
port 12 nsew signal input
rlabel metal2 s 18050 159200 18106 160000 6 io_in[11]
port 13 nsew signal input
rlabel metal2 s 19614 159200 19670 160000 6 io_in[12]
port 14 nsew signal input
rlabel metal2 s 21270 159200 21326 160000 6 io_in[13]
port 15 nsew signal input
rlabel metal2 s 22834 159200 22890 160000 6 io_in[14]
port 16 nsew signal input
rlabel metal2 s 24398 159200 24454 160000 6 io_in[15]
port 17 nsew signal input
rlabel metal2 s 25962 159200 26018 160000 6 io_in[16]
port 18 nsew signal input
rlabel metal2 s 27526 159200 27582 160000 6 io_in[17]
port 19 nsew signal input
rlabel metal2 s 29090 159200 29146 160000 6 io_in[18]
port 20 nsew signal input
rlabel metal2 s 30746 159200 30802 160000 6 io_in[19]
port 21 nsew signal input
rlabel metal2 s 2318 159200 2374 160000 6 io_in[1]
port 22 nsew signal input
rlabel metal2 s 32310 159200 32366 160000 6 io_in[20]
port 23 nsew signal input
rlabel metal2 s 33874 159200 33930 160000 6 io_in[21]
port 24 nsew signal input
rlabel metal2 s 35438 159200 35494 160000 6 io_in[22]
port 25 nsew signal input
rlabel metal2 s 37002 159200 37058 160000 6 io_in[23]
port 26 nsew signal input
rlabel metal2 s 38566 159200 38622 160000 6 io_in[24]
port 27 nsew signal input
rlabel metal2 s 40130 159200 40186 160000 6 io_in[25]
port 28 nsew signal input
rlabel metal2 s 41786 159200 41842 160000 6 io_in[26]
port 29 nsew signal input
rlabel metal2 s 43350 159200 43406 160000 6 io_in[27]
port 30 nsew signal input
rlabel metal2 s 44914 159200 44970 160000 6 io_in[28]
port 31 nsew signal input
rlabel metal2 s 46478 159200 46534 160000 6 io_in[29]
port 32 nsew signal input
rlabel metal2 s 3882 159200 3938 160000 6 io_in[2]
port 33 nsew signal input
rlabel metal2 s 48042 159200 48098 160000 6 io_in[30]
port 34 nsew signal input
rlabel metal2 s 49606 159200 49662 160000 6 io_in[31]
port 35 nsew signal input
rlabel metal2 s 51262 159200 51318 160000 6 io_in[32]
port 36 nsew signal input
rlabel metal2 s 52826 159200 52882 160000 6 io_in[33]
port 37 nsew signal input
rlabel metal2 s 54390 159200 54446 160000 6 io_in[34]
port 38 nsew signal input
rlabel metal2 s 55954 159200 56010 160000 6 io_in[35]
port 39 nsew signal input
rlabel metal2 s 57518 159200 57574 160000 6 io_in[36]
port 40 nsew signal input
rlabel metal2 s 59082 159200 59138 160000 6 io_in[37]
port 41 nsew signal input
rlabel metal2 s 5446 159200 5502 160000 6 io_in[3]
port 42 nsew signal input
rlabel metal2 s 7010 159200 7066 160000 6 io_in[4]
port 43 nsew signal input
rlabel metal2 s 8574 159200 8630 160000 6 io_in[5]
port 44 nsew signal input
rlabel metal2 s 10138 159200 10194 160000 6 io_in[6]
port 45 nsew signal input
rlabel metal2 s 11794 159200 11850 160000 6 io_in[7]
port 46 nsew signal input
rlabel metal2 s 13358 159200 13414 160000 6 io_in[8]
port 47 nsew signal input
rlabel metal2 s 14922 159200 14978 160000 6 io_in[9]
port 48 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 io_oeb[0]
port 49 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 io_oeb[10]
port 50 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 io_oeb[11]
port 51 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 io_oeb[12]
port 52 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 io_oeb[13]
port 53 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 io_oeb[14]
port 54 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 io_oeb[15]
port 55 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 io_oeb[16]
port 56 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 io_oeb[17]
port 57 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 io_oeb[18]
port 58 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 io_oeb[19]
port 59 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 io_oeb[1]
port 60 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 io_oeb[20]
port 61 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 io_oeb[21]
port 62 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 io_oeb[22]
port 63 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 io_oeb[23]
port 64 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 io_oeb[24]
port 65 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 io_oeb[25]
port 66 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 io_oeb[26]
port 67 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 io_oeb[27]
port 68 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 io_oeb[28]
port 69 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 io_oeb[29]
port 70 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 io_oeb[2]
port 71 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 io_oeb[30]
port 72 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 io_oeb[31]
port 73 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 io_oeb[32]
port 74 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 io_oeb[33]
port 75 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 io_oeb[34]
port 76 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 io_oeb[35]
port 77 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 io_oeb[36]
port 78 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 io_oeb[37]
port 79 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 io_oeb[3]
port 80 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 io_oeb[4]
port 81 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 io_oeb[5]
port 82 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 io_oeb[6]
port 83 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 io_oeb[7]
port 84 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 io_oeb[8]
port 85 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 60738 159200 60794 160000 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 76470 159200 76526 160000 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 78034 159200 78090 160000 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 79598 159200 79654 160000 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 81254 159200 81310 160000 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 82818 159200 82874 160000 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 84382 159200 84438 160000 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 85946 159200 86002 160000 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 87510 159200 87566 160000 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 89074 159200 89130 160000 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 90730 159200 90786 160000 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 62302 159200 62358 160000 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 92294 159200 92350 160000 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 93858 159200 93914 160000 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 95422 159200 95478 160000 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 96986 159200 97042 160000 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 98550 159200 98606 160000 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 100114 159200 100170 160000 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 101770 159200 101826 160000 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 103334 159200 103390 160000 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 104898 159200 104954 160000 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 106462 159200 106518 160000 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 63866 159200 63922 160000 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 108026 159200 108082 160000 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 109590 159200 109646 160000 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 111246 159200 111302 160000 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 112810 159200 112866 160000 6 io_out[33]
port 113 nsew signal output
rlabel metal2 s 114374 159200 114430 160000 6 io_out[34]
port 114 nsew signal output
rlabel metal2 s 115938 159200 115994 160000 6 io_out[35]
port 115 nsew signal output
rlabel metal2 s 117502 159200 117558 160000 6 io_out[36]
port 116 nsew signal output
rlabel metal2 s 119066 159200 119122 160000 6 io_out[37]
port 117 nsew signal output
rlabel metal2 s 65430 159200 65486 160000 6 io_out[3]
port 118 nsew signal output
rlabel metal2 s 66994 159200 67050 160000 6 io_out[4]
port 119 nsew signal output
rlabel metal2 s 68558 159200 68614 160000 6 io_out[5]
port 120 nsew signal output
rlabel metal2 s 70122 159200 70178 160000 6 io_out[6]
port 121 nsew signal output
rlabel metal2 s 71778 159200 71834 160000 6 io_out[7]
port 122 nsew signal output
rlabel metal2 s 73342 159200 73398 160000 6 io_out[8]
port 123 nsew signal output
rlabel metal2 s 74906 159200 74962 160000 6 io_out[9]
port 124 nsew signal output
rlabel metal3 s 119200 66648 120000 66768 6 jtag_tck
port 125 nsew signal output
rlabel metal3 s 119200 93304 120000 93424 6 jtag_tdi
port 126 nsew signal output
rlabel metal3 s 119200 119960 120000 120080 6 jtag_tdo
port 127 nsew signal input
rlabel metal3 s 119200 146616 120000 146736 6 jtag_tms
port 128 nsew signal output
rlabel metal3 s 119200 13336 120000 13456 6 probe_blink[0]
port 129 nsew signal output
rlabel metal3 s 119200 39992 120000 40112 6 probe_blink[1]
port 130 nsew signal output
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 131 nsew power input
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 131 nsew power input
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 131 nsew power input
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 131 nsew power input
rlabel metal2 s 108118 0 108174 800 6 vga_b[0]
port 132 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 vga_b[1]
port 133 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 vga_g[0]
port 134 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 vga_g[1]
port 135 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 vga_hsync
port 136 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 vga_r[0]
port 137 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 vga_r[1]
port 138 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 vga_vsync
port 139 nsew signal input
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 140 nsew ground input
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 140 nsew ground input
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 140 nsew ground input
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 140 nsew ground input
rlabel metal3 s 0 688 800 808 6 wb_ack_o
port 141 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 wb_adr_i[0]
port 142 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 wb_adr_i[10]
port 143 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 wb_adr_i[11]
port 144 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 wb_adr_i[12]
port 145 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 wb_adr_i[13]
port 146 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 wb_adr_i[14]
port 147 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 wb_adr_i[15]
port 148 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 wb_adr_i[16]
port 149 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 wb_adr_i[17]
port 150 nsew signal input
rlabel metal3 s 0 106224 800 106344 6 wb_adr_i[18]
port 151 nsew signal input
rlabel metal3 s 0 110984 800 111104 6 wb_adr_i[19]
port 152 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 wb_adr_i[1]
port 153 nsew signal input
rlabel metal3 s 0 115744 800 115864 6 wb_adr_i[20]
port 154 nsew signal input
rlabel metal3 s 0 120640 800 120760 6 wb_adr_i[21]
port 155 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 wb_adr_i[22]
port 156 nsew signal input
rlabel metal3 s 0 130160 800 130280 6 wb_adr_i[23]
port 157 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 wb_adr_i[2]
port 158 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 wb_adr_i[3]
port 159 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 wb_adr_i[4]
port 160 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 wb_adr_i[5]
port 161 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 wb_adr_i[6]
port 162 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 wb_adr_i[7]
port 163 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 wb_adr_i[8]
port 164 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 wb_adr_i[9]
port 165 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wb_clk_i
port 166 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 wb_cyc_i
port 167 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 wb_data_i[0]
port 168 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 wb_data_i[10]
port 169 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 wb_data_i[11]
port 170 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 wb_data_i[12]
port 171 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 wb_data_i[13]
port 172 nsew signal input
rlabel metal3 s 0 88544 800 88664 6 wb_data_i[14]
port 173 nsew signal input
rlabel metal3 s 0 93440 800 93560 6 wb_data_i[15]
port 174 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 wb_data_i[16]
port 175 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 wb_data_i[17]
port 176 nsew signal input
rlabel metal3 s 0 107720 800 107840 6 wb_data_i[18]
port 177 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 wb_data_i[19]
port 178 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 wb_data_i[1]
port 179 nsew signal input
rlabel metal3 s 0 117376 800 117496 6 wb_data_i[20]
port 180 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 wb_data_i[21]
port 181 nsew signal input
rlabel metal3 s 0 127032 800 127152 6 wb_data_i[22]
port 182 nsew signal input
rlabel metal3 s 0 131792 800 131912 6 wb_data_i[23]
port 183 nsew signal input
rlabel metal3 s 0 134920 800 135040 6 wb_data_i[24]
port 184 nsew signal input
rlabel metal3 s 0 138184 800 138304 6 wb_data_i[25]
port 185 nsew signal input
rlabel metal3 s 0 141312 800 141432 6 wb_data_i[26]
port 186 nsew signal input
rlabel metal3 s 0 144576 800 144696 6 wb_data_i[27]
port 187 nsew signal input
rlabel metal3 s 0 147704 800 147824 6 wb_data_i[28]
port 188 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 wb_data_i[29]
port 189 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 wb_data_i[2]
port 190 nsew signal input
rlabel metal3 s 0 154096 800 154216 6 wb_data_i[30]
port 191 nsew signal input
rlabel metal3 s 0 157360 800 157480 6 wb_data_i[31]
port 192 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wb_data_i[3]
port 193 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 wb_data_i[4]
port 194 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 wb_data_i[5]
port 195 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 wb_data_i[6]
port 196 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 wb_data_i[7]
port 197 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 wb_data_i[8]
port 198 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 wb_data_i[9]
port 199 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 wb_data_o[0]
port 200 nsew signal output
rlabel metal3 s 0 71000 800 71120 6 wb_data_o[10]
port 201 nsew signal output
rlabel metal3 s 0 75760 800 75880 6 wb_data_o[11]
port 202 nsew signal output
rlabel metal3 s 0 80656 800 80776 6 wb_data_o[12]
port 203 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 wb_data_o[13]
port 204 nsew signal output
rlabel metal3 s 0 90176 800 90296 6 wb_data_o[14]
port 205 nsew signal output
rlabel metal3 s 0 94936 800 95056 6 wb_data_o[15]
port 206 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 wb_data_o[16]
port 207 nsew signal output
rlabel metal3 s 0 104592 800 104712 6 wb_data_o[17]
port 208 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 wb_data_o[18]
port 209 nsew signal output
rlabel metal3 s 0 114112 800 114232 6 wb_data_o[19]
port 210 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 wb_data_o[1]
port 211 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 wb_data_o[20]
port 212 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 wb_data_o[21]
port 213 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 wb_data_o[22]
port 214 nsew signal output
rlabel metal3 s 0 133424 800 133544 6 wb_data_o[23]
port 215 nsew signal output
rlabel metal3 s 0 136552 800 136672 6 wb_data_o[24]
port 216 nsew signal output
rlabel metal3 s 0 139816 800 139936 6 wb_data_o[25]
port 217 nsew signal output
rlabel metal3 s 0 142944 800 143064 6 wb_data_o[26]
port 218 nsew signal output
rlabel metal3 s 0 146208 800 146328 6 wb_data_o[27]
port 219 nsew signal output
rlabel metal3 s 0 149336 800 149456 6 wb_data_o[28]
port 220 nsew signal output
rlabel metal3 s 0 152600 800 152720 6 wb_data_o[29]
port 221 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 wb_data_o[2]
port 222 nsew signal output
rlabel metal3 s 0 155728 800 155848 6 wb_data_o[30]
port 223 nsew signal output
rlabel metal3 s 0 158992 800 159112 6 wb_data_o[31]
port 224 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 wb_data_o[3]
port 225 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 wb_data_o[4]
port 226 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 wb_data_o[5]
port 227 nsew signal output
rlabel metal3 s 0 51824 800 51944 6 wb_data_o[6]
port 228 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 wb_data_o[7]
port 229 nsew signal output
rlabel metal3 s 0 61344 800 61464 6 wb_data_o[8]
port 230 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 wb_data_o[9]
port 231 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 wb_error_o
port 232 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 wb_rst_i
port 233 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 wb_sel_i[0]
port 234 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 wb_sel_i[1]
port 235 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 wb_sel_i[2]
port 236 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 wb_sel_i[3]
port 237 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 wb_stall_o
port 238 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 wb_stb_i
port 239 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 wb_we_i
port 240 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 50598442
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripherals_Flat/runs/Peripherals_Flat/results/finishing/Peripherals.magic.gds
string GDS_START 1119466
<< end >>

