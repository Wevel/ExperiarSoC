VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Video
  CLASS BLOCK ;
  FOREIGN Video ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 500.000 ;
  PIN sram0_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END sram0_addr0[0]
  PIN sram0_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END sram0_addr0[1]
  PIN sram0_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END sram0_addr0[2]
  PIN sram0_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END sram0_addr0[3]
  PIN sram0_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END sram0_addr0[4]
  PIN sram0_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END sram0_addr0[5]
  PIN sram0_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END sram0_addr0[6]
  PIN sram0_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END sram0_addr0[7]
  PIN sram0_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END sram0_addr0[8]
  PIN sram0_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END sram0_addr1[0]
  PIN sram0_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END sram0_addr1[1]
  PIN sram0_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END sram0_addr1[2]
  PIN sram0_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END sram0_addr1[3]
  PIN sram0_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END sram0_addr1[4]
  PIN sram0_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END sram0_addr1[5]
  PIN sram0_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END sram0_addr1[6]
  PIN sram0_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END sram0_addr1[7]
  PIN sram0_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END sram0_addr1[8]
  PIN sram0_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END sram0_clk0
  PIN sram0_clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END sram0_clk1
  PIN sram0_csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END sram0_csb0[0]
  PIN sram0_csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END sram0_csb0[1]
  PIN sram0_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END sram0_csb1[0]
  PIN sram0_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END sram0_csb1[1]
  PIN sram0_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END sram0_din0[0]
  PIN sram0_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END sram0_din0[10]
  PIN sram0_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END sram0_din0[11]
  PIN sram0_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END sram0_din0[12]
  PIN sram0_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END sram0_din0[13]
  PIN sram0_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END sram0_din0[14]
  PIN sram0_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END sram0_din0[15]
  PIN sram0_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END sram0_din0[16]
  PIN sram0_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END sram0_din0[17]
  PIN sram0_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END sram0_din0[18]
  PIN sram0_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END sram0_din0[19]
  PIN sram0_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END sram0_din0[1]
  PIN sram0_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END sram0_din0[20]
  PIN sram0_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END sram0_din0[21]
  PIN sram0_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END sram0_din0[22]
  PIN sram0_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END sram0_din0[23]
  PIN sram0_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END sram0_din0[24]
  PIN sram0_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END sram0_din0[25]
  PIN sram0_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END sram0_din0[26]
  PIN sram0_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END sram0_din0[27]
  PIN sram0_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END sram0_din0[28]
  PIN sram0_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END sram0_din0[29]
  PIN sram0_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END sram0_din0[2]
  PIN sram0_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END sram0_din0[30]
  PIN sram0_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END sram0_din0[31]
  PIN sram0_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END sram0_din0[3]
  PIN sram0_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END sram0_din0[4]
  PIN sram0_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END sram0_din0[5]
  PIN sram0_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END sram0_din0[6]
  PIN sram0_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END sram0_din0[7]
  PIN sram0_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END sram0_din0[8]
  PIN sram0_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END sram0_din0[9]
  PIN sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END sram0_dout0[0]
  PIN sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END sram0_dout0[10]
  PIN sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END sram0_dout0[11]
  PIN sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END sram0_dout0[12]
  PIN sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END sram0_dout0[13]
  PIN sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END sram0_dout0[14]
  PIN sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END sram0_dout0[15]
  PIN sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END sram0_dout0[16]
  PIN sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.080 4.000 376.680 ;
    END
  END sram0_dout0[17]
  PIN sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END sram0_dout0[18]
  PIN sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END sram0_dout0[19]
  PIN sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END sram0_dout0[1]
  PIN sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END sram0_dout0[20]
  PIN sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END sram0_dout0[21]
  PIN sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END sram0_dout0[22]
  PIN sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END sram0_dout0[23]
  PIN sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END sram0_dout0[24]
  PIN sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END sram0_dout0[25]
  PIN sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END sram0_dout0[26]
  PIN sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END sram0_dout0[27]
  PIN sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END sram0_dout0[28]
  PIN sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END sram0_dout0[29]
  PIN sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END sram0_dout0[2]
  PIN sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END sram0_dout0[30]
  PIN sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END sram0_dout0[31]
  PIN sram0_dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END sram0_dout0[32]
  PIN sram0_dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END sram0_dout0[33]
  PIN sram0_dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.960 4.000 421.560 ;
    END
  END sram0_dout0[34]
  PIN sram0_dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END sram0_dout0[35]
  PIN sram0_dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.400 4.000 427.000 ;
    END
  END sram0_dout0[36]
  PIN sram0_dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END sram0_dout0[37]
  PIN sram0_dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END sram0_dout0[38]
  PIN sram0_dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END sram0_dout0[39]
  PIN sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END sram0_dout0[3]
  PIN sram0_dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END sram0_dout0[40]
  PIN sram0_dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END sram0_dout0[41]
  PIN sram0_dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END sram0_dout0[42]
  PIN sram0_dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END sram0_dout0[43]
  PIN sram0_dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END sram0_dout0[44]
  PIN sram0_dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END sram0_dout0[45]
  PIN sram0_dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END sram0_dout0[46]
  PIN sram0_dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.960 4.000 455.560 ;
    END
  END sram0_dout0[47]
  PIN sram0_dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END sram0_dout0[48]
  PIN sram0_dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 460.400 4.000 461.000 ;
    END
  END sram0_dout0[49]
  PIN sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END sram0_dout0[4]
  PIN sram0_dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END sram0_dout0[50]
  PIN sram0_dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END sram0_dout0[51]
  PIN sram0_dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END sram0_dout0[52]
  PIN sram0_dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END sram0_dout0[53]
  PIN sram0_dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END sram0_dout0[54]
  PIN sram0_dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END sram0_dout0[55]
  PIN sram0_dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END sram0_dout0[56]
  PIN sram0_dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END sram0_dout0[57]
  PIN sram0_dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END sram0_dout0[58]
  PIN sram0_dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END sram0_dout0[59]
  PIN sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END sram0_dout0[5]
  PIN sram0_dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END sram0_dout0[60]
  PIN sram0_dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END sram0_dout0[61]
  PIN sram0_dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END sram0_dout0[62]
  PIN sram0_dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END sram0_dout0[63]
  PIN sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END sram0_dout0[6]
  PIN sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END sram0_dout0[7]
  PIN sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END sram0_dout0[8]
  PIN sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END sram0_dout0[9]
  PIN sram0_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END sram0_dout1[0]
  PIN sram0_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END sram0_dout1[10]
  PIN sram0_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END sram0_dout1[11]
  PIN sram0_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END sram0_dout1[12]
  PIN sram0_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END sram0_dout1[13]
  PIN sram0_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END sram0_dout1[14]
  PIN sram0_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END sram0_dout1[15]
  PIN sram0_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END sram0_dout1[16]
  PIN sram0_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END sram0_dout1[17]
  PIN sram0_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END sram0_dout1[18]
  PIN sram0_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END sram0_dout1[19]
  PIN sram0_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END sram0_dout1[1]
  PIN sram0_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END sram0_dout1[20]
  PIN sram0_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END sram0_dout1[21]
  PIN sram0_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END sram0_dout1[22]
  PIN sram0_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END sram0_dout1[23]
  PIN sram0_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END sram0_dout1[24]
  PIN sram0_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END sram0_dout1[25]
  PIN sram0_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END sram0_dout1[26]
  PIN sram0_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END sram0_dout1[27]
  PIN sram0_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END sram0_dout1[28]
  PIN sram0_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END sram0_dout1[29]
  PIN sram0_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END sram0_dout1[2]
  PIN sram0_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END sram0_dout1[30]
  PIN sram0_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END sram0_dout1[31]
  PIN sram0_dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END sram0_dout1[32]
  PIN sram0_dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END sram0_dout1[33]
  PIN sram0_dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END sram0_dout1[34]
  PIN sram0_dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END sram0_dout1[35]
  PIN sram0_dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END sram0_dout1[36]
  PIN sram0_dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END sram0_dout1[37]
  PIN sram0_dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END sram0_dout1[38]
  PIN sram0_dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END sram0_dout1[39]
  PIN sram0_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END sram0_dout1[3]
  PIN sram0_dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END sram0_dout1[40]
  PIN sram0_dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END sram0_dout1[41]
  PIN sram0_dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END sram0_dout1[42]
  PIN sram0_dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END sram0_dout1[43]
  PIN sram0_dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END sram0_dout1[44]
  PIN sram0_dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END sram0_dout1[45]
  PIN sram0_dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END sram0_dout1[46]
  PIN sram0_dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END sram0_dout1[47]
  PIN sram0_dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END sram0_dout1[48]
  PIN sram0_dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END sram0_dout1[49]
  PIN sram0_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END sram0_dout1[4]
  PIN sram0_dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END sram0_dout1[50]
  PIN sram0_dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END sram0_dout1[51]
  PIN sram0_dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END sram0_dout1[52]
  PIN sram0_dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END sram0_dout1[53]
  PIN sram0_dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END sram0_dout1[54]
  PIN sram0_dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END sram0_dout1[55]
  PIN sram0_dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END sram0_dout1[56]
  PIN sram0_dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END sram0_dout1[57]
  PIN sram0_dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END sram0_dout1[58]
  PIN sram0_dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END sram0_dout1[59]
  PIN sram0_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END sram0_dout1[5]
  PIN sram0_dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END sram0_dout1[60]
  PIN sram0_dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END sram0_dout1[61]
  PIN sram0_dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END sram0_dout1[62]
  PIN sram0_dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END sram0_dout1[63]
  PIN sram0_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END sram0_dout1[6]
  PIN sram0_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END sram0_dout1[7]
  PIN sram0_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END sram0_dout1[8]
  PIN sram0_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END sram0_dout1[9]
  PIN sram0_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END sram0_web0
  PIN sram0_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END sram0_wmask0[0]
  PIN sram0_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END sram0_wmask0[1]
  PIN sram0_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END sram0_wmask0[2]
  PIN sram0_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END sram0_wmask0[3]
  PIN sram1_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 222.400 350.000 223.000 ;
    END
  END sram1_addr0[0]
  PIN sram1_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 225.120 350.000 225.720 ;
    END
  END sram1_addr0[1]
  PIN sram1_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 227.840 350.000 228.440 ;
    END
  END sram1_addr0[2]
  PIN sram1_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 230.560 350.000 231.160 ;
    END
  END sram1_addr0[3]
  PIN sram1_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 233.280 350.000 233.880 ;
    END
  END sram1_addr0[4]
  PIN sram1_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 236.000 350.000 236.600 ;
    END
  END sram1_addr0[5]
  PIN sram1_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 238.720 350.000 239.320 ;
    END
  END sram1_addr0[6]
  PIN sram1_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 240.760 350.000 241.360 ;
    END
  END sram1_addr0[7]
  PIN sram1_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 243.480 350.000 244.080 ;
    END
  END sram1_addr0[8]
  PIN sram1_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 8.200 350.000 8.800 ;
    END
  END sram1_addr1[0]
  PIN sram1_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 10.920 350.000 11.520 ;
    END
  END sram1_addr1[1]
  PIN sram1_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 13.640 350.000 14.240 ;
    END
  END sram1_addr1[2]
  PIN sram1_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 16.360 350.000 16.960 ;
    END
  END sram1_addr1[3]
  PIN sram1_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 19.080 350.000 19.680 ;
    END
  END sram1_addr1[4]
  PIN sram1_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 21.800 350.000 22.400 ;
    END
  END sram1_addr1[5]
  PIN sram1_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 24.520 350.000 25.120 ;
    END
  END sram1_addr1[6]
  PIN sram1_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 26.560 350.000 27.160 ;
    END
  END sram1_addr1[7]
  PIN sram1_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 29.280 350.000 29.880 ;
    END
  END sram1_addr1[8]
  PIN sram1_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 201.320 350.000 201.920 ;
    END
  END sram1_clk0
  PIN sram1_clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 0.720 350.000 1.320 ;
    END
  END sram1_clk1
  PIN sram1_csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 204.040 350.000 204.640 ;
    END
  END sram1_csb0[0]
  PIN sram1_csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 206.760 350.000 207.360 ;
    END
  END sram1_csb0[1]
  PIN sram1_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 2.760 350.000 3.360 ;
    END
  END sram1_csb1[0]
  PIN sram1_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 5.480 350.000 6.080 ;
    END
  END sram1_csb1[1]
  PIN sram1_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 246.200 350.000 246.800 ;
    END
  END sram1_din0[0]
  PIN sram1_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 272.720 350.000 273.320 ;
    END
  END sram1_din0[10]
  PIN sram1_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 275.440 350.000 276.040 ;
    END
  END sram1_din0[11]
  PIN sram1_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 278.160 350.000 278.760 ;
    END
  END sram1_din0[12]
  PIN sram1_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 280.880 350.000 281.480 ;
    END
  END sram1_din0[13]
  PIN sram1_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 283.600 350.000 284.200 ;
    END
  END sram1_din0[14]
  PIN sram1_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 286.320 350.000 286.920 ;
    END
  END sram1_din0[15]
  PIN sram1_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 288.360 350.000 288.960 ;
    END
  END sram1_din0[16]
  PIN sram1_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 291.080 350.000 291.680 ;
    END
  END sram1_din0[17]
  PIN sram1_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 293.800 350.000 294.400 ;
    END
  END sram1_din0[18]
  PIN sram1_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 296.520 350.000 297.120 ;
    END
  END sram1_din0[19]
  PIN sram1_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 248.920 350.000 249.520 ;
    END
  END sram1_din0[1]
  PIN sram1_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 299.240 350.000 299.840 ;
    END
  END sram1_din0[20]
  PIN sram1_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 301.960 350.000 302.560 ;
    END
  END sram1_din0[21]
  PIN sram1_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 304.680 350.000 305.280 ;
    END
  END sram1_din0[22]
  PIN sram1_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 307.400 350.000 308.000 ;
    END
  END sram1_din0[23]
  PIN sram1_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 310.120 350.000 310.720 ;
    END
  END sram1_din0[24]
  PIN sram1_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 312.160 350.000 312.760 ;
    END
  END sram1_din0[25]
  PIN sram1_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 314.880 350.000 315.480 ;
    END
  END sram1_din0[26]
  PIN sram1_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 317.600 350.000 318.200 ;
    END
  END sram1_din0[27]
  PIN sram1_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 320.320 350.000 320.920 ;
    END
  END sram1_din0[28]
  PIN sram1_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 323.040 350.000 323.640 ;
    END
  END sram1_din0[29]
  PIN sram1_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 251.640 350.000 252.240 ;
    END
  END sram1_din0[2]
  PIN sram1_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 325.760 350.000 326.360 ;
    END
  END sram1_din0[30]
  PIN sram1_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 328.480 350.000 329.080 ;
    END
  END sram1_din0[31]
  PIN sram1_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 254.360 350.000 254.960 ;
    END
  END sram1_din0[3]
  PIN sram1_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 257.080 350.000 257.680 ;
    END
  END sram1_din0[4]
  PIN sram1_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 259.800 350.000 260.400 ;
    END
  END sram1_din0[5]
  PIN sram1_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 262.520 350.000 263.120 ;
    END
  END sram1_din0[6]
  PIN sram1_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 264.560 350.000 265.160 ;
    END
  END sram1_din0[7]
  PIN sram1_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 267.280 350.000 267.880 ;
    END
  END sram1_din0[8]
  PIN sram1_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 270.000 350.000 270.600 ;
    END
  END sram1_din0[9]
  PIN sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 331.200 350.000 331.800 ;
    END
  END sram1_dout0[0]
  PIN sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 357.720 350.000 358.320 ;
    END
  END sram1_dout0[10]
  PIN sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 359.760 350.000 360.360 ;
    END
  END sram1_dout0[11]
  PIN sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 362.480 350.000 363.080 ;
    END
  END sram1_dout0[12]
  PIN sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 365.200 350.000 365.800 ;
    END
  END sram1_dout0[13]
  PIN sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 367.920 350.000 368.520 ;
    END
  END sram1_dout0[14]
  PIN sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 370.640 350.000 371.240 ;
    END
  END sram1_dout0[15]
  PIN sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 373.360 350.000 373.960 ;
    END
  END sram1_dout0[16]
  PIN sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 376.080 350.000 376.680 ;
    END
  END sram1_dout0[17]
  PIN sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 378.800 350.000 379.400 ;
    END
  END sram1_dout0[18]
  PIN sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 381.520 350.000 382.120 ;
    END
  END sram1_dout0[19]
  PIN sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 333.920 350.000 334.520 ;
    END
  END sram1_dout0[1]
  PIN sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 383.560 350.000 384.160 ;
    END
  END sram1_dout0[20]
  PIN sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 386.280 350.000 386.880 ;
    END
  END sram1_dout0[21]
  PIN sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 389.000 350.000 389.600 ;
    END
  END sram1_dout0[22]
  PIN sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 391.720 350.000 392.320 ;
    END
  END sram1_dout0[23]
  PIN sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 394.440 350.000 395.040 ;
    END
  END sram1_dout0[24]
  PIN sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 397.160 350.000 397.760 ;
    END
  END sram1_dout0[25]
  PIN sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 399.880 350.000 400.480 ;
    END
  END sram1_dout0[26]
  PIN sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 402.600 350.000 403.200 ;
    END
  END sram1_dout0[27]
  PIN sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 405.320 350.000 405.920 ;
    END
  END sram1_dout0[28]
  PIN sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 407.360 350.000 407.960 ;
    END
  END sram1_dout0[29]
  PIN sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 335.960 350.000 336.560 ;
    END
  END sram1_dout0[2]
  PIN sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 410.080 350.000 410.680 ;
    END
  END sram1_dout0[30]
  PIN sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 412.800 350.000 413.400 ;
    END
  END sram1_dout0[31]
  PIN sram1_dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 415.520 350.000 416.120 ;
    END
  END sram1_dout0[32]
  PIN sram1_dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 418.240 350.000 418.840 ;
    END
  END sram1_dout0[33]
  PIN sram1_dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 420.960 350.000 421.560 ;
    END
  END sram1_dout0[34]
  PIN sram1_dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 423.680 350.000 424.280 ;
    END
  END sram1_dout0[35]
  PIN sram1_dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 426.400 350.000 427.000 ;
    END
  END sram1_dout0[36]
  PIN sram1_dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 429.120 350.000 429.720 ;
    END
  END sram1_dout0[37]
  PIN sram1_dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 431.160 350.000 431.760 ;
    END
  END sram1_dout0[38]
  PIN sram1_dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 433.880 350.000 434.480 ;
    END
  END sram1_dout0[39]
  PIN sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 338.680 350.000 339.280 ;
    END
  END sram1_dout0[3]
  PIN sram1_dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 436.600 350.000 437.200 ;
    END
  END sram1_dout0[40]
  PIN sram1_dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 439.320 350.000 439.920 ;
    END
  END sram1_dout0[41]
  PIN sram1_dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 442.040 350.000 442.640 ;
    END
  END sram1_dout0[42]
  PIN sram1_dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 444.760 350.000 445.360 ;
    END
  END sram1_dout0[43]
  PIN sram1_dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 447.480 350.000 448.080 ;
    END
  END sram1_dout0[44]
  PIN sram1_dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 450.200 350.000 450.800 ;
    END
  END sram1_dout0[45]
  PIN sram1_dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 452.920 350.000 453.520 ;
    END
  END sram1_dout0[46]
  PIN sram1_dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 454.960 350.000 455.560 ;
    END
  END sram1_dout0[47]
  PIN sram1_dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 457.680 350.000 458.280 ;
    END
  END sram1_dout0[48]
  PIN sram1_dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 460.400 350.000 461.000 ;
    END
  END sram1_dout0[49]
  PIN sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 341.400 350.000 342.000 ;
    END
  END sram1_dout0[4]
  PIN sram1_dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 463.120 350.000 463.720 ;
    END
  END sram1_dout0[50]
  PIN sram1_dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 465.840 350.000 466.440 ;
    END
  END sram1_dout0[51]
  PIN sram1_dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 468.560 350.000 469.160 ;
    END
  END sram1_dout0[52]
  PIN sram1_dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 471.280 350.000 471.880 ;
    END
  END sram1_dout0[53]
  PIN sram1_dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 474.000 350.000 474.600 ;
    END
  END sram1_dout0[54]
  PIN sram1_dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 476.720 350.000 477.320 ;
    END
  END sram1_dout0[55]
  PIN sram1_dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 478.760 350.000 479.360 ;
    END
  END sram1_dout0[56]
  PIN sram1_dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 481.480 350.000 482.080 ;
    END
  END sram1_dout0[57]
  PIN sram1_dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 484.200 350.000 484.800 ;
    END
  END sram1_dout0[58]
  PIN sram1_dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 486.920 350.000 487.520 ;
    END
  END sram1_dout0[59]
  PIN sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 344.120 350.000 344.720 ;
    END
  END sram1_dout0[5]
  PIN sram1_dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 489.640 350.000 490.240 ;
    END
  END sram1_dout0[60]
  PIN sram1_dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 492.360 350.000 492.960 ;
    END
  END sram1_dout0[61]
  PIN sram1_dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 495.080 350.000 495.680 ;
    END
  END sram1_dout0[62]
  PIN sram1_dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 497.800 350.000 498.400 ;
    END
  END sram1_dout0[63]
  PIN sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 346.840 350.000 347.440 ;
    END
  END sram1_dout0[6]
  PIN sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 349.560 350.000 350.160 ;
    END
  END sram1_dout0[7]
  PIN sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 352.280 350.000 352.880 ;
    END
  END sram1_dout0[8]
  PIN sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 355.000 350.000 355.600 ;
    END
  END sram1_dout0[9]
  PIN sram1_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 32.000 350.000 32.600 ;
    END
  END sram1_dout1[0]
  PIN sram1_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 58.520 350.000 59.120 ;
    END
  END sram1_dout1[10]
  PIN sram1_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 61.240 350.000 61.840 ;
    END
  END sram1_dout1[11]
  PIN sram1_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 63.960 350.000 64.560 ;
    END
  END sram1_dout1[12]
  PIN sram1_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 66.680 350.000 67.280 ;
    END
  END sram1_dout1[13]
  PIN sram1_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 69.400 350.000 70.000 ;
    END
  END sram1_dout1[14]
  PIN sram1_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 72.120 350.000 72.720 ;
    END
  END sram1_dout1[15]
  PIN sram1_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 74.160 350.000 74.760 ;
    END
  END sram1_dout1[16]
  PIN sram1_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 76.880 350.000 77.480 ;
    END
  END sram1_dout1[17]
  PIN sram1_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 79.600 350.000 80.200 ;
    END
  END sram1_dout1[18]
  PIN sram1_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 82.320 350.000 82.920 ;
    END
  END sram1_dout1[19]
  PIN sram1_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 34.720 350.000 35.320 ;
    END
  END sram1_dout1[1]
  PIN sram1_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 85.040 350.000 85.640 ;
    END
  END sram1_dout1[20]
  PIN sram1_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 87.760 350.000 88.360 ;
    END
  END sram1_dout1[21]
  PIN sram1_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 90.480 350.000 91.080 ;
    END
  END sram1_dout1[22]
  PIN sram1_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 93.200 350.000 93.800 ;
    END
  END sram1_dout1[23]
  PIN sram1_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 95.920 350.000 96.520 ;
    END
  END sram1_dout1[24]
  PIN sram1_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 97.960 350.000 98.560 ;
    END
  END sram1_dout1[25]
  PIN sram1_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 100.680 350.000 101.280 ;
    END
  END sram1_dout1[26]
  PIN sram1_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 103.400 350.000 104.000 ;
    END
  END sram1_dout1[27]
  PIN sram1_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 106.120 350.000 106.720 ;
    END
  END sram1_dout1[28]
  PIN sram1_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 108.840 350.000 109.440 ;
    END
  END sram1_dout1[29]
  PIN sram1_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 37.440 350.000 38.040 ;
    END
  END sram1_dout1[2]
  PIN sram1_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 111.560 350.000 112.160 ;
    END
  END sram1_dout1[30]
  PIN sram1_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 114.280 350.000 114.880 ;
    END
  END sram1_dout1[31]
  PIN sram1_dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 117.000 350.000 117.600 ;
    END
  END sram1_dout1[32]
  PIN sram1_dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 119.720 350.000 120.320 ;
    END
  END sram1_dout1[33]
  PIN sram1_dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 121.760 350.000 122.360 ;
    END
  END sram1_dout1[34]
  PIN sram1_dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 124.480 350.000 125.080 ;
    END
  END sram1_dout1[35]
  PIN sram1_dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 127.200 350.000 127.800 ;
    END
  END sram1_dout1[36]
  PIN sram1_dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 129.920 350.000 130.520 ;
    END
  END sram1_dout1[37]
  PIN sram1_dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 132.640 350.000 133.240 ;
    END
  END sram1_dout1[38]
  PIN sram1_dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 135.360 350.000 135.960 ;
    END
  END sram1_dout1[39]
  PIN sram1_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 40.160 350.000 40.760 ;
    END
  END sram1_dout1[3]
  PIN sram1_dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 138.080 350.000 138.680 ;
    END
  END sram1_dout1[40]
  PIN sram1_dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 140.800 350.000 141.400 ;
    END
  END sram1_dout1[41]
  PIN sram1_dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 143.520 350.000 144.120 ;
    END
  END sram1_dout1[42]
  PIN sram1_dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 145.560 350.000 146.160 ;
    END
  END sram1_dout1[43]
  PIN sram1_dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 148.280 350.000 148.880 ;
    END
  END sram1_dout1[44]
  PIN sram1_dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 151.000 350.000 151.600 ;
    END
  END sram1_dout1[45]
  PIN sram1_dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 153.720 350.000 154.320 ;
    END
  END sram1_dout1[46]
  PIN sram1_dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 156.440 350.000 157.040 ;
    END
  END sram1_dout1[47]
  PIN sram1_dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 159.160 350.000 159.760 ;
    END
  END sram1_dout1[48]
  PIN sram1_dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 161.880 350.000 162.480 ;
    END
  END sram1_dout1[49]
  PIN sram1_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 42.880 350.000 43.480 ;
    END
  END sram1_dout1[4]
  PIN sram1_dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 164.600 350.000 165.200 ;
    END
  END sram1_dout1[50]
  PIN sram1_dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 167.320 350.000 167.920 ;
    END
  END sram1_dout1[51]
  PIN sram1_dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 169.360 350.000 169.960 ;
    END
  END sram1_dout1[52]
  PIN sram1_dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 172.080 350.000 172.680 ;
    END
  END sram1_dout1[53]
  PIN sram1_dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 174.800 350.000 175.400 ;
    END
  END sram1_dout1[54]
  PIN sram1_dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 177.520 350.000 178.120 ;
    END
  END sram1_dout1[55]
  PIN sram1_dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 180.240 350.000 180.840 ;
    END
  END sram1_dout1[56]
  PIN sram1_dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 182.960 350.000 183.560 ;
    END
  END sram1_dout1[57]
  PIN sram1_dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 185.680 350.000 186.280 ;
    END
  END sram1_dout1[58]
  PIN sram1_dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 188.400 350.000 189.000 ;
    END
  END sram1_dout1[59]
  PIN sram1_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 45.600 350.000 46.200 ;
    END
  END sram1_dout1[5]
  PIN sram1_dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 191.120 350.000 191.720 ;
    END
  END sram1_dout1[60]
  PIN sram1_dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 193.160 350.000 193.760 ;
    END
  END sram1_dout1[61]
  PIN sram1_dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 195.880 350.000 196.480 ;
    END
  END sram1_dout1[62]
  PIN sram1_dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 198.600 350.000 199.200 ;
    END
  END sram1_dout1[63]
  PIN sram1_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 48.320 350.000 48.920 ;
    END
  END sram1_dout1[6]
  PIN sram1_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 50.360 350.000 50.960 ;
    END
  END sram1_dout1[7]
  PIN sram1_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 53.080 350.000 53.680 ;
    END
  END sram1_dout1[8]
  PIN sram1_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 55.800 350.000 56.400 ;
    END
  END sram1_dout1[9]
  PIN sram1_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 209.480 350.000 210.080 ;
    END
  END sram1_web0
  PIN sram1_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 212.200 350.000 212.800 ;
    END
  END sram1_wmask0[0]
  PIN sram1_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 214.920 350.000 215.520 ;
    END
  END sram1_wmask0[1]
  PIN sram1_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 216.960 350.000 217.560 ;
    END
  END sram1_wmask0[2]
  PIN sram1_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 219.680 350.000 220.280 ;
    END
  END sram1_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END vga_vsync
  PIN video_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END video_irq[0]
  PIN video_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 496.000 175.170 500.000 ;
    END
  END video_irq[1]
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 4.000 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 486.965 ;
      LAYER met1 ;
        RECT 1.450 7.860 348.610 487.120 ;
      LAYER met2 ;
        RECT 1.480 495.720 174.610 498.285 ;
        RECT 175.450 495.720 348.580 498.285 ;
        RECT 1.480 4.280 348.580 495.720 ;
        RECT 2.030 0.270 3.950 4.280 ;
        RECT 4.790 0.270 7.170 4.280 ;
        RECT 8.010 0.270 10.390 4.280 ;
        RECT 11.230 0.270 13.610 4.280 ;
        RECT 14.450 0.270 16.830 4.280 ;
        RECT 17.670 0.270 20.050 4.280 ;
        RECT 20.890 0.270 23.270 4.280 ;
        RECT 24.110 0.270 26.490 4.280 ;
        RECT 27.330 0.270 29.710 4.280 ;
        RECT 30.550 0.270 32.930 4.280 ;
        RECT 33.770 0.270 36.150 4.280 ;
        RECT 36.990 0.270 39.370 4.280 ;
        RECT 40.210 0.270 42.590 4.280 ;
        RECT 43.430 0.270 45.810 4.280 ;
        RECT 46.650 0.270 49.030 4.280 ;
        RECT 49.870 0.270 52.250 4.280 ;
        RECT 53.090 0.270 55.470 4.280 ;
        RECT 56.310 0.270 58.690 4.280 ;
        RECT 59.530 0.270 61.910 4.280 ;
        RECT 62.750 0.270 65.130 4.280 ;
        RECT 65.970 0.270 68.350 4.280 ;
        RECT 69.190 0.270 71.570 4.280 ;
        RECT 72.410 0.270 74.790 4.280 ;
        RECT 75.630 0.270 78.010 4.280 ;
        RECT 78.850 0.270 81.230 4.280 ;
        RECT 82.070 0.270 84.450 4.280 ;
        RECT 85.290 0.270 87.670 4.280 ;
        RECT 88.510 0.270 90.890 4.280 ;
        RECT 91.730 0.270 94.110 4.280 ;
        RECT 94.950 0.270 97.330 4.280 ;
        RECT 98.170 0.270 100.550 4.280 ;
        RECT 101.390 0.270 103.770 4.280 ;
        RECT 104.610 0.270 106.990 4.280 ;
        RECT 107.830 0.270 110.210 4.280 ;
        RECT 111.050 0.270 113.430 4.280 ;
        RECT 114.270 0.270 116.650 4.280 ;
        RECT 117.490 0.270 119.870 4.280 ;
        RECT 120.710 0.270 123.090 4.280 ;
        RECT 123.930 0.270 126.310 4.280 ;
        RECT 127.150 0.270 129.530 4.280 ;
        RECT 130.370 0.270 132.750 4.280 ;
        RECT 133.590 0.270 135.970 4.280 ;
        RECT 136.810 0.270 139.190 4.280 ;
        RECT 140.030 0.270 142.410 4.280 ;
        RECT 143.250 0.270 145.630 4.280 ;
        RECT 146.470 0.270 148.850 4.280 ;
        RECT 149.690 0.270 152.070 4.280 ;
        RECT 152.910 0.270 155.290 4.280 ;
        RECT 156.130 0.270 158.510 4.280 ;
        RECT 159.350 0.270 161.730 4.280 ;
        RECT 162.570 0.270 164.950 4.280 ;
        RECT 165.790 0.270 168.170 4.280 ;
        RECT 169.010 0.270 171.390 4.280 ;
        RECT 172.230 0.270 174.610 4.280 ;
        RECT 175.450 0.270 177.370 4.280 ;
        RECT 178.210 0.270 180.590 4.280 ;
        RECT 181.430 0.270 183.810 4.280 ;
        RECT 184.650 0.270 187.030 4.280 ;
        RECT 187.870 0.270 190.250 4.280 ;
        RECT 191.090 0.270 193.470 4.280 ;
        RECT 194.310 0.270 196.690 4.280 ;
        RECT 197.530 0.270 199.910 4.280 ;
        RECT 200.750 0.270 203.130 4.280 ;
        RECT 203.970 0.270 206.350 4.280 ;
        RECT 207.190 0.270 209.570 4.280 ;
        RECT 210.410 0.270 212.790 4.280 ;
        RECT 213.630 0.270 216.010 4.280 ;
        RECT 216.850 0.270 219.230 4.280 ;
        RECT 220.070 0.270 222.450 4.280 ;
        RECT 223.290 0.270 225.670 4.280 ;
        RECT 226.510 0.270 228.890 4.280 ;
        RECT 229.730 0.270 232.110 4.280 ;
        RECT 232.950 0.270 235.330 4.280 ;
        RECT 236.170 0.270 238.550 4.280 ;
        RECT 239.390 0.270 241.770 4.280 ;
        RECT 242.610 0.270 244.990 4.280 ;
        RECT 245.830 0.270 248.210 4.280 ;
        RECT 249.050 0.270 251.430 4.280 ;
        RECT 252.270 0.270 254.650 4.280 ;
        RECT 255.490 0.270 257.870 4.280 ;
        RECT 258.710 0.270 261.090 4.280 ;
        RECT 261.930 0.270 264.310 4.280 ;
        RECT 265.150 0.270 267.530 4.280 ;
        RECT 268.370 0.270 270.750 4.280 ;
        RECT 271.590 0.270 273.970 4.280 ;
        RECT 274.810 0.270 277.190 4.280 ;
        RECT 278.030 0.270 280.410 4.280 ;
        RECT 281.250 0.270 283.630 4.280 ;
        RECT 284.470 0.270 286.850 4.280 ;
        RECT 287.690 0.270 290.070 4.280 ;
        RECT 290.910 0.270 293.290 4.280 ;
        RECT 294.130 0.270 296.510 4.280 ;
        RECT 297.350 0.270 299.730 4.280 ;
        RECT 300.570 0.270 302.950 4.280 ;
        RECT 303.790 0.270 306.170 4.280 ;
        RECT 307.010 0.270 309.390 4.280 ;
        RECT 310.230 0.270 312.610 4.280 ;
        RECT 313.450 0.270 315.830 4.280 ;
        RECT 316.670 0.270 319.050 4.280 ;
        RECT 319.890 0.270 322.270 4.280 ;
        RECT 323.110 0.270 325.490 4.280 ;
        RECT 326.330 0.270 328.710 4.280 ;
        RECT 329.550 0.270 331.930 4.280 ;
        RECT 332.770 0.270 335.150 4.280 ;
        RECT 335.990 0.270 338.370 4.280 ;
        RECT 339.210 0.270 341.590 4.280 ;
        RECT 342.430 0.270 344.810 4.280 ;
        RECT 345.650 0.270 348.030 4.280 ;
      LAYER met3 ;
        RECT 4.400 497.400 345.600 498.265 ;
        RECT 4.000 496.080 346.000 497.400 ;
        RECT 4.400 494.680 345.600 496.080 ;
        RECT 4.000 493.360 346.000 494.680 ;
        RECT 4.400 491.960 345.600 493.360 ;
        RECT 4.000 490.640 346.000 491.960 ;
        RECT 4.400 489.240 345.600 490.640 ;
        RECT 4.000 487.920 346.000 489.240 ;
        RECT 4.400 486.520 345.600 487.920 ;
        RECT 4.000 485.200 346.000 486.520 ;
        RECT 4.400 483.800 345.600 485.200 ;
        RECT 4.000 482.480 346.000 483.800 ;
        RECT 4.400 481.080 345.600 482.480 ;
        RECT 4.000 479.760 346.000 481.080 ;
        RECT 4.400 478.360 345.600 479.760 ;
        RECT 4.000 477.720 346.000 478.360 ;
        RECT 4.400 476.320 345.600 477.720 ;
        RECT 4.000 475.000 346.000 476.320 ;
        RECT 4.400 473.600 345.600 475.000 ;
        RECT 4.000 472.280 346.000 473.600 ;
        RECT 4.400 470.880 345.600 472.280 ;
        RECT 4.000 469.560 346.000 470.880 ;
        RECT 4.400 468.160 345.600 469.560 ;
        RECT 4.000 466.840 346.000 468.160 ;
        RECT 4.400 465.440 345.600 466.840 ;
        RECT 4.000 464.120 346.000 465.440 ;
        RECT 4.400 462.720 345.600 464.120 ;
        RECT 4.000 461.400 346.000 462.720 ;
        RECT 4.400 460.000 345.600 461.400 ;
        RECT 4.000 458.680 346.000 460.000 ;
        RECT 4.400 457.280 345.600 458.680 ;
        RECT 4.000 455.960 346.000 457.280 ;
        RECT 4.400 454.560 345.600 455.960 ;
        RECT 4.000 453.920 346.000 454.560 ;
        RECT 4.400 452.520 345.600 453.920 ;
        RECT 4.000 451.200 346.000 452.520 ;
        RECT 4.400 449.800 345.600 451.200 ;
        RECT 4.000 448.480 346.000 449.800 ;
        RECT 4.400 447.080 345.600 448.480 ;
        RECT 4.000 445.760 346.000 447.080 ;
        RECT 4.400 444.360 345.600 445.760 ;
        RECT 4.000 443.040 346.000 444.360 ;
        RECT 4.400 441.640 345.600 443.040 ;
        RECT 4.000 440.320 346.000 441.640 ;
        RECT 4.400 438.920 345.600 440.320 ;
        RECT 4.000 437.600 346.000 438.920 ;
        RECT 4.400 436.200 345.600 437.600 ;
        RECT 4.000 434.880 346.000 436.200 ;
        RECT 4.400 433.480 345.600 434.880 ;
        RECT 4.000 432.160 346.000 433.480 ;
        RECT 4.400 430.760 345.600 432.160 ;
        RECT 4.000 430.120 346.000 430.760 ;
        RECT 4.400 428.720 345.600 430.120 ;
        RECT 4.000 427.400 346.000 428.720 ;
        RECT 4.400 426.000 345.600 427.400 ;
        RECT 4.000 424.680 346.000 426.000 ;
        RECT 4.400 423.280 345.600 424.680 ;
        RECT 4.000 421.960 346.000 423.280 ;
        RECT 4.400 420.560 345.600 421.960 ;
        RECT 4.000 419.240 346.000 420.560 ;
        RECT 4.400 417.840 345.600 419.240 ;
        RECT 4.000 416.520 346.000 417.840 ;
        RECT 4.400 415.120 345.600 416.520 ;
        RECT 4.000 413.800 346.000 415.120 ;
        RECT 4.400 412.400 345.600 413.800 ;
        RECT 4.000 411.080 346.000 412.400 ;
        RECT 4.400 409.680 345.600 411.080 ;
        RECT 4.000 408.360 346.000 409.680 ;
        RECT 4.400 406.960 345.600 408.360 ;
        RECT 4.000 406.320 346.000 406.960 ;
        RECT 4.400 404.920 345.600 406.320 ;
        RECT 4.000 403.600 346.000 404.920 ;
        RECT 4.400 402.200 345.600 403.600 ;
        RECT 4.000 400.880 346.000 402.200 ;
        RECT 4.400 399.480 345.600 400.880 ;
        RECT 4.000 398.160 346.000 399.480 ;
        RECT 4.400 396.760 345.600 398.160 ;
        RECT 4.000 395.440 346.000 396.760 ;
        RECT 4.400 394.040 345.600 395.440 ;
        RECT 4.000 392.720 346.000 394.040 ;
        RECT 4.400 391.320 345.600 392.720 ;
        RECT 4.000 390.000 346.000 391.320 ;
        RECT 4.400 388.600 345.600 390.000 ;
        RECT 4.000 387.280 346.000 388.600 ;
        RECT 4.400 385.880 345.600 387.280 ;
        RECT 4.000 384.560 346.000 385.880 ;
        RECT 4.400 383.160 345.600 384.560 ;
        RECT 4.000 382.520 346.000 383.160 ;
        RECT 4.400 381.120 345.600 382.520 ;
        RECT 4.000 379.800 346.000 381.120 ;
        RECT 4.400 378.400 345.600 379.800 ;
        RECT 4.000 377.080 346.000 378.400 ;
        RECT 4.400 375.680 345.600 377.080 ;
        RECT 4.000 374.360 346.000 375.680 ;
        RECT 4.400 372.960 345.600 374.360 ;
        RECT 4.000 371.640 346.000 372.960 ;
        RECT 4.400 370.240 345.600 371.640 ;
        RECT 4.000 368.920 346.000 370.240 ;
        RECT 4.400 367.520 345.600 368.920 ;
        RECT 4.000 366.200 346.000 367.520 ;
        RECT 4.400 364.800 345.600 366.200 ;
        RECT 4.000 363.480 346.000 364.800 ;
        RECT 4.400 362.080 345.600 363.480 ;
        RECT 4.000 360.760 346.000 362.080 ;
        RECT 4.400 359.360 345.600 360.760 ;
        RECT 4.000 358.720 346.000 359.360 ;
        RECT 4.400 357.320 345.600 358.720 ;
        RECT 4.000 356.000 346.000 357.320 ;
        RECT 4.400 354.600 345.600 356.000 ;
        RECT 4.000 353.280 346.000 354.600 ;
        RECT 4.400 351.880 345.600 353.280 ;
        RECT 4.000 350.560 346.000 351.880 ;
        RECT 4.400 349.160 345.600 350.560 ;
        RECT 4.000 347.840 346.000 349.160 ;
        RECT 4.400 346.440 345.600 347.840 ;
        RECT 4.000 345.120 346.000 346.440 ;
        RECT 4.400 343.720 345.600 345.120 ;
        RECT 4.000 342.400 346.000 343.720 ;
        RECT 4.400 341.000 345.600 342.400 ;
        RECT 4.000 339.680 346.000 341.000 ;
        RECT 4.400 338.280 345.600 339.680 ;
        RECT 4.000 336.960 346.000 338.280 ;
        RECT 4.400 335.560 345.600 336.960 ;
        RECT 4.000 334.920 346.000 335.560 ;
        RECT 4.400 333.520 345.600 334.920 ;
        RECT 4.000 332.200 346.000 333.520 ;
        RECT 4.400 330.800 345.600 332.200 ;
        RECT 4.000 329.480 346.000 330.800 ;
        RECT 4.400 328.080 345.600 329.480 ;
        RECT 4.000 326.760 346.000 328.080 ;
        RECT 4.400 325.360 345.600 326.760 ;
        RECT 4.000 324.040 346.000 325.360 ;
        RECT 4.400 322.640 345.600 324.040 ;
        RECT 4.000 321.320 346.000 322.640 ;
        RECT 4.400 319.920 345.600 321.320 ;
        RECT 4.000 318.600 346.000 319.920 ;
        RECT 4.400 317.200 345.600 318.600 ;
        RECT 4.000 315.880 346.000 317.200 ;
        RECT 4.400 314.480 345.600 315.880 ;
        RECT 4.000 313.160 346.000 314.480 ;
        RECT 4.400 311.760 345.600 313.160 ;
        RECT 4.000 311.120 346.000 311.760 ;
        RECT 4.400 309.720 345.600 311.120 ;
        RECT 4.000 308.400 346.000 309.720 ;
        RECT 4.400 307.000 345.600 308.400 ;
        RECT 4.000 305.680 346.000 307.000 ;
        RECT 4.400 304.280 345.600 305.680 ;
        RECT 4.000 302.960 346.000 304.280 ;
        RECT 4.400 301.560 345.600 302.960 ;
        RECT 4.000 300.240 346.000 301.560 ;
        RECT 4.400 298.840 345.600 300.240 ;
        RECT 4.000 297.520 346.000 298.840 ;
        RECT 4.400 296.120 345.600 297.520 ;
        RECT 4.000 294.800 346.000 296.120 ;
        RECT 4.400 293.400 345.600 294.800 ;
        RECT 4.000 292.080 346.000 293.400 ;
        RECT 4.400 290.680 345.600 292.080 ;
        RECT 4.000 289.360 346.000 290.680 ;
        RECT 4.400 287.960 345.600 289.360 ;
        RECT 4.000 287.320 346.000 287.960 ;
        RECT 4.400 285.920 345.600 287.320 ;
        RECT 4.000 284.600 346.000 285.920 ;
        RECT 4.400 283.200 345.600 284.600 ;
        RECT 4.000 281.880 346.000 283.200 ;
        RECT 4.400 280.480 345.600 281.880 ;
        RECT 4.000 279.160 346.000 280.480 ;
        RECT 4.400 277.760 345.600 279.160 ;
        RECT 4.000 276.440 346.000 277.760 ;
        RECT 4.400 275.040 345.600 276.440 ;
        RECT 4.000 273.720 346.000 275.040 ;
        RECT 4.400 272.320 345.600 273.720 ;
        RECT 4.000 271.000 346.000 272.320 ;
        RECT 4.400 269.600 345.600 271.000 ;
        RECT 4.000 268.280 346.000 269.600 ;
        RECT 4.400 266.880 345.600 268.280 ;
        RECT 4.000 265.560 346.000 266.880 ;
        RECT 4.400 264.160 345.600 265.560 ;
        RECT 4.000 263.520 346.000 264.160 ;
        RECT 4.400 262.120 345.600 263.520 ;
        RECT 4.000 260.800 346.000 262.120 ;
        RECT 4.400 259.400 345.600 260.800 ;
        RECT 4.000 258.080 346.000 259.400 ;
        RECT 4.400 256.680 345.600 258.080 ;
        RECT 4.000 255.360 346.000 256.680 ;
        RECT 4.400 253.960 345.600 255.360 ;
        RECT 4.000 252.640 346.000 253.960 ;
        RECT 4.400 251.240 345.600 252.640 ;
        RECT 4.000 249.920 346.000 251.240 ;
        RECT 4.400 248.520 345.600 249.920 ;
        RECT 4.000 247.200 346.000 248.520 ;
        RECT 4.400 245.800 345.600 247.200 ;
        RECT 4.000 244.480 346.000 245.800 ;
        RECT 4.400 243.080 345.600 244.480 ;
        RECT 4.000 241.760 346.000 243.080 ;
        RECT 4.400 240.360 345.600 241.760 ;
        RECT 4.000 239.720 346.000 240.360 ;
        RECT 4.400 238.320 345.600 239.720 ;
        RECT 4.000 237.000 346.000 238.320 ;
        RECT 4.400 235.600 345.600 237.000 ;
        RECT 4.000 234.280 346.000 235.600 ;
        RECT 4.400 232.880 345.600 234.280 ;
        RECT 4.000 231.560 346.000 232.880 ;
        RECT 4.400 230.160 345.600 231.560 ;
        RECT 4.000 228.840 346.000 230.160 ;
        RECT 4.400 227.440 345.600 228.840 ;
        RECT 4.000 226.120 346.000 227.440 ;
        RECT 4.400 224.720 345.600 226.120 ;
        RECT 4.000 223.400 346.000 224.720 ;
        RECT 4.400 222.000 345.600 223.400 ;
        RECT 4.000 220.680 346.000 222.000 ;
        RECT 4.400 219.280 345.600 220.680 ;
        RECT 4.000 217.960 346.000 219.280 ;
        RECT 4.400 216.560 345.600 217.960 ;
        RECT 4.000 215.920 346.000 216.560 ;
        RECT 4.400 214.520 345.600 215.920 ;
        RECT 4.000 213.200 346.000 214.520 ;
        RECT 4.400 211.800 345.600 213.200 ;
        RECT 4.000 210.480 346.000 211.800 ;
        RECT 4.400 209.080 345.600 210.480 ;
        RECT 4.000 207.760 346.000 209.080 ;
        RECT 4.400 206.360 345.600 207.760 ;
        RECT 4.000 205.040 346.000 206.360 ;
        RECT 4.400 203.640 345.600 205.040 ;
        RECT 4.000 202.320 346.000 203.640 ;
        RECT 4.400 200.920 345.600 202.320 ;
        RECT 4.000 199.600 346.000 200.920 ;
        RECT 4.400 198.200 345.600 199.600 ;
        RECT 4.000 196.880 346.000 198.200 ;
        RECT 4.400 195.480 345.600 196.880 ;
        RECT 4.000 194.160 346.000 195.480 ;
        RECT 4.400 192.760 345.600 194.160 ;
        RECT 4.000 192.120 346.000 192.760 ;
        RECT 4.400 190.720 345.600 192.120 ;
        RECT 4.000 189.400 346.000 190.720 ;
        RECT 4.400 188.000 345.600 189.400 ;
        RECT 4.000 186.680 346.000 188.000 ;
        RECT 4.400 185.280 345.600 186.680 ;
        RECT 4.000 183.960 346.000 185.280 ;
        RECT 4.400 182.560 345.600 183.960 ;
        RECT 4.000 181.240 346.000 182.560 ;
        RECT 4.400 179.840 345.600 181.240 ;
        RECT 4.000 178.520 346.000 179.840 ;
        RECT 4.400 177.120 345.600 178.520 ;
        RECT 4.000 175.800 346.000 177.120 ;
        RECT 4.400 174.400 345.600 175.800 ;
        RECT 4.000 173.080 346.000 174.400 ;
        RECT 4.400 171.680 345.600 173.080 ;
        RECT 4.000 170.360 346.000 171.680 ;
        RECT 4.400 168.960 345.600 170.360 ;
        RECT 4.000 168.320 346.000 168.960 ;
        RECT 4.400 166.920 345.600 168.320 ;
        RECT 4.000 165.600 346.000 166.920 ;
        RECT 4.400 164.200 345.600 165.600 ;
        RECT 4.000 162.880 346.000 164.200 ;
        RECT 4.400 161.480 345.600 162.880 ;
        RECT 4.000 160.160 346.000 161.480 ;
        RECT 4.400 158.760 345.600 160.160 ;
        RECT 4.000 157.440 346.000 158.760 ;
        RECT 4.400 156.040 345.600 157.440 ;
        RECT 4.000 154.720 346.000 156.040 ;
        RECT 4.400 153.320 345.600 154.720 ;
        RECT 4.000 152.000 346.000 153.320 ;
        RECT 4.400 150.600 345.600 152.000 ;
        RECT 4.000 149.280 346.000 150.600 ;
        RECT 4.400 147.880 345.600 149.280 ;
        RECT 4.000 146.560 346.000 147.880 ;
        RECT 4.400 145.160 345.600 146.560 ;
        RECT 4.000 144.520 346.000 145.160 ;
        RECT 4.400 143.120 345.600 144.520 ;
        RECT 4.000 141.800 346.000 143.120 ;
        RECT 4.400 140.400 345.600 141.800 ;
        RECT 4.000 139.080 346.000 140.400 ;
        RECT 4.400 137.680 345.600 139.080 ;
        RECT 4.000 136.360 346.000 137.680 ;
        RECT 4.400 134.960 345.600 136.360 ;
        RECT 4.000 133.640 346.000 134.960 ;
        RECT 4.400 132.240 345.600 133.640 ;
        RECT 4.000 130.920 346.000 132.240 ;
        RECT 4.400 129.520 345.600 130.920 ;
        RECT 4.000 128.200 346.000 129.520 ;
        RECT 4.400 126.800 345.600 128.200 ;
        RECT 4.000 125.480 346.000 126.800 ;
        RECT 4.400 124.080 345.600 125.480 ;
        RECT 4.000 122.760 346.000 124.080 ;
        RECT 4.400 121.360 345.600 122.760 ;
        RECT 4.000 120.720 346.000 121.360 ;
        RECT 4.400 119.320 345.600 120.720 ;
        RECT 4.000 118.000 346.000 119.320 ;
        RECT 4.400 116.600 345.600 118.000 ;
        RECT 4.000 115.280 346.000 116.600 ;
        RECT 4.400 113.880 345.600 115.280 ;
        RECT 4.000 112.560 346.000 113.880 ;
        RECT 4.400 111.160 345.600 112.560 ;
        RECT 4.000 109.840 346.000 111.160 ;
        RECT 4.400 108.440 345.600 109.840 ;
        RECT 4.000 107.120 346.000 108.440 ;
        RECT 4.400 105.720 345.600 107.120 ;
        RECT 4.000 104.400 346.000 105.720 ;
        RECT 4.400 103.000 345.600 104.400 ;
        RECT 4.000 101.680 346.000 103.000 ;
        RECT 4.400 100.280 345.600 101.680 ;
        RECT 4.000 98.960 346.000 100.280 ;
        RECT 4.400 97.560 345.600 98.960 ;
        RECT 4.000 96.920 346.000 97.560 ;
        RECT 4.400 95.520 345.600 96.920 ;
        RECT 4.000 94.200 346.000 95.520 ;
        RECT 4.400 92.800 345.600 94.200 ;
        RECT 4.000 91.480 346.000 92.800 ;
        RECT 4.400 90.080 345.600 91.480 ;
        RECT 4.000 88.760 346.000 90.080 ;
        RECT 4.400 87.360 345.600 88.760 ;
        RECT 4.000 86.040 346.000 87.360 ;
        RECT 4.400 84.640 345.600 86.040 ;
        RECT 4.000 83.320 346.000 84.640 ;
        RECT 4.400 81.920 345.600 83.320 ;
        RECT 4.000 80.600 346.000 81.920 ;
        RECT 4.400 79.200 345.600 80.600 ;
        RECT 4.000 77.880 346.000 79.200 ;
        RECT 4.400 76.480 345.600 77.880 ;
        RECT 4.000 75.160 346.000 76.480 ;
        RECT 4.400 73.760 345.600 75.160 ;
        RECT 4.000 73.120 346.000 73.760 ;
        RECT 4.400 71.720 345.600 73.120 ;
        RECT 4.000 70.400 346.000 71.720 ;
        RECT 4.400 69.000 345.600 70.400 ;
        RECT 4.000 67.680 346.000 69.000 ;
        RECT 4.400 66.280 345.600 67.680 ;
        RECT 4.000 64.960 346.000 66.280 ;
        RECT 4.400 63.560 345.600 64.960 ;
        RECT 4.000 62.240 346.000 63.560 ;
        RECT 4.400 60.840 345.600 62.240 ;
        RECT 4.000 59.520 346.000 60.840 ;
        RECT 4.400 58.120 345.600 59.520 ;
        RECT 4.000 56.800 346.000 58.120 ;
        RECT 4.400 55.400 345.600 56.800 ;
        RECT 4.000 54.080 346.000 55.400 ;
        RECT 4.400 52.680 345.600 54.080 ;
        RECT 4.000 51.360 346.000 52.680 ;
        RECT 4.400 49.960 345.600 51.360 ;
        RECT 4.000 49.320 346.000 49.960 ;
        RECT 4.400 47.920 345.600 49.320 ;
        RECT 4.000 46.600 346.000 47.920 ;
        RECT 4.400 45.200 345.600 46.600 ;
        RECT 4.000 43.880 346.000 45.200 ;
        RECT 4.400 42.480 345.600 43.880 ;
        RECT 4.000 41.160 346.000 42.480 ;
        RECT 4.400 39.760 345.600 41.160 ;
        RECT 4.000 38.440 346.000 39.760 ;
        RECT 4.400 37.040 345.600 38.440 ;
        RECT 4.000 35.720 346.000 37.040 ;
        RECT 4.400 34.320 345.600 35.720 ;
        RECT 4.000 33.000 346.000 34.320 ;
        RECT 4.400 31.600 345.600 33.000 ;
        RECT 4.000 30.280 346.000 31.600 ;
        RECT 4.400 28.880 345.600 30.280 ;
        RECT 4.000 27.560 346.000 28.880 ;
        RECT 4.400 26.160 345.600 27.560 ;
        RECT 4.000 25.520 346.000 26.160 ;
        RECT 4.400 24.120 345.600 25.520 ;
        RECT 4.000 22.800 346.000 24.120 ;
        RECT 4.400 21.400 345.600 22.800 ;
        RECT 4.000 20.080 346.000 21.400 ;
        RECT 4.400 18.680 345.600 20.080 ;
        RECT 4.000 17.360 346.000 18.680 ;
        RECT 4.400 15.960 345.600 17.360 ;
        RECT 4.000 14.640 346.000 15.960 ;
        RECT 4.400 13.240 345.600 14.640 ;
        RECT 4.000 11.920 346.000 13.240 ;
        RECT 4.400 10.520 345.600 11.920 ;
        RECT 4.000 9.200 346.000 10.520 ;
        RECT 4.400 7.800 345.600 9.200 ;
        RECT 4.000 6.480 346.000 7.800 ;
        RECT 4.400 5.080 345.600 6.480 ;
        RECT 4.000 3.760 346.000 5.080 ;
        RECT 4.400 2.360 345.600 3.760 ;
        RECT 4.000 1.720 346.000 2.360 ;
        RECT 4.400 0.855 345.600 1.720 ;
      LAYER met4 ;
        RECT 7.655 132.095 20.640 468.345 ;
        RECT 23.040 132.095 97.440 468.345 ;
        RECT 99.840 132.095 174.240 468.345 ;
        RECT 176.640 132.095 251.040 468.345 ;
        RECT 253.440 132.095 327.840 468.345 ;
        RECT 330.240 132.095 335.505 468.345 ;
  END
END Video
END LIBRARY

