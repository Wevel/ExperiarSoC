VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Peripherals
  CLASS BLOCK ;
  FOREIGN Peripherals ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 750.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 746.000 2.670 750.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 746.000 147.110 750.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 746.000 161.830 750.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 746.000 176.090 750.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 746.000 190.810 750.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 746.000 205.070 750.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 746.000 219.790 750.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 746.000 234.050 750.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 746.000 248.770 750.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 746.000 263.030 750.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 746.000 277.750 750.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 746.000 16.930 750.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 746.000 292.010 750.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 746.000 306.270 750.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 746.000 320.990 750.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 746.000 335.250 750.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 746.000 349.970 750.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 746.000 364.230 750.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 746.000 378.950 750.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 746.000 393.210 750.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 746.000 407.930 750.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 746.000 422.190 750.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 746.000 31.190 750.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 746.000 436.910 750.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 746.000 451.170 750.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 746.000 465.890 750.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 746.000 480.150 750.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 746.000 494.870 750.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 746.000 509.130 750.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 746.000 523.850 750.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 746.000 538.110 750.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 746.000 45.910 750.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 746.000 60.170 750.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 746.000 74.890 750.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 746.000 89.150 750.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 746.000 103.870 750.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 746.000 118.130 750.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 746.000 132.850 750.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 746.000 7.270 750.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 746.000 152.170 750.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 746.000 166.430 750.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 746.000 181.150 750.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 746.000 195.410 750.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 746.000 210.130 750.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 746.000 224.390 750.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 746.000 239.110 750.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 746.000 253.370 750.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 746.000 268.090 750.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 746.000 282.350 750.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 746.000 21.530 750.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 746.000 296.610 750.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 746.000 311.330 750.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 746.000 325.590 750.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 746.000 340.310 750.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 746.000 354.570 750.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 746.000 369.290 750.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 746.000 383.550 750.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 746.000 398.270 750.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 746.000 412.530 750.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 746.000 427.250 750.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 746.000 36.250 750.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 746.000 441.510 750.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 746.000 456.230 750.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 746.000 470.490 750.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 746.000 485.210 750.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 746.000 499.470 750.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 746.000 514.190 750.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 746.000 528.450 750.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 746.000 543.170 750.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 746.000 50.510 750.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 746.000 65.230 750.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 746.000 79.490 750.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 746.000 94.210 750.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 746.000 108.470 750.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 746.000 123.190 750.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 746.000 137.450 750.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 746.000 11.870 750.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 746.000 156.770 750.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 746.000 171.490 750.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 746.000 185.750 750.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 746.000 200.470 750.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 746.000 214.730 750.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 746.000 229.450 750.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 746.000 243.710 750.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 746.000 258.430 750.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 746.000 272.690 750.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 746.000 286.950 750.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 746.000 26.590 750.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 746.000 301.670 750.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 746.000 315.930 750.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 746.000 330.650 750.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 746.000 344.910 750.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 746.000 359.630 750.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 746.000 373.890 750.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 746.000 388.610 750.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 746.000 402.870 750.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 746.000 417.590 750.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 746.000 431.850 750.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 746.000 40.850 750.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 746.000 446.570 750.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 746.000 460.830 750.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 746.000 475.550 750.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 746.000 489.810 750.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 746.000 504.530 750.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 746.000 518.790 750.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 746.000 533.510 750.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 746.000 547.770 750.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 746.000 55.570 750.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 746.000 69.830 750.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 746.000 84.550 750.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 746.000 98.810 750.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 746.000 113.530 750.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 746.000 127.790 750.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 746.000 142.510 750.000 ;
    END
  END io_out[9]
  PIN la_blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 187.040 550.000 187.640 ;
    END
  END la_blink[0]
  PIN la_blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 561.720 550.000 562.320 ;
    END
  END la_blink[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 737.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 737.360 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.760 4.000 496.360 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.760 4.000 564.360 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.800 4.000 617.400 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.280 4.000 692.880 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.920 4.000 708.520 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.600 4.000 420.200 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.720 4.000 443.320 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.720 4.000 511.320 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.880 4.000 655.480 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 4.000 745.920 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END wb_data_o[9]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 544.180 737.205 ;
      LAYER met1 ;
        RECT 2.370 10.640 547.790 737.760 ;
      LAYER met2 ;
        RECT 2.950 745.720 6.710 746.370 ;
        RECT 7.550 745.720 11.310 746.370 ;
        RECT 12.150 745.720 16.370 746.370 ;
        RECT 17.210 745.720 20.970 746.370 ;
        RECT 21.810 745.720 26.030 746.370 ;
        RECT 26.870 745.720 30.630 746.370 ;
        RECT 31.470 745.720 35.690 746.370 ;
        RECT 36.530 745.720 40.290 746.370 ;
        RECT 41.130 745.720 45.350 746.370 ;
        RECT 46.190 745.720 49.950 746.370 ;
        RECT 50.790 745.720 55.010 746.370 ;
        RECT 55.850 745.720 59.610 746.370 ;
        RECT 60.450 745.720 64.670 746.370 ;
        RECT 65.510 745.720 69.270 746.370 ;
        RECT 70.110 745.720 74.330 746.370 ;
        RECT 75.170 745.720 78.930 746.370 ;
        RECT 79.770 745.720 83.990 746.370 ;
        RECT 84.830 745.720 88.590 746.370 ;
        RECT 89.430 745.720 93.650 746.370 ;
        RECT 94.490 745.720 98.250 746.370 ;
        RECT 99.090 745.720 103.310 746.370 ;
        RECT 104.150 745.720 107.910 746.370 ;
        RECT 108.750 745.720 112.970 746.370 ;
        RECT 113.810 745.720 117.570 746.370 ;
        RECT 118.410 745.720 122.630 746.370 ;
        RECT 123.470 745.720 127.230 746.370 ;
        RECT 128.070 745.720 132.290 746.370 ;
        RECT 133.130 745.720 136.890 746.370 ;
        RECT 137.730 745.720 141.950 746.370 ;
        RECT 142.790 745.720 146.550 746.370 ;
        RECT 147.390 745.720 151.610 746.370 ;
        RECT 152.450 745.720 156.210 746.370 ;
        RECT 157.050 745.720 161.270 746.370 ;
        RECT 162.110 745.720 165.870 746.370 ;
        RECT 166.710 745.720 170.930 746.370 ;
        RECT 171.770 745.720 175.530 746.370 ;
        RECT 176.370 745.720 180.590 746.370 ;
        RECT 181.430 745.720 185.190 746.370 ;
        RECT 186.030 745.720 190.250 746.370 ;
        RECT 191.090 745.720 194.850 746.370 ;
        RECT 195.690 745.720 199.910 746.370 ;
        RECT 200.750 745.720 204.510 746.370 ;
        RECT 205.350 745.720 209.570 746.370 ;
        RECT 210.410 745.720 214.170 746.370 ;
        RECT 215.010 745.720 219.230 746.370 ;
        RECT 220.070 745.720 223.830 746.370 ;
        RECT 224.670 745.720 228.890 746.370 ;
        RECT 229.730 745.720 233.490 746.370 ;
        RECT 234.330 745.720 238.550 746.370 ;
        RECT 239.390 745.720 243.150 746.370 ;
        RECT 243.990 745.720 248.210 746.370 ;
        RECT 249.050 745.720 252.810 746.370 ;
        RECT 253.650 745.720 257.870 746.370 ;
        RECT 258.710 745.720 262.470 746.370 ;
        RECT 263.310 745.720 267.530 746.370 ;
        RECT 268.370 745.720 272.130 746.370 ;
        RECT 272.970 745.720 277.190 746.370 ;
        RECT 278.030 745.720 281.790 746.370 ;
        RECT 282.630 745.720 286.390 746.370 ;
        RECT 287.230 745.720 291.450 746.370 ;
        RECT 292.290 745.720 296.050 746.370 ;
        RECT 296.890 745.720 301.110 746.370 ;
        RECT 301.950 745.720 305.710 746.370 ;
        RECT 306.550 745.720 310.770 746.370 ;
        RECT 311.610 745.720 315.370 746.370 ;
        RECT 316.210 745.720 320.430 746.370 ;
        RECT 321.270 745.720 325.030 746.370 ;
        RECT 325.870 745.720 330.090 746.370 ;
        RECT 330.930 745.720 334.690 746.370 ;
        RECT 335.530 745.720 339.750 746.370 ;
        RECT 340.590 745.720 344.350 746.370 ;
        RECT 345.190 745.720 349.410 746.370 ;
        RECT 350.250 745.720 354.010 746.370 ;
        RECT 354.850 745.720 359.070 746.370 ;
        RECT 359.910 745.720 363.670 746.370 ;
        RECT 364.510 745.720 368.730 746.370 ;
        RECT 369.570 745.720 373.330 746.370 ;
        RECT 374.170 745.720 378.390 746.370 ;
        RECT 379.230 745.720 382.990 746.370 ;
        RECT 383.830 745.720 388.050 746.370 ;
        RECT 388.890 745.720 392.650 746.370 ;
        RECT 393.490 745.720 397.710 746.370 ;
        RECT 398.550 745.720 402.310 746.370 ;
        RECT 403.150 745.720 407.370 746.370 ;
        RECT 408.210 745.720 411.970 746.370 ;
        RECT 412.810 745.720 417.030 746.370 ;
        RECT 417.870 745.720 421.630 746.370 ;
        RECT 422.470 745.720 426.690 746.370 ;
        RECT 427.530 745.720 431.290 746.370 ;
        RECT 432.130 745.720 436.350 746.370 ;
        RECT 437.190 745.720 440.950 746.370 ;
        RECT 441.790 745.720 446.010 746.370 ;
        RECT 446.850 745.720 450.610 746.370 ;
        RECT 451.450 745.720 455.670 746.370 ;
        RECT 456.510 745.720 460.270 746.370 ;
        RECT 461.110 745.720 465.330 746.370 ;
        RECT 466.170 745.720 469.930 746.370 ;
        RECT 470.770 745.720 474.990 746.370 ;
        RECT 475.830 745.720 479.590 746.370 ;
        RECT 480.430 745.720 484.650 746.370 ;
        RECT 485.490 745.720 489.250 746.370 ;
        RECT 490.090 745.720 494.310 746.370 ;
        RECT 495.150 745.720 498.910 746.370 ;
        RECT 499.750 745.720 503.970 746.370 ;
        RECT 504.810 745.720 508.570 746.370 ;
        RECT 509.410 745.720 513.630 746.370 ;
        RECT 514.470 745.720 518.230 746.370 ;
        RECT 519.070 745.720 523.290 746.370 ;
        RECT 524.130 745.720 527.890 746.370 ;
        RECT 528.730 745.720 532.950 746.370 ;
        RECT 533.790 745.720 537.550 746.370 ;
        RECT 538.390 745.720 542.610 746.370 ;
        RECT 543.450 745.720 547.210 746.370 ;
        RECT 2.400 3.555 547.760 745.720 ;
      LAYER met3 ;
        RECT 4.400 744.920 546.000 745.785 ;
        RECT 4.000 738.840 546.000 744.920 ;
        RECT 4.400 737.440 546.000 738.840 ;
        RECT 4.000 731.360 546.000 737.440 ;
        RECT 4.400 729.960 546.000 731.360 ;
        RECT 4.000 723.880 546.000 729.960 ;
        RECT 4.400 722.480 546.000 723.880 ;
        RECT 4.000 716.400 546.000 722.480 ;
        RECT 4.400 715.000 546.000 716.400 ;
        RECT 4.000 708.920 546.000 715.000 ;
        RECT 4.400 707.520 546.000 708.920 ;
        RECT 4.000 701.440 546.000 707.520 ;
        RECT 4.400 700.040 546.000 701.440 ;
        RECT 4.000 693.280 546.000 700.040 ;
        RECT 4.400 691.880 546.000 693.280 ;
        RECT 4.000 685.800 546.000 691.880 ;
        RECT 4.400 684.400 546.000 685.800 ;
        RECT 4.000 678.320 546.000 684.400 ;
        RECT 4.400 676.920 546.000 678.320 ;
        RECT 4.000 670.840 546.000 676.920 ;
        RECT 4.400 669.440 546.000 670.840 ;
        RECT 4.000 663.360 546.000 669.440 ;
        RECT 4.400 661.960 546.000 663.360 ;
        RECT 4.000 655.880 546.000 661.960 ;
        RECT 4.400 654.480 546.000 655.880 ;
        RECT 4.000 648.400 546.000 654.480 ;
        RECT 4.400 647.000 546.000 648.400 ;
        RECT 4.000 640.240 546.000 647.000 ;
        RECT 4.400 638.840 546.000 640.240 ;
        RECT 4.000 632.760 546.000 638.840 ;
        RECT 4.400 631.360 546.000 632.760 ;
        RECT 4.000 625.280 546.000 631.360 ;
        RECT 4.400 623.880 546.000 625.280 ;
        RECT 4.000 617.800 546.000 623.880 ;
        RECT 4.400 616.400 546.000 617.800 ;
        RECT 4.000 610.320 546.000 616.400 ;
        RECT 4.400 608.920 546.000 610.320 ;
        RECT 4.000 602.840 546.000 608.920 ;
        RECT 4.400 601.440 546.000 602.840 ;
        RECT 4.000 595.360 546.000 601.440 ;
        RECT 4.400 593.960 546.000 595.360 ;
        RECT 4.000 587.200 546.000 593.960 ;
        RECT 4.400 585.800 546.000 587.200 ;
        RECT 4.000 579.720 546.000 585.800 ;
        RECT 4.400 578.320 546.000 579.720 ;
        RECT 4.000 572.240 546.000 578.320 ;
        RECT 4.400 570.840 546.000 572.240 ;
        RECT 4.000 564.760 546.000 570.840 ;
        RECT 4.400 563.360 546.000 564.760 ;
        RECT 4.000 562.720 546.000 563.360 ;
        RECT 4.000 561.320 545.600 562.720 ;
        RECT 4.000 557.280 546.000 561.320 ;
        RECT 4.400 555.880 546.000 557.280 ;
        RECT 4.000 549.800 546.000 555.880 ;
        RECT 4.400 548.400 546.000 549.800 ;
        RECT 4.000 542.320 546.000 548.400 ;
        RECT 4.400 540.920 546.000 542.320 ;
        RECT 4.000 534.160 546.000 540.920 ;
        RECT 4.400 532.760 546.000 534.160 ;
        RECT 4.000 526.680 546.000 532.760 ;
        RECT 4.400 525.280 546.000 526.680 ;
        RECT 4.000 519.200 546.000 525.280 ;
        RECT 4.400 517.800 546.000 519.200 ;
        RECT 4.000 511.720 546.000 517.800 ;
        RECT 4.400 510.320 546.000 511.720 ;
        RECT 4.000 504.240 546.000 510.320 ;
        RECT 4.400 502.840 546.000 504.240 ;
        RECT 4.000 496.760 546.000 502.840 ;
        RECT 4.400 495.360 546.000 496.760 ;
        RECT 4.000 489.280 546.000 495.360 ;
        RECT 4.400 487.880 546.000 489.280 ;
        RECT 4.000 481.120 546.000 487.880 ;
        RECT 4.400 479.720 546.000 481.120 ;
        RECT 4.000 473.640 546.000 479.720 ;
        RECT 4.400 472.240 546.000 473.640 ;
        RECT 4.000 466.160 546.000 472.240 ;
        RECT 4.400 464.760 546.000 466.160 ;
        RECT 4.000 458.680 546.000 464.760 ;
        RECT 4.400 457.280 546.000 458.680 ;
        RECT 4.000 451.200 546.000 457.280 ;
        RECT 4.400 449.800 546.000 451.200 ;
        RECT 4.000 443.720 546.000 449.800 ;
        RECT 4.400 442.320 546.000 443.720 ;
        RECT 4.000 436.240 546.000 442.320 ;
        RECT 4.400 434.840 546.000 436.240 ;
        RECT 4.000 428.080 546.000 434.840 ;
        RECT 4.400 426.680 546.000 428.080 ;
        RECT 4.000 420.600 546.000 426.680 ;
        RECT 4.400 419.200 546.000 420.600 ;
        RECT 4.000 413.120 546.000 419.200 ;
        RECT 4.400 411.720 546.000 413.120 ;
        RECT 4.000 405.640 546.000 411.720 ;
        RECT 4.400 404.240 546.000 405.640 ;
        RECT 4.000 398.160 546.000 404.240 ;
        RECT 4.400 396.760 546.000 398.160 ;
        RECT 4.000 390.680 546.000 396.760 ;
        RECT 4.400 389.280 546.000 390.680 ;
        RECT 4.000 383.200 546.000 389.280 ;
        RECT 4.400 381.800 546.000 383.200 ;
        RECT 4.000 375.040 546.000 381.800 ;
        RECT 4.400 373.640 546.000 375.040 ;
        RECT 4.000 367.560 546.000 373.640 ;
        RECT 4.400 366.160 546.000 367.560 ;
        RECT 4.000 360.080 546.000 366.160 ;
        RECT 4.400 358.680 546.000 360.080 ;
        RECT 4.000 352.600 546.000 358.680 ;
        RECT 4.400 351.200 546.000 352.600 ;
        RECT 4.000 345.120 546.000 351.200 ;
        RECT 4.400 343.720 546.000 345.120 ;
        RECT 4.000 337.640 546.000 343.720 ;
        RECT 4.400 336.240 546.000 337.640 ;
        RECT 4.000 330.160 546.000 336.240 ;
        RECT 4.400 328.760 546.000 330.160 ;
        RECT 4.000 322.000 546.000 328.760 ;
        RECT 4.400 320.600 546.000 322.000 ;
        RECT 4.000 314.520 546.000 320.600 ;
        RECT 4.400 313.120 546.000 314.520 ;
        RECT 4.000 307.040 546.000 313.120 ;
        RECT 4.400 305.640 546.000 307.040 ;
        RECT 4.000 299.560 546.000 305.640 ;
        RECT 4.400 298.160 546.000 299.560 ;
        RECT 4.000 292.080 546.000 298.160 ;
        RECT 4.400 290.680 546.000 292.080 ;
        RECT 4.000 284.600 546.000 290.680 ;
        RECT 4.400 283.200 546.000 284.600 ;
        RECT 4.000 277.120 546.000 283.200 ;
        RECT 4.400 275.720 546.000 277.120 ;
        RECT 4.000 268.960 546.000 275.720 ;
        RECT 4.400 267.560 546.000 268.960 ;
        RECT 4.000 261.480 546.000 267.560 ;
        RECT 4.400 260.080 546.000 261.480 ;
        RECT 4.000 254.000 546.000 260.080 ;
        RECT 4.400 252.600 546.000 254.000 ;
        RECT 4.000 246.520 546.000 252.600 ;
        RECT 4.400 245.120 546.000 246.520 ;
        RECT 4.000 239.040 546.000 245.120 ;
        RECT 4.400 237.640 546.000 239.040 ;
        RECT 4.000 231.560 546.000 237.640 ;
        RECT 4.400 230.160 546.000 231.560 ;
        RECT 4.000 224.080 546.000 230.160 ;
        RECT 4.400 222.680 546.000 224.080 ;
        RECT 4.000 215.920 546.000 222.680 ;
        RECT 4.400 214.520 546.000 215.920 ;
        RECT 4.000 208.440 546.000 214.520 ;
        RECT 4.400 207.040 546.000 208.440 ;
        RECT 4.000 200.960 546.000 207.040 ;
        RECT 4.400 199.560 546.000 200.960 ;
        RECT 4.000 193.480 546.000 199.560 ;
        RECT 4.400 192.080 546.000 193.480 ;
        RECT 4.000 188.040 546.000 192.080 ;
        RECT 4.000 186.640 545.600 188.040 ;
        RECT 4.000 186.000 546.000 186.640 ;
        RECT 4.400 184.600 546.000 186.000 ;
        RECT 4.000 178.520 546.000 184.600 ;
        RECT 4.400 177.120 546.000 178.520 ;
        RECT 4.000 171.040 546.000 177.120 ;
        RECT 4.400 169.640 546.000 171.040 ;
        RECT 4.000 162.880 546.000 169.640 ;
        RECT 4.400 161.480 546.000 162.880 ;
        RECT 4.000 155.400 546.000 161.480 ;
        RECT 4.400 154.000 546.000 155.400 ;
        RECT 4.000 147.920 546.000 154.000 ;
        RECT 4.400 146.520 546.000 147.920 ;
        RECT 4.000 140.440 546.000 146.520 ;
        RECT 4.400 139.040 546.000 140.440 ;
        RECT 4.000 132.960 546.000 139.040 ;
        RECT 4.400 131.560 546.000 132.960 ;
        RECT 4.000 125.480 546.000 131.560 ;
        RECT 4.400 124.080 546.000 125.480 ;
        RECT 4.000 118.000 546.000 124.080 ;
        RECT 4.400 116.600 546.000 118.000 ;
        RECT 4.000 109.840 546.000 116.600 ;
        RECT 4.400 108.440 546.000 109.840 ;
        RECT 4.000 102.360 546.000 108.440 ;
        RECT 4.400 100.960 546.000 102.360 ;
        RECT 4.000 94.880 546.000 100.960 ;
        RECT 4.400 93.480 546.000 94.880 ;
        RECT 4.000 87.400 546.000 93.480 ;
        RECT 4.400 86.000 546.000 87.400 ;
        RECT 4.000 79.920 546.000 86.000 ;
        RECT 4.400 78.520 546.000 79.920 ;
        RECT 4.000 72.440 546.000 78.520 ;
        RECT 4.400 71.040 546.000 72.440 ;
        RECT 4.000 64.960 546.000 71.040 ;
        RECT 4.400 63.560 546.000 64.960 ;
        RECT 4.000 56.800 546.000 63.560 ;
        RECT 4.400 55.400 546.000 56.800 ;
        RECT 4.000 49.320 546.000 55.400 ;
        RECT 4.400 47.920 546.000 49.320 ;
        RECT 4.000 41.840 546.000 47.920 ;
        RECT 4.400 40.440 546.000 41.840 ;
        RECT 4.000 34.360 546.000 40.440 ;
        RECT 4.400 32.960 546.000 34.360 ;
        RECT 4.000 26.880 546.000 32.960 ;
        RECT 4.400 25.480 546.000 26.880 ;
        RECT 4.000 19.400 546.000 25.480 ;
        RECT 4.400 18.000 546.000 19.400 ;
        RECT 4.000 11.920 546.000 18.000 ;
        RECT 4.400 10.520 546.000 11.920 ;
        RECT 4.000 4.440 546.000 10.520 ;
        RECT 4.400 3.575 546.000 4.440 ;
      LAYER met4 ;
        RECT 8.575 19.895 20.640 735.585 ;
        RECT 23.040 19.895 97.440 735.585 ;
        RECT 99.840 19.895 174.240 735.585 ;
        RECT 176.640 19.895 251.040 735.585 ;
        RECT 253.440 19.895 327.840 735.585 ;
        RECT 330.240 19.895 404.640 735.585 ;
        RECT 407.040 19.895 481.440 735.585 ;
        RECT 483.840 19.895 529.625 735.585 ;
  END
END Peripherals
END LIBRARY

