magic
tech sky130A
magscale 1 2
timestamp 1654452354
<< viali >>
rect 2329 39593 2363 39627
rect 3065 39593 3099 39627
rect 3985 39593 4019 39627
rect 27169 39593 27203 39627
rect 41429 39593 41463 39627
rect 48973 39593 49007 39627
rect 56425 39593 56459 39627
rect 19257 39457 19291 39491
rect 1409 39389 1443 39423
rect 2145 39389 2179 39423
rect 2881 39389 2915 39423
rect 3801 39389 3835 39423
rect 26985 39389 27019 39423
rect 33793 39389 33827 39423
rect 56241 39389 56275 39423
rect 1593 39253 1627 39287
rect 4445 39253 4479 39287
rect 33977 39253 34011 39287
rect 35081 39049 35115 39083
rect 1409 38913 1443 38947
rect 35265 38913 35299 38947
rect 1593 38709 1627 38743
rect 1593 38505 1627 38539
rect 1409 38301 1443 38335
rect 1409 37825 1443 37859
rect 1593 37621 1627 37655
rect 1409 36737 1443 36771
rect 1593 36601 1627 36635
rect 1409 36125 1443 36159
rect 1593 35989 1627 36023
rect 1869 34969 1903 35003
rect 1961 34901 1995 34935
rect 1593 34697 1627 34731
rect 2145 34697 2179 34731
rect 1409 34561 1443 34595
rect 2329 34561 2363 34595
rect 1409 33949 1443 33983
rect 1593 33813 1627 33847
rect 1869 33473 1903 33507
rect 2881 33473 2915 33507
rect 2053 33337 2087 33371
rect 2697 33269 2731 33303
rect 1409 32861 1443 32895
rect 1593 32725 1627 32759
rect 1409 32385 1443 32419
rect 1593 32181 1627 32215
rect 1409 31909 1443 31943
rect 1593 31773 1627 31807
rect 1869 31297 1903 31331
rect 2145 31093 2179 31127
rect 1593 30889 1627 30923
rect 2145 30821 2179 30855
rect 1409 30685 1443 30719
rect 2329 30685 2363 30719
rect 2973 30685 3007 30719
rect 4813 30685 4847 30719
rect 2789 30549 2823 30583
rect 4629 30549 4663 30583
rect 2789 30345 2823 30379
rect 1409 30209 1443 30243
rect 2697 30209 2731 30243
rect 4712 30209 4746 30243
rect 2973 30141 3007 30175
rect 4445 30141 4479 30175
rect 1593 30005 1627 30039
rect 2329 30005 2363 30039
rect 5825 30005 5859 30039
rect 6837 29801 6871 29835
rect 7205 29801 7239 29835
rect 4261 29733 4295 29767
rect 4813 29665 4847 29699
rect 1869 29597 1903 29631
rect 4629 29597 4663 29631
rect 4721 29597 4755 29631
rect 6929 29597 6963 29631
rect 7021 29597 7055 29631
rect 7941 29597 7975 29631
rect 2136 29529 2170 29563
rect 6745 29529 6779 29563
rect 3249 29461 3283 29495
rect 7757 29461 7791 29495
rect 3433 29257 3467 29291
rect 8217 29257 8251 29291
rect 1869 29189 1903 29223
rect 2697 29121 2731 29155
rect 3617 29121 3651 29155
rect 4261 29121 4295 29155
rect 7104 29121 7138 29155
rect 6837 29053 6871 29087
rect 2145 28985 2179 29019
rect 2881 28985 2915 29019
rect 4077 28985 4111 29019
rect 3893 28713 3927 28747
rect 6929 28713 6963 28747
rect 15485 28713 15519 28747
rect 4537 28577 4571 28611
rect 7389 28577 7423 28611
rect 7573 28577 7607 28611
rect 4353 28509 4387 28543
rect 7297 28509 7331 28543
rect 10701 28509 10735 28543
rect 10885 28509 10919 28543
rect 10977 28509 11011 28543
rect 14105 28509 14139 28543
rect 16681 28509 16715 28543
rect 1869 28441 1903 28475
rect 14372 28441 14406 28475
rect 16948 28441 16982 28475
rect 2145 28373 2179 28407
rect 4261 28373 4295 28407
rect 10517 28373 10551 28407
rect 18061 28373 18095 28407
rect 13829 28169 13863 28203
rect 14657 28169 14691 28203
rect 15025 28169 15059 28203
rect 17049 28169 17083 28203
rect 17417 28169 17451 28203
rect 4436 28101 4470 28135
rect 9864 28101 9898 28135
rect 1409 28033 1443 28067
rect 2421 28033 2455 28067
rect 3065 28033 3099 28067
rect 4169 28033 4203 28067
rect 6837 28033 6871 28067
rect 9597 28033 9631 28067
rect 12449 28033 12483 28067
rect 12716 28033 12750 28067
rect 14841 28033 14875 28067
rect 15117 28033 15151 28067
rect 17233 28033 17267 28067
rect 17509 28033 17543 28067
rect 5549 27897 5583 27931
rect 10977 27897 11011 27931
rect 1593 27829 1627 27863
rect 2237 27829 2271 27863
rect 2881 27829 2915 27863
rect 6653 27829 6687 27863
rect 6745 27625 6779 27659
rect 12909 27625 12943 27659
rect 7205 27489 7239 27523
rect 7389 27489 7423 27523
rect 9689 27489 9723 27523
rect 1869 27421 1903 27455
rect 2136 27421 2170 27455
rect 13093 27421 13127 27455
rect 13369 27421 13403 27455
rect 9956 27353 9990 27387
rect 13277 27353 13311 27387
rect 3249 27285 3283 27319
rect 7113 27285 7147 27319
rect 11069 27285 11103 27319
rect 2329 27081 2363 27115
rect 2789 27081 2823 27115
rect 7757 27081 7791 27115
rect 10517 27081 10551 27115
rect 10885 27081 10919 27115
rect 1501 27013 1535 27047
rect 2697 27013 2731 27047
rect 6644 27013 6678 27047
rect 17049 27013 17083 27047
rect 3709 26945 3743 26979
rect 10701 26945 10735 26979
rect 10977 26945 11011 26979
rect 16865 26945 16899 26979
rect 17141 26945 17175 26979
rect 2973 26877 3007 26911
rect 6377 26877 6411 26911
rect 1777 26809 1811 26843
rect 3525 26741 3559 26775
rect 16681 26741 16715 26775
rect 5181 26537 5215 26571
rect 16681 26537 16715 26571
rect 18521 26537 18555 26571
rect 3065 26469 3099 26503
rect 1409 26333 1443 26367
rect 2145 26333 2179 26367
rect 3249 26333 3283 26367
rect 3801 26333 3835 26367
rect 4057 26333 4091 26367
rect 15301 26333 15335 26367
rect 15568 26333 15602 26367
rect 17141 26333 17175 26367
rect 17408 26265 17442 26299
rect 1593 26197 1627 26231
rect 2329 26197 2363 26231
rect 3065 25993 3099 26027
rect 3525 25993 3559 26027
rect 8769 25993 8803 26027
rect 13921 25993 13955 26027
rect 17325 25993 17359 26027
rect 17693 25993 17727 26027
rect 3433 25925 3467 25959
rect 4629 25925 4663 25959
rect 1409 25857 1443 25891
rect 2329 25857 2363 25891
rect 4445 25857 4479 25891
rect 7389 25857 7423 25891
rect 7656 25857 7690 25891
rect 9597 25857 9631 25891
rect 9864 25857 9898 25891
rect 12541 25857 12575 25891
rect 12808 25857 12842 25891
rect 14637 25857 14671 25891
rect 17509 25857 17543 25891
rect 17785 25857 17819 25891
rect 3709 25789 3743 25823
rect 14381 25789 14415 25823
rect 1593 25721 1627 25755
rect 2145 25653 2179 25687
rect 10977 25653 11011 25687
rect 15761 25653 15795 25687
rect 9597 25449 9631 25483
rect 10885 25449 10919 25483
rect 13093 25449 13127 25483
rect 7297 25381 7331 25415
rect 1869 25313 1903 25347
rect 5917 25313 5951 25347
rect 8953 25245 8987 25279
rect 9046 25245 9080 25279
rect 9321 25245 9355 25279
rect 9459 25245 9493 25279
rect 10241 25245 10275 25279
rect 10389 25245 10423 25279
rect 10517 25245 10551 25279
rect 10609 25245 10643 25279
rect 10706 25245 10740 25279
rect 12449 25245 12483 25279
rect 12542 25245 12576 25279
rect 12817 25245 12851 25279
rect 12914 25245 12948 25279
rect 17141 25245 17175 25279
rect 17417 25245 17451 25279
rect 2136 25177 2170 25211
rect 6184 25177 6218 25211
rect 7849 25177 7883 25211
rect 9229 25177 9263 25211
rect 12173 25177 12207 25211
rect 12725 25177 12759 25211
rect 17325 25177 17359 25211
rect 3249 25109 3283 25143
rect 8125 25109 8159 25143
rect 16957 25109 16991 25143
rect 2329 24905 2363 24939
rect 1685 24837 1719 24871
rect 9045 24837 9079 24871
rect 16948 24837 16982 24871
rect 1409 24769 1443 24803
rect 2513 24769 2547 24803
rect 3157 24769 3191 24803
rect 3801 24769 3835 24803
rect 4077 24769 4111 24803
rect 8769 24769 8803 24803
rect 8862 24769 8896 24803
rect 9137 24769 9171 24803
rect 9275 24769 9309 24803
rect 11805 24769 11839 24803
rect 11989 24769 12023 24803
rect 12633 24769 12667 24803
rect 12726 24769 12760 24803
rect 12909 24769 12943 24803
rect 13001 24769 13035 24803
rect 13098 24769 13132 24803
rect 3893 24701 3927 24735
rect 12357 24701 12391 24735
rect 16681 24701 16715 24735
rect 13277 24633 13311 24667
rect 2973 24565 3007 24599
rect 3801 24565 3835 24599
rect 4261 24565 4295 24599
rect 9413 24565 9447 24599
rect 18061 24565 18095 24599
rect 2237 24361 2271 24395
rect 5181 24361 5215 24395
rect 2697 24225 2731 24259
rect 2881 24225 2915 24259
rect 12817 24225 12851 24259
rect 1409 24157 1443 24191
rect 2605 24157 2639 24191
rect 3808 24157 3842 24191
rect 12541 24157 12575 24191
rect 15485 24157 15519 24191
rect 4068 24089 4102 24123
rect 14565 24089 14599 24123
rect 14749 24089 14783 24123
rect 15752 24089 15786 24123
rect 1593 24021 1627 24055
rect 16865 24021 16899 24055
rect 2421 23817 2455 23851
rect 3433 23817 3467 23851
rect 8861 23817 8895 23851
rect 9965 23817 9999 23851
rect 15669 23817 15703 23851
rect 7748 23749 7782 23783
rect 10793 23749 10827 23783
rect 16037 23749 16071 23783
rect 1409 23681 1443 23715
rect 2605 23681 2639 23715
rect 4353 23681 4387 23715
rect 9321 23681 9355 23715
rect 9414 23681 9448 23715
rect 9597 23681 9631 23715
rect 9689 23681 9723 23715
rect 9827 23681 9861 23715
rect 11529 23681 11563 23715
rect 11796 23681 11830 23715
rect 15853 23681 15887 23715
rect 16129 23681 16163 23715
rect 3525 23613 3559 23647
rect 3617 23613 3651 23647
rect 7481 23613 7515 23647
rect 3065 23545 3099 23579
rect 4537 23545 4571 23579
rect 10977 23545 11011 23579
rect 1593 23477 1627 23511
rect 12909 23477 12943 23511
rect 2053 23273 2087 23307
rect 8401 23273 8435 23307
rect 11897 23273 11931 23307
rect 14105 23137 14139 23171
rect 17417 23137 17451 23171
rect 17509 23137 17543 23171
rect 1593 23069 1627 23103
rect 2237 23069 2271 23103
rect 7021 23069 7055 23103
rect 10517 23069 10551 23103
rect 11253 23069 11287 23103
rect 11346 23069 11380 23103
rect 11618 23069 11652 23103
rect 11718 23069 11752 23103
rect 17325 23069 17359 23103
rect 17601 23069 17635 23103
rect 19993 23069 20027 23103
rect 24409 23069 24443 23103
rect 27629 23069 27663 23103
rect 33241 23069 33275 23103
rect 33517 23069 33551 23103
rect 7288 23001 7322 23035
rect 11529 23001 11563 23035
rect 14350 23001 14384 23035
rect 20260 23001 20294 23035
rect 24676 23001 24710 23035
rect 27896 23001 27930 23035
rect 1409 22933 1443 22967
rect 10701 22933 10735 22967
rect 15485 22933 15519 22967
rect 17141 22933 17175 22967
rect 21373 22933 21407 22967
rect 25789 22933 25823 22967
rect 29009 22933 29043 22967
rect 33057 22933 33091 22967
rect 33425 22933 33459 22967
rect 2973 22729 3007 22763
rect 5181 22729 5215 22763
rect 9321 22729 9355 22763
rect 14105 22729 14139 22763
rect 14473 22729 14507 22763
rect 17601 22729 17635 22763
rect 20821 22729 20855 22763
rect 24685 22729 24719 22763
rect 25053 22729 25087 22763
rect 27997 22729 28031 22763
rect 28365 22729 28399 22763
rect 13461 22661 13495 22695
rect 21189 22661 21223 22695
rect 33302 22661 33336 22695
rect 1409 22593 1443 22627
rect 3065 22593 3099 22627
rect 3801 22593 3835 22627
rect 4057 22593 4091 22627
rect 8677 22593 8711 22627
rect 8825 22593 8859 22627
rect 8953 22593 8987 22627
rect 9045 22593 9079 22627
rect 9183 22593 9217 22627
rect 13645 22593 13679 22627
rect 14289 22593 14323 22627
rect 14565 22593 14599 22627
rect 17877 22593 17911 22627
rect 18061 22593 18095 22627
rect 21005 22593 21039 22627
rect 21281 22593 21315 22627
rect 24869 22593 24903 22627
rect 25145 22593 25179 22627
rect 28181 22593 28215 22627
rect 28457 22593 28491 22627
rect 30472 22593 30506 22627
rect 3157 22525 3191 22559
rect 17785 22525 17819 22559
rect 17969 22525 18003 22559
rect 30205 22525 30239 22559
rect 33057 22525 33091 22559
rect 1593 22389 1627 22423
rect 2605 22389 2639 22423
rect 31585 22389 31619 22423
rect 34437 22389 34471 22423
rect 3801 22185 3835 22219
rect 17785 22185 17819 22219
rect 25513 22185 25547 22219
rect 25697 22185 25731 22219
rect 30849 22185 30883 22219
rect 33241 22185 33275 22219
rect 2053 22049 2087 22083
rect 15761 22049 15795 22083
rect 15945 22049 15979 22083
rect 16129 22049 16163 22083
rect 16958 22049 16992 22083
rect 17233 22049 17267 22083
rect 17969 22049 18003 22083
rect 18153 22049 18187 22083
rect 20453 22049 20487 22083
rect 29653 22049 29687 22083
rect 31125 22049 31159 22083
rect 32229 22049 32263 22083
rect 32873 22049 32907 22083
rect 1869 21981 1903 22015
rect 2881 21981 2915 22015
rect 3985 21981 4019 22015
rect 11345 21981 11379 22015
rect 11621 21981 11655 22015
rect 16037 21981 16071 22015
rect 16221 21981 16255 22015
rect 17049 21981 17083 22015
rect 17141 21981 17175 22015
rect 18061 21981 18095 22015
rect 18245 21981 18279 22015
rect 22477 21981 22511 22015
rect 24593 21981 24627 22015
rect 24869 21981 24903 22015
rect 29561 21981 29595 22015
rect 29745 21981 29779 22015
rect 31033 21981 31067 22015
rect 31217 21981 31251 22015
rect 31309 21981 31343 22015
rect 32965 21981 32999 22015
rect 20720 21913 20754 21947
rect 22744 21913 22778 21947
rect 24409 21913 24443 21947
rect 25329 21913 25363 21947
rect 31861 21913 31895 21947
rect 32045 21913 32079 21947
rect 2697 21845 2731 21879
rect 16773 21845 16807 21879
rect 21833 21845 21867 21879
rect 23857 21845 23891 21879
rect 24777 21845 24811 21879
rect 25529 21845 25563 21879
rect 7665 21641 7699 21675
rect 10885 21641 10919 21675
rect 17141 21641 17175 21675
rect 21833 21641 21867 21675
rect 22201 21641 22235 21675
rect 26157 21641 26191 21675
rect 29561 21641 29595 21675
rect 32505 21641 32539 21675
rect 2942 21573 2976 21607
rect 4905 21573 4939 21607
rect 24777 21573 24811 21607
rect 24993 21573 25027 21607
rect 25789 21573 25823 21607
rect 26019 21539 26053 21573
rect 1409 21505 1443 21539
rect 5089 21505 5123 21539
rect 7481 21505 7515 21539
rect 7757 21505 7791 21539
rect 9772 21505 9806 21539
rect 14105 21505 14139 21539
rect 17325 21505 17359 21539
rect 17417 21505 17451 21539
rect 18429 21505 18463 21539
rect 18521 21505 18555 21539
rect 22017 21505 22051 21539
rect 22293 21505 22327 21539
rect 27896 21505 27930 21539
rect 29469 21505 29503 21539
rect 29653 21505 29687 21539
rect 32321 21505 32355 21539
rect 32505 21505 32539 21539
rect 35265 21505 35299 21539
rect 2697 21437 2731 21471
rect 9505 21437 9539 21471
rect 17509 21437 17543 21471
rect 17601 21437 17635 21471
rect 18337 21437 18371 21471
rect 18613 21437 18647 21471
rect 27629 21437 27663 21471
rect 1593 21301 1627 21335
rect 4077 21301 4111 21335
rect 5273 21301 5307 21335
rect 7297 21301 7331 21335
rect 14197 21301 14231 21335
rect 18153 21301 18187 21335
rect 24685 21301 24719 21335
rect 24961 21301 24995 21335
rect 25145 21301 25179 21335
rect 25513 21301 25547 21335
rect 25973 21301 26007 21335
rect 29009 21301 29043 21335
rect 35081 21301 35115 21335
rect 2513 21097 2547 21131
rect 7665 21097 7699 21131
rect 10149 21097 10183 21131
rect 19257 21097 19291 21131
rect 27905 21097 27939 21131
rect 36553 21097 36587 21131
rect 1961 21029 1995 21063
rect 15117 21029 15151 21063
rect 17785 21029 17819 21063
rect 2973 20961 3007 20995
rect 3157 20961 3191 20995
rect 14473 20961 14507 20995
rect 15393 20961 15427 20995
rect 15485 20961 15519 20995
rect 18153 20961 18187 20995
rect 19441 20961 19475 20995
rect 19625 20961 19659 20995
rect 19717 20961 19751 20995
rect 33425 20961 33459 20995
rect 33609 20961 33643 20995
rect 35173 20961 35207 20995
rect 2881 20893 2915 20927
rect 6285 20893 6319 20927
rect 6552 20893 6586 20927
rect 10333 20893 10367 20927
rect 10609 20893 10643 20927
rect 11805 20893 11839 20927
rect 13277 20893 13311 20927
rect 13553 20893 13587 20927
rect 14289 20893 14323 20927
rect 14382 20893 14416 20927
rect 14565 20893 14599 20927
rect 15301 20893 15335 20927
rect 15577 20893 15611 20927
rect 17969 20893 18003 20927
rect 18061 20893 18095 20927
rect 18245 20893 18279 20927
rect 19533 20893 19567 20927
rect 28089 20893 28123 20927
rect 28273 20893 28307 20927
rect 28365 20893 28399 20927
rect 28825 20893 28859 20927
rect 29009 20893 29043 20927
rect 33333 20893 33367 20927
rect 33517 20893 33551 20927
rect 35440 20893 35474 20927
rect 37381 20893 37415 20927
rect 37657 20893 37691 20927
rect 1685 20825 1719 20859
rect 10517 20825 10551 20859
rect 28917 20825 28951 20859
rect 11989 20757 12023 20791
rect 13093 20757 13127 20791
rect 13461 20757 13495 20791
rect 14105 20757 14139 20791
rect 33149 20757 33183 20791
rect 37197 20757 37231 20791
rect 37565 20757 37599 20791
rect 2973 20553 3007 20587
rect 3709 20553 3743 20587
rect 8493 20553 8527 20587
rect 14105 20553 14139 20587
rect 15485 20553 15519 20587
rect 18613 20553 18647 20587
rect 33057 20553 33091 20587
rect 33701 20553 33735 20587
rect 33885 20553 33919 20587
rect 34897 20553 34931 20587
rect 12992 20485 13026 20519
rect 25237 20485 25271 20519
rect 25421 20485 25455 20519
rect 28733 20485 28767 20519
rect 28933 20485 28967 20519
rect 32689 20485 32723 20519
rect 33517 20485 33551 20519
rect 37626 20485 37660 20519
rect 1409 20417 1443 20451
rect 2881 20417 2915 20451
rect 3893 20417 3927 20451
rect 7380 20417 7414 20451
rect 12725 20417 12759 20451
rect 15669 20417 15703 20451
rect 15853 20417 15887 20451
rect 15945 20417 15979 20451
rect 17601 20417 17635 20451
rect 18798 20417 18832 20451
rect 18889 20417 18923 20451
rect 19901 20417 19935 20451
rect 20168 20417 20202 20451
rect 23029 20417 23063 20451
rect 23296 20417 23330 20451
rect 25697 20417 25731 20451
rect 32420 20417 32454 20451
rect 32506 20417 32540 20451
rect 32781 20417 32815 20451
rect 32919 20417 32953 20451
rect 33793 20417 33827 20451
rect 34529 20417 34563 20451
rect 34713 20417 34747 20451
rect 3157 20349 3191 20383
rect 7113 20349 7147 20383
rect 15761 20349 15795 20383
rect 17325 20349 17359 20383
rect 18981 20349 19015 20383
rect 19073 20349 19107 20383
rect 37381 20349 37415 20383
rect 24409 20281 24443 20315
rect 29101 20281 29135 20315
rect 1593 20213 1627 20247
rect 2513 20213 2547 20247
rect 21281 20213 21315 20247
rect 24869 20213 24903 20247
rect 25421 20213 25455 20247
rect 28917 20213 28951 20247
rect 34069 20213 34103 20247
rect 38761 20213 38795 20247
rect 7849 20009 7883 20043
rect 20729 20009 20763 20043
rect 22017 20009 22051 20043
rect 22201 20009 22235 20043
rect 23397 20009 23431 20043
rect 24961 20009 24995 20043
rect 28641 20009 28675 20043
rect 30113 20009 30147 20043
rect 32413 20009 32447 20043
rect 33517 20009 33551 20043
rect 37013 20009 37047 20043
rect 37565 20009 37599 20043
rect 10241 19873 10275 19907
rect 11989 19873 12023 19907
rect 15301 19873 15335 19907
rect 16589 19873 16623 19907
rect 37933 19873 37967 19907
rect 1409 19805 1443 19839
rect 2789 19805 2823 19839
rect 5089 19805 5123 19839
rect 8033 19805 8067 19839
rect 8309 19805 8343 19839
rect 11713 19805 11747 19839
rect 15025 19805 15059 19839
rect 16313 19805 16347 19839
rect 17601 19805 17635 19839
rect 17877 19805 17911 19839
rect 20913 19805 20947 19839
rect 21097 19805 21131 19839
rect 21189 19805 21223 19839
rect 23581 19805 23615 19839
rect 23765 19805 23799 19839
rect 23857 19805 23891 19839
rect 26525 19805 26559 19839
rect 28641 19805 28675 19839
rect 28917 19805 28951 19839
rect 29837 19805 29871 19839
rect 31769 19805 31803 19839
rect 31917 19805 31951 19839
rect 32045 19805 32079 19839
rect 32275 19805 32309 19839
rect 32873 19805 32907 19839
rect 33021 19805 33055 19839
rect 33338 19805 33372 19839
rect 36921 19805 36955 19839
rect 37105 19805 37139 19839
rect 37749 19805 37783 19839
rect 38025 19805 38059 19839
rect 10057 19737 10091 19771
rect 21465 19737 21499 19771
rect 21833 19737 21867 19771
rect 22049 19737 22083 19771
rect 24869 19737 24903 19771
rect 26792 19737 26826 19771
rect 29561 19737 29595 19771
rect 29929 19737 29963 19771
rect 32137 19737 32171 19771
rect 33149 19737 33183 19771
rect 33241 19737 33275 19771
rect 1593 19669 1627 19703
rect 2605 19669 2639 19703
rect 4905 19669 4939 19703
rect 8217 19669 8251 19703
rect 9689 19669 9723 19703
rect 10149 19669 10183 19703
rect 27905 19669 27939 19703
rect 28825 19669 28859 19703
rect 29745 19669 29779 19703
rect 3985 19465 4019 19499
rect 10977 19465 11011 19499
rect 14013 19465 14047 19499
rect 18337 19465 18371 19499
rect 22038 19465 22072 19499
rect 22201 19465 22235 19499
rect 24409 19465 24443 19499
rect 26985 19465 27019 19499
rect 33701 19465 33735 19499
rect 33885 19465 33919 19499
rect 2850 19397 2884 19431
rect 4712 19397 4746 19431
rect 21833 19397 21867 19431
rect 32413 19397 32447 19431
rect 1409 19329 1443 19363
rect 4445 19329 4479 19363
rect 9597 19329 9631 19363
rect 9864 19329 9898 19363
rect 13369 19329 13403 19363
rect 15209 19329 15243 19363
rect 15485 19329 15519 19363
rect 18613 19329 18647 19363
rect 24225 19329 24259 19363
rect 27445 19329 27479 19363
rect 27997 19329 28031 19363
rect 28181 19329 28215 19363
rect 28641 19329 28675 19363
rect 28917 19329 28951 19363
rect 32126 19329 32160 19363
rect 32230 19329 32264 19363
rect 32505 19329 32539 19363
rect 32643 19329 32677 19363
rect 33333 19329 33367 19363
rect 44097 19329 44131 19363
rect 2605 19261 2639 19295
rect 13553 19261 13587 19295
rect 14198 19261 14232 19295
rect 14290 19261 14324 19295
rect 14381 19261 14415 19295
rect 14473 19261 14507 19295
rect 15025 19261 15059 19295
rect 15301 19261 15335 19295
rect 15393 19261 15427 19295
rect 17049 19261 17083 19295
rect 17325 19261 17359 19295
rect 18522 19261 18556 19295
rect 18705 19261 18739 19295
rect 18797 19261 18831 19295
rect 27169 19261 27203 19295
rect 27261 19261 27295 19295
rect 27353 19261 27387 19295
rect 37841 19261 37875 19295
rect 38117 19261 38151 19295
rect 28089 19193 28123 19227
rect 32781 19193 32815 19227
rect 1593 19125 1627 19159
rect 5825 19125 5859 19159
rect 22017 19125 22051 19159
rect 33701 19125 33735 19159
rect 43913 19125 43947 19159
rect 2973 18921 3007 18955
rect 4905 18921 4939 18955
rect 15669 18921 15703 18955
rect 27537 18921 27571 18955
rect 33241 18921 33275 18955
rect 41245 18921 41279 18955
rect 9873 18853 9907 18887
rect 15853 18853 15887 18887
rect 1593 18785 1627 18819
rect 5549 18785 5583 18819
rect 14289 18785 14323 18819
rect 18429 18785 18463 18819
rect 18521 18785 18555 18819
rect 29837 18785 29871 18819
rect 39865 18785 39899 18819
rect 3985 18717 4019 18751
rect 7113 18717 7147 18751
rect 10057 18717 10091 18751
rect 11437 18717 11471 18751
rect 14565 18717 14599 18751
rect 16865 18717 16899 18751
rect 17141 18717 17175 18751
rect 18337 18717 18371 18751
rect 18613 18717 18647 18751
rect 27353 18717 27387 18751
rect 29561 18717 29595 18751
rect 32597 18717 32631 18751
rect 32745 18717 32779 18751
rect 33062 18717 33096 18751
rect 36645 18717 36679 18751
rect 36921 18717 36955 18751
rect 38117 18717 38151 18751
rect 38393 18717 38427 18751
rect 38853 18717 38887 18751
rect 39129 18717 39163 18751
rect 43085 18717 43119 18751
rect 43352 18717 43386 18751
rect 47501 18717 47535 18751
rect 1860 18649 1894 18683
rect 5365 18649 5399 18683
rect 11704 18649 11738 18683
rect 14473 18649 14507 18683
rect 15025 18649 15059 18683
rect 15485 18649 15519 18683
rect 27169 18649 27203 18683
rect 32873 18649 32907 18683
rect 32965 18649 32999 18683
rect 39037 18649 39071 18683
rect 40110 18649 40144 18683
rect 3801 18581 3835 18615
rect 5273 18581 5307 18615
rect 6929 18581 6963 18615
rect 12817 18581 12851 18615
rect 15695 18581 15729 18615
rect 18153 18581 18187 18615
rect 37933 18581 37967 18615
rect 38301 18581 38335 18615
rect 38945 18581 38979 18615
rect 44465 18581 44499 18615
rect 47317 18581 47351 18615
rect 1593 18377 1627 18411
rect 2329 18377 2363 18411
rect 2697 18377 2731 18411
rect 12633 18377 12667 18411
rect 14197 18377 14231 18411
rect 17233 18377 17267 18411
rect 19257 18377 19291 18411
rect 21005 18377 21039 18411
rect 35449 18377 35483 18411
rect 35541 18377 35575 18411
rect 43929 18377 43963 18411
rect 44097 18377 44131 18411
rect 53389 18377 53423 18411
rect 55413 18377 55447 18411
rect 7450 18309 7484 18343
rect 13001 18309 13035 18343
rect 20821 18309 20855 18343
rect 22201 18309 22235 18343
rect 27445 18309 27479 18343
rect 29837 18309 29871 18343
rect 34069 18309 34103 18343
rect 43729 18309 43763 18343
rect 47838 18309 47872 18343
rect 54278 18309 54312 18343
rect 1409 18241 1443 18275
rect 2513 18241 2547 18275
rect 2789 18241 2823 18275
rect 3433 18241 3467 18275
rect 6561 18241 6595 18275
rect 12817 18241 12851 18275
rect 13093 18241 13127 18275
rect 14473 18241 14507 18275
rect 14565 18241 14599 18275
rect 15301 18241 15335 18275
rect 17509 18241 17543 18275
rect 18429 18241 18463 18275
rect 19533 18241 19567 18275
rect 21281 18241 21315 18275
rect 22036 18241 22070 18275
rect 22290 18241 22324 18275
rect 23480 18241 23514 18275
rect 27077 18241 27111 18275
rect 29469 18241 29503 18275
rect 29617 18241 29651 18275
rect 29745 18241 29779 18275
rect 29975 18241 30009 18275
rect 31033 18241 31067 18275
rect 32689 18241 32723 18275
rect 33701 18241 33735 18275
rect 33849 18241 33883 18275
rect 33977 18241 34011 18275
rect 34166 18241 34200 18275
rect 35357 18241 35391 18275
rect 36369 18241 36403 18275
rect 36553 18241 36587 18275
rect 37565 18241 37599 18275
rect 46673 18241 46707 18275
rect 46857 18241 46891 18275
rect 47593 18241 47627 18275
rect 53573 18241 53607 18275
rect 7205 18173 7239 18207
rect 14381 18173 14415 18207
rect 14657 18173 14691 18207
rect 17417 18173 17451 18207
rect 17601 18173 17635 18207
rect 17693 18173 17727 18207
rect 18521 18173 18555 18207
rect 18613 18173 18647 18207
rect 18705 18173 18739 18207
rect 19441 18173 19475 18207
rect 19626 18173 19660 18207
rect 19717 18173 19751 18207
rect 23213 18173 23247 18207
rect 30757 18173 30791 18207
rect 32413 18173 32447 18207
rect 35725 18173 35759 18207
rect 36461 18173 36495 18207
rect 36645 18173 36679 18207
rect 37289 18173 37323 18207
rect 54033 18173 54067 18207
rect 6745 18105 6779 18139
rect 15485 18105 15519 18139
rect 18245 18105 18279 18139
rect 30113 18105 30147 18139
rect 3249 18037 3283 18071
rect 8585 18037 8619 18071
rect 21005 18037 21039 18071
rect 21833 18037 21867 18071
rect 24593 18037 24627 18071
rect 27445 18037 27479 18071
rect 27629 18037 27663 18071
rect 34345 18037 34379 18071
rect 35633 18037 35667 18071
rect 36185 18037 36219 18071
rect 43913 18037 43947 18071
rect 47041 18037 47075 18071
rect 48973 18037 49007 18071
rect 6377 17833 6411 17867
rect 33885 17833 33919 17867
rect 37657 17833 37691 17867
rect 43913 17833 43947 17867
rect 47041 17833 47075 17867
rect 47225 17833 47259 17867
rect 22109 17765 22143 17799
rect 24409 17765 24443 17799
rect 6837 17697 6871 17731
rect 6929 17697 6963 17731
rect 8953 17697 8987 17731
rect 16313 17697 16347 17731
rect 17509 17697 17543 17731
rect 31125 17697 31159 17731
rect 31401 17697 31435 17731
rect 37197 17697 37231 17731
rect 37841 17697 37875 17731
rect 37933 17697 37967 17731
rect 44189 17697 44223 17731
rect 44281 17697 44315 17731
rect 1409 17629 1443 17663
rect 2145 17629 2179 17663
rect 3801 17629 3835 17663
rect 14565 17629 14599 17663
rect 16037 17629 16071 17663
rect 17233 17629 17267 17663
rect 20729 17629 20763 17663
rect 20996 17629 21030 17663
rect 24593 17629 24627 17663
rect 24869 17629 24903 17663
rect 25513 17629 25547 17663
rect 26157 17629 26191 17663
rect 29561 17629 29595 17663
rect 29654 17629 29688 17663
rect 30026 17629 30060 17663
rect 33241 17629 33275 17663
rect 33389 17629 33423 17663
rect 33747 17629 33781 17663
rect 36737 17629 36771 17663
rect 36829 17629 36863 17663
rect 38025 17629 38059 17663
rect 38117 17629 38151 17663
rect 40785 17629 40819 17663
rect 42625 17629 42659 17663
rect 42809 17629 42843 17663
rect 43085 17629 43119 17663
rect 44097 17629 44131 17663
rect 44373 17629 44407 17663
rect 47685 17629 47719 17663
rect 47869 17629 47903 17663
rect 4046 17561 4080 17595
rect 5733 17561 5767 17595
rect 9198 17561 9232 17595
rect 25329 17561 25363 17595
rect 26402 17561 26436 17595
rect 29837 17561 29871 17595
rect 29929 17561 29963 17595
rect 33517 17561 33551 17595
rect 33609 17561 33643 17595
rect 37105 17561 37139 17595
rect 41052 17561 41086 17595
rect 46857 17561 46891 17595
rect 47073 17561 47107 17595
rect 47777 17561 47811 17595
rect 1593 17493 1627 17527
rect 2329 17493 2363 17527
rect 5181 17493 5215 17527
rect 5825 17493 5859 17527
rect 6745 17493 6779 17527
rect 10333 17493 10367 17527
rect 14841 17493 14875 17527
rect 24777 17493 24811 17527
rect 25697 17493 25731 17527
rect 27537 17493 27571 17527
rect 30205 17493 30239 17527
rect 36553 17493 36587 17527
rect 37013 17493 37047 17527
rect 42165 17493 42199 17527
rect 42993 17493 43027 17527
rect 3801 17289 3835 17323
rect 4169 17289 4203 17323
rect 7021 17289 7055 17323
rect 7849 17289 7883 17323
rect 13185 17289 13219 17323
rect 16681 17289 16715 17323
rect 18705 17289 18739 17323
rect 36569 17289 36603 17323
rect 42533 17289 42567 17323
rect 44189 17289 44223 17323
rect 12817 17221 12851 17255
rect 13001 17221 13035 17255
rect 33517 17221 33551 17255
rect 33609 17221 33643 17255
rect 36369 17221 36403 17255
rect 44097 17221 44131 17255
rect 44281 17221 44315 17255
rect 1869 17153 1903 17187
rect 2881 17153 2915 17187
rect 3985 17153 4019 17187
rect 4261 17153 4295 17187
rect 8033 17153 8067 17187
rect 16865 17153 16899 17187
rect 17141 17153 17175 17187
rect 18061 17153 18095 17187
rect 18981 17153 19015 17187
rect 19073 17153 19107 17187
rect 26157 17153 26191 17187
rect 29193 17153 29227 17187
rect 29286 17153 29320 17187
rect 29469 17153 29503 17187
rect 29561 17153 29595 17187
rect 29699 17153 29733 17187
rect 32137 17153 32171 17187
rect 33241 17153 33275 17187
rect 33334 17153 33368 17187
rect 33747 17153 33781 17187
rect 42441 17153 42475 17187
rect 44373 17153 44407 17187
rect 51457 17153 51491 17187
rect 7113 17085 7147 17119
rect 7205 17085 7239 17119
rect 13737 17085 13771 17119
rect 14013 17085 14047 17119
rect 15025 17085 15059 17119
rect 15301 17085 15335 17119
rect 16957 17085 16991 17119
rect 17049 17085 17083 17119
rect 17877 17085 17911 17119
rect 17969 17085 18003 17119
rect 18153 17085 18187 17119
rect 18889 17085 18923 17119
rect 19165 17085 19199 17119
rect 30297 17085 30331 17119
rect 30573 17085 30607 17119
rect 2697 17017 2731 17051
rect 6653 17017 6687 17051
rect 33885 17017 33919 17051
rect 2145 16949 2179 16983
rect 13001 16949 13035 16983
rect 17693 16949 17727 16983
rect 25973 16949 26007 16983
rect 29837 16949 29871 16983
rect 32321 16949 32355 16983
rect 36553 16949 36587 16983
rect 36737 16949 36771 16983
rect 51273 16949 51307 16983
rect 14381 16745 14415 16779
rect 24593 16745 24627 16779
rect 25145 16745 25179 16779
rect 29009 16745 29043 16779
rect 31677 16745 31711 16779
rect 46121 16745 46155 16779
rect 46949 16745 46983 16779
rect 28457 16677 28491 16711
rect 40693 16677 40727 16711
rect 45109 16677 45143 16711
rect 46581 16677 46615 16711
rect 1593 16609 1627 16643
rect 12173 16609 12207 16643
rect 16129 16609 16163 16643
rect 16865 16609 16899 16643
rect 16957 16609 16991 16643
rect 17141 16609 17175 16643
rect 17693 16609 17727 16643
rect 17969 16609 18003 16643
rect 20269 16609 20303 16643
rect 37565 16609 37599 16643
rect 42533 16609 42567 16643
rect 47869 16609 47903 16643
rect 50813 16609 50847 16643
rect 53389 16609 53423 16643
rect 6929 16541 6963 16575
rect 10977 16541 11011 16575
rect 17049 16541 17083 16575
rect 28733 16541 28767 16575
rect 28825 16541 28859 16575
rect 29745 16541 29779 16575
rect 30021 16541 30055 16575
rect 31033 16541 31067 16575
rect 31181 16541 31215 16575
rect 31309 16541 31343 16575
rect 31498 16541 31532 16575
rect 35173 16541 35207 16575
rect 35265 16541 35299 16575
rect 36047 16541 36081 16575
rect 36182 16541 36216 16575
rect 24639 16507 24673 16541
rect 36277 16538 36311 16572
rect 36461 16541 36495 16575
rect 37105 16541 37139 16575
rect 40877 16541 40911 16575
rect 41153 16541 41187 16575
rect 41337 16541 41371 16575
rect 41797 16541 41831 16575
rect 41981 16541 42015 16575
rect 42257 16541 42291 16575
rect 42625 16541 42659 16575
rect 45293 16541 45327 16575
rect 45845 16541 45879 16575
rect 45937 16541 45971 16575
rect 51080 16541 51114 16575
rect 1860 16473 1894 16507
rect 12440 16473 12474 16507
rect 14197 16473 14231 16507
rect 15209 16473 15243 16507
rect 15393 16473 15427 16507
rect 15945 16473 15979 16507
rect 20536 16473 20570 16507
rect 24409 16473 24443 16507
rect 25697 16473 25731 16507
rect 28641 16473 28675 16507
rect 31401 16473 31435 16507
rect 37810 16473 37844 16507
rect 45017 16473 45051 16507
rect 45201 16473 45235 16507
rect 48114 16473 48148 16507
rect 53634 16473 53668 16507
rect 2973 16405 3007 16439
rect 6745 16405 6779 16439
rect 11069 16405 11103 16439
rect 13553 16405 13587 16439
rect 14381 16405 14415 16439
rect 14565 16405 14599 16439
rect 16681 16405 16715 16439
rect 21649 16405 21683 16439
rect 24777 16405 24811 16439
rect 25789 16405 25823 16439
rect 35817 16405 35851 16439
rect 36921 16405 36955 16439
rect 38945 16405 38979 16439
rect 42809 16405 42843 16439
rect 46949 16405 46983 16439
rect 47133 16405 47167 16439
rect 49249 16405 49283 16439
rect 52193 16405 52227 16439
rect 54769 16405 54803 16439
rect 2329 16201 2363 16235
rect 2697 16201 2731 16235
rect 12357 16201 12391 16235
rect 17969 16201 18003 16235
rect 21833 16201 21867 16235
rect 22201 16201 22235 16235
rect 28181 16201 28215 16235
rect 36737 16201 36771 16235
rect 40601 16201 40635 16235
rect 46765 16201 46799 16235
rect 47685 16201 47719 16235
rect 51733 16201 51767 16235
rect 1869 16133 1903 16167
rect 30021 16133 30055 16167
rect 35624 16133 35658 16167
rect 46581 16133 46615 16167
rect 51365 16133 51399 16167
rect 51581 16133 51615 16167
rect 53205 16133 53239 16167
rect 54217 16133 54251 16167
rect 1501 16065 1535 16099
rect 2513 16065 2547 16099
rect 2789 16065 2823 16099
rect 4537 16065 4571 16099
rect 7001 16065 7035 16099
rect 9597 16065 9631 16099
rect 9864 16065 9898 16099
rect 11713 16065 11747 16099
rect 12541 16065 12575 16099
rect 15945 16065 15979 16099
rect 16957 16065 16991 16099
rect 18153 16065 18187 16099
rect 18245 16065 18279 16099
rect 18429 16065 18463 16099
rect 22017 16065 22051 16099
rect 22293 16065 22327 16099
rect 23213 16065 23247 16099
rect 23480 16065 23514 16099
rect 28365 16065 28399 16099
rect 28549 16065 28583 16099
rect 28641 16065 28675 16099
rect 29653 16065 29687 16099
rect 29801 16065 29835 16099
rect 29929 16065 29963 16099
rect 30118 16065 30152 16099
rect 32597 16065 32631 16099
rect 32864 16065 32898 16099
rect 35357 16065 35391 16099
rect 40325 16065 40359 16099
rect 40417 16065 40451 16099
rect 43637 16065 43671 16099
rect 46397 16065 46431 16099
rect 47869 16065 47903 16099
rect 53389 16065 53423 16099
rect 53481 16065 53515 16099
rect 53941 16065 53975 16099
rect 6745 15997 6779 16031
rect 11529 15997 11563 16031
rect 16681 15997 16715 16031
rect 18337 15997 18371 16031
rect 28457 15997 28491 16031
rect 54217 15997 54251 16031
rect 53205 15929 53239 15963
rect 4353 15861 4387 15895
rect 8125 15861 8159 15895
rect 10977 15861 11011 15895
rect 11897 15861 11931 15895
rect 16037 15861 16071 15895
rect 24593 15861 24627 15895
rect 30297 15861 30331 15895
rect 33977 15861 34011 15895
rect 43729 15861 43763 15895
rect 51549 15861 51583 15895
rect 54033 15861 54067 15895
rect 23029 15657 23063 15691
rect 23581 15657 23615 15691
rect 23765 15657 23799 15691
rect 24409 15657 24443 15691
rect 43177 15657 43211 15691
rect 43913 15657 43947 15691
rect 52285 15657 52319 15691
rect 52929 15657 52963 15691
rect 6561 15589 6595 15623
rect 10609 15589 10643 15623
rect 11897 15589 11931 15623
rect 17417 15589 17451 15623
rect 7113 15521 7147 15555
rect 16405 15521 16439 15555
rect 17693 15521 17727 15555
rect 25973 15521 26007 15555
rect 32689 15521 32723 15555
rect 42533 15521 42567 15555
rect 43018 15521 43052 15555
rect 53205 15521 53239 15555
rect 1409 15453 1443 15487
rect 2329 15453 2363 15487
rect 4077 15453 4111 15487
rect 4344 15453 4378 15487
rect 10793 15453 10827 15487
rect 10885 15453 10919 15487
rect 11069 15453 11103 15487
rect 11161 15453 11195 15487
rect 13185 15453 13219 15487
rect 13369 15453 13403 15487
rect 16129 15453 16163 15487
rect 17601 15453 17635 15487
rect 17785 15453 17819 15487
rect 17877 15453 17911 15487
rect 20177 15453 20211 15487
rect 24593 15453 24627 15487
rect 24869 15453 24903 15487
rect 29653 15453 29687 15487
rect 29745 15453 29779 15487
rect 32781 15453 32815 15487
rect 42809 15453 42843 15487
rect 43729 15453 43763 15487
rect 44005 15453 44039 15487
rect 48053 15453 48087 15487
rect 52193 15453 52227 15487
rect 52469 15453 52503 15487
rect 53113 15453 53147 15487
rect 53297 15453 53331 15487
rect 53389 15453 53423 15487
rect 53941 15453 53975 15487
rect 55689 15453 55723 15487
rect 55873 15453 55907 15487
rect 7021 15385 7055 15419
rect 11713 15385 11747 15419
rect 20444 15385 20478 15419
rect 23397 15385 23431 15419
rect 23581 15385 23615 15419
rect 26240 15385 26274 15419
rect 43637 15385 43671 15419
rect 44097 15385 44131 15419
rect 52377 15385 52411 15419
rect 1593 15317 1627 15351
rect 2145 15317 2179 15351
rect 5457 15317 5491 15351
rect 6929 15317 6963 15351
rect 13277 15317 13311 15351
rect 21557 15317 21591 15351
rect 24777 15317 24811 15351
rect 27353 15317 27387 15351
rect 29929 15317 29963 15351
rect 33149 15317 33183 15351
rect 42901 15317 42935 15351
rect 47869 15317 47903 15351
rect 54171 15317 54205 15351
rect 55781 15317 55815 15351
rect 4537 15113 4571 15147
rect 11529 15113 11563 15147
rect 12725 15113 12759 15147
rect 17877 15113 17911 15147
rect 21833 15113 21867 15147
rect 23489 15113 23523 15147
rect 23949 15113 23983 15147
rect 24685 15113 24719 15147
rect 25881 15113 25915 15147
rect 29193 15113 29227 15147
rect 30941 15113 30975 15147
rect 32873 15113 32907 15147
rect 41613 15113 41647 15147
rect 45017 15113 45051 15147
rect 57345 15113 57379 15147
rect 13185 15045 13219 15079
rect 22201 15045 22235 15079
rect 23029 15045 23063 15079
rect 24317 15045 24351 15079
rect 33517 15045 33551 15079
rect 39037 15045 39071 15079
rect 39129 15045 39163 15079
rect 40969 15045 41003 15079
rect 43904 15045 43938 15079
rect 47860 15045 47894 15079
rect 50261 15045 50295 15079
rect 55413 15045 55447 15079
rect 56210 15045 56244 15079
rect 24547 15011 24581 15045
rect 1409 14977 1443 15011
rect 2329 14977 2363 15011
rect 4905 14977 4939 15011
rect 7573 14977 7607 15011
rect 7665 14977 7699 15011
rect 7849 14977 7883 15011
rect 7941 14977 7975 15011
rect 11897 14977 11931 15011
rect 13093 14977 13127 15011
rect 17325 14977 17359 15011
rect 18061 14977 18095 15011
rect 18153 14977 18187 15011
rect 18245 14977 18279 15011
rect 22017 14977 22051 15011
rect 22293 14977 22327 15011
rect 22845 14977 22879 15011
rect 23673 14977 23707 15011
rect 26341 14977 26375 15011
rect 26985 14977 27019 15011
rect 27169 14977 27203 15011
rect 29009 14977 29043 15011
rect 29285 14977 29319 15011
rect 29929 14977 29963 15011
rect 30113 14977 30147 15011
rect 30757 14977 30791 15011
rect 30941 14977 30975 15011
rect 33149 14977 33183 15011
rect 33425 14977 33459 15011
rect 38761 14977 38795 15011
rect 40601 14977 40635 15011
rect 40785 14977 40819 15011
rect 41429 14977 41463 15011
rect 41613 14977 41647 15011
rect 51089 14977 51123 15011
rect 52929 14977 52963 15011
rect 53021 14977 53055 15011
rect 55229 14977 55263 15011
rect 4997 14909 5031 14943
rect 5181 14909 5215 14943
rect 11989 14909 12023 14943
rect 12081 14909 12115 14943
rect 13277 14909 13311 14943
rect 17049 14909 17083 14943
rect 17141 14909 17175 14943
rect 17233 14909 17267 14943
rect 18337 14909 18371 14943
rect 26065 14909 26099 14943
rect 26157 14909 26191 14943
rect 26249 14909 26283 14943
rect 30021 14909 30055 14943
rect 30205 14909 30239 14943
rect 33057 14909 33091 14943
rect 38669 14909 38703 14943
rect 43637 14909 43671 14943
rect 47593 14909 47627 14943
rect 52745 14909 52779 14943
rect 53113 14909 53147 14943
rect 53205 14909 53239 14943
rect 55045 14909 55079 14943
rect 55965 14909 55999 14943
rect 2145 14841 2179 14875
rect 16865 14841 16899 14875
rect 27077 14841 27111 14875
rect 28825 14841 28859 14875
rect 49893 14841 49927 14875
rect 50445 14841 50479 14875
rect 1593 14773 1627 14807
rect 7389 14773 7423 14807
rect 24501 14773 24535 14807
rect 29745 14773 29779 14807
rect 38485 14773 38519 14807
rect 48973 14773 49007 14807
rect 50261 14773 50295 14807
rect 50905 14773 50939 14807
rect 2973 14569 3007 14603
rect 8033 14569 8067 14603
rect 14105 14569 14139 14603
rect 14473 14569 14507 14603
rect 17325 14569 17359 14603
rect 26341 14569 26375 14603
rect 28411 14569 28445 14603
rect 30941 14569 30975 14603
rect 47593 14569 47627 14603
rect 47777 14569 47811 14603
rect 52193 14569 52227 14603
rect 55413 14569 55447 14603
rect 55505 14569 55539 14603
rect 35541 14501 35575 14535
rect 36829 14501 36863 14535
rect 41705 14501 41739 14535
rect 48605 14501 48639 14535
rect 7941 14433 7975 14467
rect 16589 14433 16623 14467
rect 17601 14433 17635 14467
rect 17785 14433 17819 14467
rect 37933 14433 37967 14467
rect 42717 14433 42751 14467
rect 50813 14433 50847 14467
rect 55597 14433 55631 14467
rect 1593 14365 1627 14399
rect 6837 14365 6871 14399
rect 7113 14365 7147 14399
rect 8033 14365 8067 14399
rect 8953 14365 8987 14399
rect 9137 14365 9171 14399
rect 14289 14365 14323 14399
rect 14565 14365 14599 14399
rect 16497 14365 16531 14399
rect 16681 14365 16715 14399
rect 16773 14365 16807 14399
rect 17509 14365 17543 14399
rect 17694 14365 17728 14399
rect 25973 14365 26007 14399
rect 28181 14365 28215 14399
rect 29561 14365 29595 14399
rect 29828 14365 29862 14399
rect 38200 14365 38234 14399
rect 41705 14365 41739 14399
rect 41981 14365 42015 14399
rect 48237 14365 48271 14399
rect 49065 14365 49099 14399
rect 49249 14365 49283 14399
rect 51069 14365 51103 14399
rect 55321 14365 55355 14399
rect 1860 14297 1894 14331
rect 7573 14297 7607 14331
rect 26157 14297 26191 14331
rect 35357 14297 35391 14331
rect 36553 14297 36587 14331
rect 42533 14297 42567 14331
rect 47409 14297 47443 14331
rect 48421 14297 48455 14331
rect 6653 14229 6687 14263
rect 7021 14229 7055 14263
rect 8217 14229 8251 14263
rect 9321 14229 9355 14263
rect 16313 14229 16347 14263
rect 39313 14229 39347 14263
rect 41889 14229 41923 14263
rect 47619 14229 47653 14263
rect 49157 14229 49191 14263
rect 2329 14025 2363 14059
rect 2697 14025 2731 14059
rect 14473 14025 14507 14059
rect 17693 14025 17727 14059
rect 20821 14025 20855 14059
rect 23305 14025 23339 14059
rect 23791 14025 23825 14059
rect 24609 14025 24643 14059
rect 26065 14025 26099 14059
rect 35541 14025 35575 14059
rect 36461 14025 36495 14059
rect 37841 14025 37875 14059
rect 53113 14025 53147 14059
rect 54033 14025 54067 14059
rect 54217 14025 54251 14059
rect 7757 13957 7791 13991
rect 9781 13957 9815 13991
rect 14105 13957 14139 13991
rect 14305 13957 14339 13991
rect 23581 13957 23615 13991
rect 24409 13957 24443 13991
rect 37749 13957 37783 13991
rect 52745 13957 52779 13991
rect 53849 13957 53883 13991
rect 1409 13889 1443 13923
rect 2513 13889 2547 13923
rect 2789 13889 2823 13923
rect 10793 13889 10827 13923
rect 16957 13889 16991 13923
rect 17049 13889 17083 13923
rect 17877 13889 17911 13923
rect 18061 13889 18095 13923
rect 19441 13889 19475 13923
rect 19708 13889 19742 13923
rect 25697 13889 25731 13923
rect 33241 13889 33275 13923
rect 33497 13889 33531 13923
rect 35357 13889 35391 13923
rect 36277 13889 36311 13923
rect 38577 13889 38611 13923
rect 38761 13889 38795 13923
rect 40417 13889 40451 13923
rect 42881 13889 42915 13923
rect 45661 13889 45695 13923
rect 45845 13889 45879 13923
rect 47777 13889 47811 13923
rect 52929 13889 52963 13923
rect 53021 13889 53055 13923
rect 54125 13889 54159 13923
rect 8125 13821 8159 13855
rect 8493 13821 8527 13855
rect 10609 13821 10643 13855
rect 10977 13821 11011 13855
rect 16681 13821 16715 13855
rect 16865 13821 16899 13855
rect 17141 13821 17175 13855
rect 17969 13821 18003 13855
rect 18153 13821 18187 13855
rect 36093 13821 36127 13855
rect 38669 13821 38703 13855
rect 40693 13821 40727 13855
rect 42625 13821 42659 13855
rect 47869 13821 47903 13855
rect 8033 13753 8067 13787
rect 9965 13753 9999 13787
rect 23949 13753 23983 13787
rect 24777 13753 24811 13787
rect 34621 13753 34655 13787
rect 48145 13753 48179 13787
rect 1593 13685 1627 13719
rect 7922 13685 7956 13719
rect 14289 13685 14323 13719
rect 23765 13685 23799 13719
rect 24593 13685 24627 13719
rect 26065 13685 26099 13719
rect 26249 13685 26283 13719
rect 44005 13685 44039 13719
rect 46029 13685 46063 13719
rect 53297 13685 53331 13719
rect 54401 13685 54435 13719
rect 6929 13481 6963 13515
rect 7205 13481 7239 13515
rect 10241 13481 10275 13515
rect 19993 13481 20027 13515
rect 22109 13481 22143 13515
rect 23121 13481 23155 13515
rect 23581 13481 23615 13515
rect 30573 13481 30607 13515
rect 33333 13481 33367 13515
rect 36553 13481 36587 13515
rect 37289 13481 37323 13515
rect 41429 13481 41463 13515
rect 42809 13481 42843 13515
rect 51181 13481 51215 13515
rect 54585 13481 54619 13515
rect 55689 13481 55723 13515
rect 57713 13481 57747 13515
rect 7389 13413 7423 13447
rect 8217 13413 8251 13447
rect 23765 13413 23799 13447
rect 51365 13413 51399 13447
rect 54769 13413 54803 13447
rect 3801 13345 3835 13379
rect 10241 13345 10275 13379
rect 11437 13345 11471 13379
rect 25145 13345 25179 13379
rect 28365 13345 28399 13379
rect 33977 13345 34011 13379
rect 46029 13345 46063 13379
rect 55321 13345 55355 13379
rect 1409 13277 1443 13311
rect 2329 13277 2363 13311
rect 7297 13277 7331 13311
rect 7665 13277 7699 13311
rect 8125 13277 8159 13311
rect 8309 13277 8343 13311
rect 10149 13277 10183 13311
rect 11713 13277 11747 13311
rect 14105 13277 14139 13311
rect 20177 13277 20211 13311
rect 20453 13277 20487 13311
rect 21281 13277 21315 13311
rect 21925 13277 21959 13311
rect 22477 13277 22511 13311
rect 24869 13277 24903 13311
rect 25789 13277 25823 13311
rect 26157 13277 26191 13311
rect 26801 13277 26835 13311
rect 28273 13277 28307 13311
rect 28457 13277 28491 13311
rect 30389 13277 30423 13311
rect 31861 13277 31895 13311
rect 33517 13277 33551 13311
rect 33609 13277 33643 13311
rect 36369 13277 36403 13311
rect 37105 13277 37139 13311
rect 38761 13277 38795 13311
rect 39037 13277 39071 13311
rect 41245 13277 41279 13311
rect 42441 13277 42475 13311
rect 42809 13277 42843 13311
rect 48513 13277 48547 13311
rect 50813 13277 50847 13311
rect 52009 13277 52043 13311
rect 53297 13277 53331 13311
rect 53481 13277 53515 13311
rect 56333 13277 56367 13311
rect 4068 13209 4102 13243
rect 14350 13209 14384 13243
rect 21097 13209 21131 13243
rect 23397 13209 23431 13243
rect 23613 13209 23647 13243
rect 25973 13209 26007 13243
rect 33885 13209 33919 13243
rect 41061 13209 41095 13243
rect 46274 13209 46308 13243
rect 53389 13209 53423 13243
rect 54401 13209 54435 13243
rect 55689 13209 55723 13243
rect 56578 13209 56612 13243
rect 1593 13141 1627 13175
rect 2145 13141 2179 13175
rect 5181 13141 5215 13175
rect 7573 13141 7607 13175
rect 10517 13141 10551 13175
rect 15485 13141 15519 13175
rect 20361 13141 20395 13175
rect 22661 13141 22695 13175
rect 26617 13141 26651 13175
rect 31677 13141 31711 13175
rect 38577 13141 38611 13175
rect 38945 13141 38979 13175
rect 42625 13141 42659 13175
rect 47409 13141 47443 13175
rect 48605 13141 48639 13175
rect 51181 13141 51215 13175
rect 51825 13141 51859 13175
rect 54601 13141 54635 13175
rect 55873 13141 55907 13175
rect 4077 12937 4111 12971
rect 4445 12937 4479 12971
rect 14197 12937 14231 12971
rect 14565 12937 14599 12971
rect 24133 12937 24167 12971
rect 25421 12937 25455 12971
rect 46029 12937 46063 12971
rect 48789 12937 48823 12971
rect 52193 12937 52227 12971
rect 55045 12937 55079 12971
rect 56057 12937 56091 12971
rect 2237 12869 2271 12903
rect 19349 12869 19383 12903
rect 30665 12869 30699 12903
rect 30865 12869 30899 12903
rect 32382 12869 32416 12903
rect 35817 12869 35851 12903
rect 38384 12869 38418 12903
rect 40693 12869 40727 12903
rect 41797 12869 41831 12903
rect 42809 12869 42843 12903
rect 51080 12869 51114 12903
rect 55413 12869 55447 12903
rect 1869 12801 1903 12835
rect 2697 12801 2731 12835
rect 3617 12801 3651 12835
rect 4261 12801 4295 12835
rect 4537 12801 4571 12835
rect 7205 12801 7239 12835
rect 7481 12801 7515 12835
rect 8217 12801 8251 12835
rect 8401 12801 8435 12835
rect 10425 12801 10459 12835
rect 10609 12801 10643 12835
rect 11529 12801 11563 12835
rect 11805 12801 11839 12835
rect 14381 12801 14415 12835
rect 14657 12801 14691 12835
rect 17141 12801 17175 12835
rect 17408 12801 17442 12835
rect 18981 12801 19015 12835
rect 19165 12801 19199 12835
rect 19441 12801 19475 12835
rect 21925 12801 21959 12835
rect 24041 12801 24075 12835
rect 24777 12801 24811 12835
rect 25605 12801 25639 12835
rect 32137 12801 32171 12835
rect 35633 12801 35667 12835
rect 38117 12801 38151 12835
rect 40601 12801 40635 12835
rect 40785 12801 40819 12835
rect 41705 12801 41739 12835
rect 42625 12801 42659 12835
rect 43453 12801 43487 12835
rect 46213 12801 46247 12835
rect 48697 12801 48731 12835
rect 48881 12801 48915 12835
rect 50813 12801 50847 12835
rect 55229 12801 55263 12835
rect 55505 12801 55539 12835
rect 56241 12801 56275 12835
rect 7297 12733 7331 12767
rect 11621 12733 11655 12767
rect 22661 12733 22695 12767
rect 22937 12733 22971 12767
rect 35449 12733 35483 12767
rect 43545 12733 43579 12767
rect 43729 12733 43763 12767
rect 7665 12665 7699 12699
rect 18521 12665 18555 12699
rect 22109 12665 22143 12699
rect 31033 12665 31067 12699
rect 42993 12665 43027 12699
rect 2881 12597 2915 12631
rect 3433 12597 3467 12631
rect 7481 12597 7515 12631
rect 8585 12597 8619 12631
rect 10609 12597 10643 12631
rect 10793 12597 10827 12631
rect 11529 12597 11563 12631
rect 11989 12597 12023 12631
rect 24869 12597 24903 12631
rect 30849 12597 30883 12631
rect 33517 12597 33551 12631
rect 39497 12597 39531 12631
rect 43637 12597 43671 12631
rect 6653 12393 6687 12427
rect 6837 12393 6871 12427
rect 7389 12393 7423 12427
rect 14979 12393 15013 12427
rect 16221 12393 16255 12427
rect 16405 12393 16439 12427
rect 20821 12393 20855 12427
rect 21281 12393 21315 12427
rect 21741 12393 21775 12427
rect 21925 12393 21959 12427
rect 23121 12393 23155 12427
rect 24593 12393 24627 12427
rect 25605 12393 25639 12427
rect 30941 12393 30975 12427
rect 31861 12393 31895 12427
rect 39865 12393 39899 12427
rect 44097 12393 44131 12427
rect 48329 12393 48363 12427
rect 50629 12393 50663 12427
rect 51825 12393 51859 12427
rect 3249 12325 3283 12359
rect 21465 12325 21499 12359
rect 34989 12325 35023 12359
rect 38669 12325 38703 12359
rect 42257 12325 42291 12359
rect 48237 12325 48271 12359
rect 52009 12325 52043 12359
rect 6561 12257 6595 12291
rect 8953 12257 8987 12291
rect 9229 12257 9263 12291
rect 11713 12257 11747 12291
rect 17233 12257 17267 12291
rect 17509 12257 17543 12291
rect 26065 12257 26099 12291
rect 29561 12257 29595 12291
rect 48421 12257 48455 12291
rect 50813 12257 50847 12291
rect 50905 12257 50939 12291
rect 55597 12257 55631 12291
rect 1869 12189 1903 12223
rect 2136 12189 2170 12223
rect 6469 12189 6503 12223
rect 7297 12189 7331 12223
rect 7665 12189 7699 12223
rect 10241 12189 10275 12223
rect 10701 12189 10735 12223
rect 11069 12189 11103 12223
rect 11437 12189 11471 12223
rect 12633 12189 12667 12223
rect 12817 12189 12851 12223
rect 14749 12189 14783 12223
rect 21925 12189 21959 12223
rect 22109 12189 22143 12223
rect 23011 12189 23045 12223
rect 25237 12189 25271 12223
rect 28825 12189 28859 12223
rect 31493 12189 31527 12223
rect 31677 12189 31711 12223
rect 35265 12189 35299 12223
rect 36185 12189 36219 12223
rect 38567 12189 38601 12223
rect 38761 12189 38795 12223
rect 38853 12189 38887 12223
rect 39865 12189 39899 12223
rect 40049 12189 40083 12223
rect 43065 12189 43099 12223
rect 43174 12186 43208 12220
rect 43269 12189 43303 12223
rect 43453 12189 43487 12223
rect 44005 12189 44039 12223
rect 48145 12189 48179 12223
rect 48605 12189 48639 12223
rect 50997 12189 51031 12223
rect 51089 12189 51123 12223
rect 55321 12189 55355 12223
rect 55413 12189 55447 12223
rect 13001 12121 13035 12155
rect 16037 12121 16071 12155
rect 21097 12121 21131 12155
rect 21313 12121 21347 12155
rect 24409 12121 24443 12155
rect 24625 12121 24659 12155
rect 25421 12121 25455 12155
rect 26332 12121 26366 12155
rect 29806 12121 29840 12155
rect 34989 12121 35023 12155
rect 41889 12121 41923 12155
rect 51641 12121 51675 12155
rect 7849 12053 7883 12087
rect 16247 12053 16281 12087
rect 24777 12053 24811 12087
rect 27445 12053 27479 12087
rect 28641 12053 28675 12087
rect 35173 12053 35207 12087
rect 35909 12053 35943 12087
rect 38393 12053 38427 12087
rect 42349 12053 42383 12087
rect 42809 12053 42843 12087
rect 47869 12053 47903 12087
rect 51841 12053 51875 12087
rect 55597 12053 55631 12087
rect 2605 11849 2639 11883
rect 10977 11849 11011 11883
rect 46581 11849 46615 11883
rect 48053 11849 48087 11883
rect 56057 11849 56091 11883
rect 5641 11781 5675 11815
rect 7481 11781 7515 11815
rect 10793 11781 10827 11815
rect 15577 11781 15611 11815
rect 24133 11781 24167 11815
rect 28457 11781 28491 11815
rect 42901 11781 42935 11815
rect 45446 11781 45480 11815
rect 53941 11781 53975 11815
rect 54125 11781 54159 11815
rect 1409 11713 1443 11747
rect 2513 11713 2547 11747
rect 3525 11713 3559 11747
rect 8677 11713 8711 11747
rect 10609 11713 10643 11747
rect 12173 11713 12207 11747
rect 13001 11713 13035 11747
rect 13185 11713 13219 11747
rect 14841 11713 14875 11747
rect 15485 11713 15519 11747
rect 17141 11713 17175 11747
rect 18981 11713 19015 11747
rect 19165 11713 19199 11747
rect 19257 11713 19291 11747
rect 22109 11713 22143 11747
rect 22293 11713 22327 11747
rect 23949 11713 23983 11747
rect 28089 11713 28123 11747
rect 29377 11713 29411 11747
rect 32505 11713 32539 11747
rect 34529 11713 34563 11747
rect 34796 11713 34830 11747
rect 36369 11713 36403 11747
rect 36461 11713 36495 11747
rect 42717 11713 42751 11747
rect 43617 11713 43651 11747
rect 45201 11713 45235 11747
rect 47961 11713 47995 11747
rect 49065 11713 49099 11747
rect 51457 11713 51491 11747
rect 54217 11713 54251 11747
rect 54933 11713 54967 11747
rect 2697 11645 2731 11679
rect 8401 11645 8435 11679
rect 15669 11645 15703 11679
rect 16865 11645 16899 11679
rect 22017 11645 22051 11679
rect 22201 11645 22235 11679
rect 29285 11645 29319 11679
rect 29469 11645 29503 11679
rect 29561 11645 29595 11679
rect 36645 11645 36679 11679
rect 43361 11645 43395 11679
rect 51549 11645 51583 11679
rect 51733 11645 51767 11679
rect 54677 11645 54711 11679
rect 2145 11577 2179 11611
rect 13093 11577 13127 11611
rect 15117 11577 15151 11611
rect 29101 11577 29135 11611
rect 32689 11577 32723 11611
rect 35909 11577 35943 11611
rect 51641 11577 51675 11611
rect 53941 11577 53975 11611
rect 1593 11509 1627 11543
rect 3341 11509 3375 11543
rect 5733 11509 5767 11543
rect 7573 11509 7607 11543
rect 18797 11509 18831 11543
rect 21833 11509 21867 11543
rect 24317 11509 24351 11543
rect 28457 11509 28491 11543
rect 28641 11509 28675 11543
rect 36553 11509 36587 11543
rect 44741 11509 44775 11543
rect 48697 11509 48731 11543
rect 5457 11305 5491 11339
rect 9505 11305 9539 11339
rect 12909 11305 12943 11339
rect 14105 11305 14139 11339
rect 17601 11305 17635 11339
rect 21557 11305 21591 11339
rect 23397 11305 23431 11339
rect 23581 11305 23615 11339
rect 34805 11305 34839 11339
rect 36093 11305 36127 11339
rect 36185 11305 36219 11339
rect 43269 11305 43303 11339
rect 47777 11305 47811 11339
rect 12357 11237 12391 11271
rect 13369 11237 13403 11271
rect 23029 11237 23063 11271
rect 35265 11237 35299 11271
rect 40785 11237 40819 11271
rect 48605 11237 48639 11271
rect 51365 11237 51399 11271
rect 4077 11169 4111 11203
rect 13093 11169 13127 11203
rect 16313 11169 16347 11203
rect 16589 11169 16623 11203
rect 18061 11169 18095 11203
rect 42901 11169 42935 11203
rect 2697 11101 2731 11135
rect 10057 11101 10091 11135
rect 10241 11101 10275 11135
rect 12173 11101 12207 11135
rect 13185 11101 13219 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 17785 11101 17819 11135
rect 17877 11101 17911 11135
rect 17969 11101 18003 11135
rect 22201 11101 22235 11135
rect 22477 11101 22511 11135
rect 24777 11101 24811 11135
rect 28181 11101 28215 11135
rect 29837 11101 29871 11135
rect 30113 11101 30147 11135
rect 34713 11101 34747 11135
rect 35081 11101 35115 11135
rect 35714 11093 35748 11127
rect 36185 11101 36219 11135
rect 36737 11101 36771 11135
rect 36921 11101 36955 11135
rect 40969 11101 41003 11135
rect 41061 11101 41095 11135
rect 42533 11101 42567 11135
rect 42717 11101 42751 11135
rect 42809 11101 42843 11135
rect 43085 11101 43119 11135
rect 47685 11101 47719 11135
rect 48421 11101 48455 11135
rect 48513 11101 48547 11135
rect 51365 11101 51399 11135
rect 51641 11101 51675 11135
rect 1869 11033 1903 11067
rect 2053 11033 2087 11067
rect 4344 11033 4378 11067
rect 9413 11033 9447 11067
rect 12909 11033 12943 11067
rect 21189 11033 21223 11067
rect 21373 11033 21407 11067
rect 22017 11033 22051 11067
rect 23397 11033 23431 11067
rect 25022 11033 25056 11067
rect 28365 11033 28399 11067
rect 28549 11033 28583 11067
rect 29561 11033 29595 11067
rect 29929 11033 29963 11067
rect 35817 11033 35851 11067
rect 40785 11033 40819 11067
rect 2513 10965 2547 10999
rect 10149 10965 10183 10999
rect 22385 10965 22419 10999
rect 26157 10965 26191 10999
rect 29745 10965 29779 10999
rect 35935 10965 35969 10999
rect 36829 10965 36863 10999
rect 51549 10965 51583 10999
rect 4905 10761 4939 10795
rect 5273 10761 5307 10795
rect 13001 10761 13035 10795
rect 15577 10761 15611 10795
rect 19533 10761 19567 10795
rect 21281 10761 21315 10795
rect 22493 10761 22527 10795
rect 22661 10761 22695 10795
rect 24685 10761 24719 10795
rect 40325 10761 40359 10795
rect 40417 10761 40451 10795
rect 49341 10761 49375 10795
rect 2320 10693 2354 10727
rect 9496 10693 9530 10727
rect 18420 10693 18454 10727
rect 22293 10693 22327 10727
rect 38669 10693 38703 10727
rect 1593 10625 1627 10659
rect 2053 10625 2087 10659
rect 5089 10625 5123 10659
rect 5365 10625 5399 10659
rect 7205 10625 7239 10659
rect 7389 10625 7423 10659
rect 7481 10625 7515 10659
rect 12357 10625 12391 10659
rect 13001 10625 13035 10659
rect 13737 10625 13771 10659
rect 15853 10625 15887 10659
rect 16037 10625 16071 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 21097 10625 21131 10659
rect 21281 10625 21315 10659
rect 24869 10625 24903 10659
rect 27905 10625 27939 10659
rect 28089 10625 28123 10659
rect 31217 10625 31251 10659
rect 38485 10625 38519 10659
rect 39129 10625 39163 10659
rect 40233 10625 40267 10659
rect 40693 10625 40727 10659
rect 48217 10625 48251 10659
rect 7021 10557 7055 10591
rect 9229 10557 9263 10591
rect 11529 10557 11563 10591
rect 12081 10557 12115 10591
rect 12541 10557 12575 10591
rect 13093 10557 13127 10591
rect 13277 10557 13311 10591
rect 15761 10557 15795 10591
rect 15945 10557 15979 10591
rect 16957 10557 16991 10591
rect 17141 10557 17175 10591
rect 18153 10557 18187 10591
rect 31125 10557 31159 10591
rect 47961 10557 47995 10591
rect 7297 10489 7331 10523
rect 10609 10489 10643 10523
rect 1409 10421 1443 10455
rect 3433 10421 3467 10455
rect 13829 10421 13863 10455
rect 16681 10421 16715 10455
rect 22477 10421 22511 10455
rect 27997 10421 28031 10455
rect 31493 10421 31527 10455
rect 39405 10421 39439 10455
rect 39589 10421 39623 10455
rect 40601 10421 40635 10455
rect 40693 10421 40727 10455
rect 2145 10217 2179 10251
rect 6285 10217 6319 10251
rect 6469 10217 6503 10251
rect 7297 10217 7331 10251
rect 7757 10217 7791 10251
rect 10149 10217 10183 10251
rect 16865 10217 16899 10251
rect 39129 10217 39163 10251
rect 42625 10217 42659 10251
rect 47593 10217 47627 10251
rect 47961 10217 47995 10251
rect 52929 10217 52963 10251
rect 7389 10149 7423 10183
rect 22661 10149 22695 10183
rect 2697 10081 2731 10115
rect 6193 10081 6227 10115
rect 7481 10081 7515 10115
rect 17049 10081 17083 10115
rect 17325 10081 17359 10115
rect 27445 10081 27479 10115
rect 30665 10081 30699 10115
rect 46305 10081 46339 10115
rect 48053 10081 48087 10115
rect 51549 10081 51583 10115
rect 2513 10013 2547 10047
rect 2605 10013 2639 10047
rect 6009 10013 6043 10047
rect 6285 10013 6319 10047
rect 6929 10013 6963 10047
rect 9873 10013 9907 10047
rect 12265 10013 12299 10047
rect 12541 10013 12575 10047
rect 13093 10013 13127 10047
rect 13461 10013 13495 10047
rect 15669 10013 15703 10047
rect 17141 10013 17175 10047
rect 17233 10013 17267 10047
rect 22017 10013 22051 10047
rect 22110 10013 22144 10047
rect 22482 10013 22516 10047
rect 24777 10013 24811 10047
rect 24925 10013 24959 10047
rect 25053 10013 25087 10047
rect 25242 10013 25276 10047
rect 30941 10013 30975 10047
rect 36185 10013 36219 10047
rect 36369 10013 36403 10047
rect 37013 10013 37047 10047
rect 37657 10013 37691 10047
rect 37841 10013 37875 10047
rect 38853 10013 38887 10047
rect 41245 10013 41279 10047
rect 41501 10013 41535 10047
rect 46121 10013 46155 10047
rect 46397 10013 46431 10047
rect 47777 10013 47811 10047
rect 51805 10013 51839 10047
rect 13553 9945 13587 9979
rect 22293 9945 22327 9979
rect 22385 9945 22419 9979
rect 25145 9945 25179 9979
rect 27712 9945 27746 9979
rect 36829 9945 36863 9979
rect 37197 9945 37231 9979
rect 15761 9877 15795 9911
rect 25421 9877 25455 9911
rect 28825 9877 28859 9911
rect 32045 9877 32079 9911
rect 36277 9877 36311 9911
rect 37749 9877 37783 9911
rect 39313 9877 39347 9911
rect 45937 9877 45971 9911
rect 2605 9673 2639 9707
rect 15485 9673 15519 9707
rect 28089 9673 28123 9707
rect 30941 9673 30975 9707
rect 42441 9673 42475 9707
rect 2513 9605 2547 9639
rect 10057 9605 10091 9639
rect 15025 9605 15059 9639
rect 22078 9605 22112 9639
rect 28641 9605 28675 9639
rect 31493 9605 31527 9639
rect 35725 9605 35759 9639
rect 39037 9605 39071 9639
rect 42809 9605 42843 9639
rect 45928 9605 45962 9639
rect 49249 9605 49283 9639
rect 49465 9605 49499 9639
rect 1409 9537 1443 9571
rect 8309 9537 8343 9571
rect 9873 9537 9907 9571
rect 12449 9537 12483 9571
rect 13277 9537 13311 9571
rect 14841 9537 14875 9571
rect 15669 9537 15703 9571
rect 15761 9537 15795 9571
rect 18337 9537 18371 9571
rect 18604 9537 18638 9571
rect 25973 9537 26007 9571
rect 28365 9537 28399 9571
rect 31217 9537 31251 9571
rect 33589 9537 33623 9571
rect 36556 9537 36590 9571
rect 37289 9537 37323 9571
rect 38945 9537 38979 9571
rect 39129 9537 39163 9571
rect 39589 9537 39623 9571
rect 39773 9537 39807 9571
rect 42625 9537 42659 9571
rect 42717 9537 42751 9571
rect 42927 9537 42961 9571
rect 2697 9469 2731 9503
rect 6929 9469 6963 9503
rect 7481 9469 7515 9503
rect 7849 9469 7883 9503
rect 13185 9469 13219 9503
rect 15853 9469 15887 9503
rect 15945 9469 15979 9503
rect 21833 9469 21867 9503
rect 24685 9469 24719 9503
rect 24961 9469 24995 9503
rect 28273 9469 28307 9503
rect 28733 9469 28767 9503
rect 31126 9469 31160 9503
rect 31585 9469 31619 9503
rect 33333 9469 33367 9503
rect 36369 9469 36403 9503
rect 43085 9469 43119 9503
rect 45661 9469 45695 9503
rect 7297 9401 7331 9435
rect 7389 9401 7423 9435
rect 8493 9401 8527 9435
rect 19717 9401 19751 9435
rect 1593 9333 1627 9367
rect 2145 9333 2179 9367
rect 10241 9333 10275 9367
rect 13553 9333 13587 9367
rect 23213 9333 23247 9367
rect 26157 9333 26191 9367
rect 34713 9333 34747 9367
rect 35817 9333 35851 9367
rect 36737 9333 36771 9367
rect 37519 9333 37553 9367
rect 39589 9333 39623 9367
rect 47041 9333 47075 9367
rect 49433 9333 49467 9367
rect 49617 9333 49651 9367
rect 5917 9129 5951 9163
rect 8217 9129 8251 9163
rect 9321 9129 9355 9163
rect 10057 9129 10091 9163
rect 10333 9129 10367 9163
rect 13553 9129 13587 9163
rect 14316 9129 14350 9163
rect 19257 9129 19291 9163
rect 25421 9129 25455 9163
rect 33333 9129 33367 9163
rect 42165 9129 42199 9163
rect 46305 9129 46339 9163
rect 50997 9129 51031 9163
rect 21925 9061 21959 9095
rect 4537 8993 4571 9027
rect 15201 8993 15235 9027
rect 16037 8993 16071 9027
rect 16405 8993 16439 9027
rect 36737 8993 36771 9027
rect 36829 8993 36863 9027
rect 37473 8993 37507 9027
rect 51549 8993 51583 9027
rect 1593 8925 1627 8959
rect 2421 8925 2455 8959
rect 3065 8925 3099 8959
rect 8217 8925 8251 8959
rect 8401 8925 8435 8959
rect 9137 8925 9171 8959
rect 9873 8925 9907 8959
rect 12909 8925 12943 8959
rect 13057 8925 13091 8959
rect 13185 8925 13219 8959
rect 13415 8925 13449 8959
rect 15301 8925 15335 8959
rect 15394 8925 15428 8959
rect 15485 8925 15519 8959
rect 16221 8925 16255 8959
rect 16313 8925 16347 8959
rect 16497 8925 16531 8959
rect 19441 8925 19475 8959
rect 19717 8925 19751 8959
rect 22109 8925 22143 8959
rect 22845 8925 22879 8959
rect 23121 8925 23155 8959
rect 24777 8925 24811 8959
rect 24870 8925 24904 8959
rect 25053 8925 25087 8959
rect 25242 8925 25276 8959
rect 27997 8925 28031 8959
rect 28641 8925 28675 8959
rect 33517 8925 33551 8959
rect 33839 8925 33873 8959
rect 33977 8925 34011 8959
rect 36645 8925 36679 8959
rect 36921 8925 36955 8959
rect 37749 8925 37783 8959
rect 38853 8925 38887 8959
rect 39037 8925 39071 8959
rect 45201 8925 45235 8959
rect 45293 8925 45327 8959
rect 45661 8925 45695 8959
rect 48237 8925 48271 8959
rect 50813 8925 50847 8959
rect 51089 8925 51123 8959
rect 4804 8857 4838 8891
rect 8953 8857 8987 8891
rect 13277 8857 13311 8891
rect 14105 8857 14139 8891
rect 25145 8857 25179 8891
rect 33609 8857 33643 8891
rect 33701 8857 33735 8891
rect 41981 8857 42015 8891
rect 42197 8857 42231 8891
rect 45385 8857 45419 8891
rect 45503 8857 45537 8891
rect 46121 8857 46155 8891
rect 46337 8857 46371 8891
rect 48504 8857 48538 8891
rect 50629 8857 50663 8891
rect 51794 8857 51828 8891
rect 1409 8789 1443 8823
rect 2237 8789 2271 8823
rect 2881 8789 2915 8823
rect 14289 8789 14323 8823
rect 14473 8789 14507 8823
rect 15025 8789 15059 8823
rect 19625 8789 19659 8823
rect 27813 8789 27847 8823
rect 28457 8789 28491 8823
rect 36461 8789 36495 8823
rect 42349 8789 42383 8823
rect 45017 8789 45051 8823
rect 46489 8789 46523 8823
rect 49617 8789 49651 8823
rect 52929 8789 52963 8823
rect 5181 8585 5215 8619
rect 19901 8585 19935 8619
rect 22477 8585 22511 8619
rect 25329 8585 25363 8619
rect 33701 8585 33735 8619
rect 39681 8585 39715 8619
rect 48605 8585 48639 8619
rect 50461 8585 50495 8619
rect 50629 8585 50663 8619
rect 2228 8517 2262 8551
rect 5549 8517 5583 8551
rect 22201 8517 22235 8551
rect 24961 8517 24995 8551
rect 27629 8517 27663 8551
rect 27813 8517 27847 8551
rect 28457 8517 28491 8551
rect 28733 8517 28767 8551
rect 28933 8517 28967 8551
rect 33333 8517 33367 8551
rect 42809 8517 42843 8551
rect 42927 8517 42961 8551
rect 44741 8517 44775 8551
rect 45017 8517 45051 8551
rect 45109 8517 45143 8551
rect 45227 8517 45261 8551
rect 50261 8517 50295 8551
rect 1961 8449 1995 8483
rect 5365 8449 5399 8483
rect 5641 8449 5675 8483
rect 16957 8449 16991 8483
rect 18521 8449 18555 8483
rect 18788 8449 18822 8483
rect 21833 8449 21867 8483
rect 21953 8449 21987 8483
rect 22109 8449 22143 8483
rect 22339 8449 22373 8483
rect 24685 8449 24719 8483
rect 24778 8449 24812 8483
rect 25053 8449 25087 8483
rect 25191 8449 25225 8483
rect 30205 8449 30239 8483
rect 30481 8449 30515 8483
rect 32137 8449 32171 8483
rect 33517 8449 33551 8483
rect 35265 8449 35299 8483
rect 36185 8449 36219 8483
rect 37749 8449 37783 8483
rect 38761 8449 38795 8483
rect 38945 8449 38979 8483
rect 39589 8449 39623 8483
rect 41613 8449 41647 8483
rect 41889 8449 41923 8483
rect 42625 8449 42659 8483
rect 42717 8449 42751 8483
rect 44925 8449 44959 8483
rect 48789 8449 48823 8483
rect 48973 8449 49007 8483
rect 49065 8449 49099 8483
rect 15301 8381 15335 8415
rect 15577 8381 15611 8415
rect 16681 8381 16715 8415
rect 35081 8381 35115 8415
rect 43085 8381 43119 8415
rect 45385 8381 45419 8415
rect 3341 8313 3375 8347
rect 27997 8313 28031 8347
rect 29101 8313 29135 8347
rect 32321 8313 32355 8347
rect 36369 8313 36403 8347
rect 37933 8313 37967 8347
rect 41797 8313 41831 8347
rect 42441 8313 42475 8347
rect 27813 8245 27847 8279
rect 28917 8245 28951 8279
rect 35449 8245 35483 8279
rect 38761 8245 38795 8279
rect 41429 8245 41463 8279
rect 50445 8245 50479 8279
rect 6009 8041 6043 8075
rect 9321 8041 9355 8075
rect 10149 8041 10183 8075
rect 13093 8041 13127 8075
rect 14289 8041 14323 8075
rect 19257 8041 19291 8075
rect 24685 8041 24719 8075
rect 25145 8041 25179 8075
rect 25504 8041 25538 8075
rect 27537 8041 27571 8075
rect 29745 8041 29779 8075
rect 46489 8041 46523 8075
rect 52929 8041 52963 8075
rect 4169 7973 4203 8007
rect 27721 7973 27755 8007
rect 33057 7973 33091 8007
rect 35081 7973 35115 8007
rect 38761 7973 38795 8007
rect 42625 7973 42659 8007
rect 1409 7905 1443 7939
rect 1685 7905 1719 7939
rect 4629 7905 4663 7939
rect 11713 7905 11747 7939
rect 15669 7905 15703 7939
rect 41245 7905 41279 7939
rect 45293 7905 45327 7939
rect 2697 7837 2731 7871
rect 8125 7837 8159 7871
rect 9045 7837 9079 7871
rect 10057 7837 10091 7871
rect 15485 7837 15519 7871
rect 15577 7837 15611 7871
rect 15761 7837 15795 7871
rect 19441 7837 19475 7871
rect 19717 7837 19751 7871
rect 28181 7837 28215 7871
rect 28457 7837 28491 7871
rect 31033 7837 31067 7871
rect 32873 7837 32907 7871
rect 34713 7837 34747 7871
rect 37841 7837 37875 7871
rect 38025 7837 38059 7871
rect 38577 7837 38611 7871
rect 41512 7837 41546 7871
rect 45017 7837 45051 7871
rect 52745 7837 52779 7871
rect 53021 7837 53055 7871
rect 3985 7769 4019 7803
rect 4896 7769 4930 7803
rect 11980 7769 12014 7803
rect 14105 7769 14139 7803
rect 14305 7769 14339 7803
rect 19625 7769 19659 7803
rect 24501 7769 24535 7803
rect 24717 7769 24751 7803
rect 25329 7769 25363 7803
rect 26249 7769 26283 7803
rect 27353 7769 27387 7803
rect 29561 7769 29595 7803
rect 31300 7769 31334 7803
rect 34897 7769 34931 7803
rect 46397 7769 46431 7803
rect 2881 7701 2915 7735
rect 8217 7701 8251 7735
rect 9505 7701 9539 7735
rect 10517 7701 10551 7735
rect 14473 7701 14507 7735
rect 15301 7701 15335 7735
rect 24869 7701 24903 7735
rect 25529 7701 25563 7735
rect 25697 7701 25731 7735
rect 26341 7701 26375 7735
rect 27563 7701 27597 7735
rect 29761 7701 29795 7735
rect 29929 7701 29963 7735
rect 32413 7701 32447 7735
rect 37933 7701 37967 7735
rect 52561 7701 52595 7735
rect 2605 7497 2639 7531
rect 5273 7497 5307 7531
rect 12633 7497 12667 7531
rect 13001 7497 13035 7531
rect 16681 7497 16715 7531
rect 19467 7497 19501 7531
rect 20469 7497 20503 7531
rect 25145 7497 25179 7531
rect 32137 7497 32171 7531
rect 54861 7497 54895 7531
rect 2513 7429 2547 7463
rect 5641 7429 5675 7463
rect 7665 7429 7699 7463
rect 11897 7429 11931 7463
rect 19257 7429 19291 7463
rect 20269 7429 20303 7463
rect 23121 7429 23155 7463
rect 24133 7429 24167 7463
rect 24349 7429 24383 7463
rect 27813 7429 27847 7463
rect 27997 7429 28031 7463
rect 28733 7429 28767 7463
rect 28933 7429 28967 7463
rect 30941 7429 30975 7463
rect 42809 7429 42843 7463
rect 43361 7429 43395 7463
rect 46213 7429 46247 7463
rect 49157 7429 49191 7463
rect 50322 7429 50356 7463
rect 53726 7429 53760 7463
rect 1501 7361 1535 7395
rect 3525 7361 3559 7395
rect 5457 7361 5491 7395
rect 5733 7361 5767 7395
rect 7757 7361 7791 7395
rect 8769 7361 8803 7395
rect 9045 7361 9079 7395
rect 10241 7361 10275 7395
rect 11529 7361 11563 7395
rect 11713 7361 11747 7395
rect 12817 7361 12851 7395
rect 13093 7361 13127 7395
rect 15577 7361 15611 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 22937 7361 22971 7395
rect 23213 7361 23247 7395
rect 25053 7361 25087 7395
rect 25697 7361 25731 7395
rect 30205 7361 30239 7395
rect 30389 7361 30423 7395
rect 31125 7361 31159 7395
rect 32321 7361 32355 7395
rect 34897 7361 34931 7395
rect 35081 7361 35115 7395
rect 35173 7361 35207 7395
rect 35265 7361 35299 7395
rect 35449 7361 35483 7395
rect 38005 7361 38039 7395
rect 42625 7361 42659 7395
rect 42717 7361 42751 7395
rect 42927 7361 42961 7395
rect 44373 7361 44407 7395
rect 44557 7361 44591 7395
rect 44649 7361 44683 7395
rect 44787 7361 44821 7395
rect 46029 7361 46063 7395
rect 46305 7361 46339 7395
rect 46397 7361 46431 7395
rect 49341 7361 49375 7395
rect 49525 7361 49559 7395
rect 53481 7361 53515 7395
rect 2697 7293 2731 7327
rect 8125 7293 8159 7327
rect 8217 7293 8251 7327
rect 10057 7293 10091 7327
rect 15301 7293 15335 7327
rect 16957 7293 16991 7327
rect 17141 7293 17175 7327
rect 32597 7293 32631 7327
rect 37749 7293 37783 7327
rect 43085 7293 43119 7327
rect 49617 7293 49651 7327
rect 50077 7293 50111 7327
rect 19625 7225 19659 7259
rect 20637 7225 20671 7259
rect 32505 7225 32539 7259
rect 1593 7157 1627 7191
rect 2145 7157 2179 7191
rect 3341 7157 3375 7191
rect 10425 7157 10459 7191
rect 19441 7157 19475 7191
rect 19901 7157 19935 7191
rect 20453 7157 20487 7191
rect 22753 7157 22787 7191
rect 24317 7157 24351 7191
rect 24501 7157 24535 7191
rect 25881 7157 25915 7191
rect 27997 7157 28031 7191
rect 28181 7157 28215 7191
rect 28917 7157 28951 7191
rect 29101 7157 29135 7191
rect 35633 7157 35667 7191
rect 39129 7157 39163 7191
rect 42441 7157 42475 7191
rect 44925 7157 44959 7191
rect 46581 7157 46615 7191
rect 51457 7157 51491 7191
rect 23489 6953 23523 6987
rect 27997 6953 28031 6987
rect 37473 6953 37507 6987
rect 30665 6885 30699 6919
rect 1685 6817 1719 6851
rect 15669 6817 15703 6851
rect 17141 6817 17175 6851
rect 17233 6817 17267 6851
rect 17417 6817 17451 6851
rect 37105 6817 37139 6851
rect 45017 6817 45051 6851
rect 1409 6749 1443 6783
rect 2881 6749 2915 6783
rect 6101 6749 6135 6783
rect 6285 6749 6319 6783
rect 6377 6749 6411 6783
rect 9413 6749 9447 6783
rect 9781 6749 9815 6783
rect 14289 6749 14323 6783
rect 14565 6749 14599 6783
rect 15945 6749 15979 6783
rect 17325 6749 17359 6783
rect 19441 6749 19475 6783
rect 19717 6749 19751 6783
rect 22109 6749 22143 6783
rect 22376 6749 22410 6783
rect 30481 6749 30515 6783
rect 32321 6749 32355 6783
rect 32597 6749 32631 6783
rect 32689 6749 32723 6783
rect 34805 6749 34839 6783
rect 35072 6749 35106 6783
rect 36737 6749 36771 6783
rect 36921 6749 36955 6783
rect 37013 6749 37047 6783
rect 37289 6749 37323 6783
rect 47133 6749 47167 6783
rect 47389 6749 47423 6783
rect 49341 6749 49375 6783
rect 49525 6749 49559 6783
rect 49617 6749 49651 6783
rect 52653 6749 52687 6783
rect 52837 6749 52871 6783
rect 52929 6749 52963 6783
rect 19625 6681 19659 6715
rect 24869 6681 24903 6715
rect 27813 6681 27847 6715
rect 32505 6681 32539 6715
rect 41337 6681 41371 6715
rect 45284 6681 45318 6715
rect 2697 6613 2731 6647
rect 5917 6613 5951 6647
rect 14105 6613 14139 6647
rect 14473 6613 14507 6647
rect 16957 6613 16991 6647
rect 19257 6613 19291 6647
rect 24961 6613 24995 6647
rect 28013 6613 28047 6647
rect 28181 6613 28215 6647
rect 32873 6613 32907 6647
rect 36185 6613 36219 6647
rect 41429 6613 41463 6647
rect 46397 6613 46431 6647
rect 48513 6613 48547 6647
rect 49157 6613 49191 6647
rect 52469 6613 52503 6647
rect 2605 6409 2639 6443
rect 15209 6409 15243 6443
rect 33517 6409 33551 6443
rect 36645 6409 36679 6443
rect 44557 6409 44591 6443
rect 46765 6409 46799 6443
rect 49157 6409 49191 6443
rect 50169 6409 50203 6443
rect 53297 6409 53331 6443
rect 6622 6341 6656 6375
rect 13360 6341 13394 6375
rect 18512 6341 18546 6375
rect 22477 6341 22511 6375
rect 22661 6341 22695 6375
rect 29469 6341 29503 6375
rect 29685 6341 29719 6375
rect 32404 6341 32438 6375
rect 44189 6341 44223 6375
rect 44281 6341 44315 6375
rect 46397 6341 46431 6375
rect 46489 6341 46523 6375
rect 48881 6341 48915 6375
rect 49893 6341 49927 6375
rect 52929 6341 52963 6375
rect 1409 6273 1443 6307
rect 2513 6273 2547 6307
rect 4997 6273 5031 6307
rect 5181 6273 5215 6307
rect 5273 6273 5307 6307
rect 8861 6273 8895 6307
rect 13093 6273 13127 6307
rect 15393 6273 15427 6307
rect 15485 6273 15519 6307
rect 15669 6273 15703 6307
rect 17049 6273 17083 6307
rect 17141 6273 17175 6307
rect 18245 6273 18279 6307
rect 22293 6273 22327 6307
rect 22385 6273 22419 6307
rect 36277 6273 36311 6307
rect 36461 6273 36495 6307
rect 39957 6273 39991 6307
rect 40141 6273 40175 6307
rect 42901 6273 42935 6307
rect 43085 6273 43119 6307
rect 44005 6273 44039 6307
rect 44373 6273 44407 6307
rect 46213 6273 46247 6307
rect 46581 6273 46615 6307
rect 48605 6273 48639 6307
rect 48789 6273 48823 6307
rect 48973 6273 49007 6307
rect 49617 6273 49651 6307
rect 49755 6273 49789 6307
rect 49985 6273 50019 6307
rect 52745 6273 52779 6307
rect 53021 6273 53055 6307
rect 53113 6273 53147 6307
rect 2697 6205 2731 6239
rect 6377 6205 6411 6239
rect 9137 6205 9171 6239
rect 15577 6205 15611 6239
rect 16865 6205 16899 6239
rect 16957 6205 16991 6239
rect 32137 6205 32171 6239
rect 40233 6205 40267 6239
rect 43177 6205 43211 6239
rect 9045 6137 9079 6171
rect 16681 6137 16715 6171
rect 22109 6137 22143 6171
rect 1593 6069 1627 6103
rect 2145 6069 2179 6103
rect 4813 6069 4847 6103
rect 7757 6069 7791 6103
rect 8677 6069 8711 6103
rect 14473 6069 14507 6103
rect 19625 6069 19659 6103
rect 29653 6069 29687 6103
rect 29837 6069 29871 6103
rect 39773 6069 39807 6103
rect 42717 6069 42751 6103
rect 5457 5865 5491 5899
rect 12265 5865 12299 5899
rect 15209 5865 15243 5899
rect 21465 5865 21499 5899
rect 29745 5865 29779 5899
rect 52561 5865 52595 5899
rect 21097 5797 21131 5831
rect 22339 5797 22373 5831
rect 32873 5797 32907 5831
rect 38301 5797 38335 5831
rect 1869 5729 1903 5763
rect 10149 5729 10183 5763
rect 10333 5729 10367 5763
rect 15577 5729 15611 5763
rect 15669 5729 15703 5763
rect 23765 5729 23799 5763
rect 26801 5729 26835 5763
rect 35541 5729 35575 5763
rect 36645 5729 36679 5763
rect 39865 5729 39899 5763
rect 42349 5729 42383 5763
rect 2136 5661 2170 5695
rect 4077 5661 4111 5695
rect 4344 5661 4378 5695
rect 8953 5661 8987 5695
rect 9137 5661 9171 5695
rect 10885 5661 10919 5695
rect 15393 5661 15427 5695
rect 15485 5661 15519 5695
rect 22109 5661 22143 5695
rect 23397 5661 23431 5695
rect 25238 5671 25272 5705
rect 25422 5661 25456 5695
rect 25697 5661 25731 5695
rect 26341 5661 26375 5695
rect 27445 5661 27479 5695
rect 27629 5661 27663 5695
rect 27747 5661 27781 5695
rect 27905 5661 27939 5695
rect 28549 5661 28583 5695
rect 28733 5661 28767 5695
rect 28851 5661 28885 5695
rect 29009 5661 29043 5695
rect 32321 5661 32355 5695
rect 32689 5661 32723 5695
rect 35725 5661 35759 5695
rect 36461 5661 36495 5695
rect 38117 5661 38151 5695
rect 40121 5661 40155 5695
rect 41889 5661 41923 5695
rect 41981 5661 42015 5695
rect 42211 5661 42245 5695
rect 42993 5661 43027 5695
rect 43295 5661 43329 5695
rect 43453 5661 43487 5695
rect 52009 5661 52043 5695
rect 52193 5661 52227 5695
rect 52377 5661 52411 5695
rect 53021 5661 53055 5695
rect 53288 5661 53322 5695
rect 11152 5593 11186 5627
rect 21465 5593 21499 5627
rect 23581 5593 23615 5627
rect 25329 5593 25363 5627
rect 25539 5593 25573 5627
rect 26434 5593 26468 5627
rect 26525 5593 26559 5627
rect 26663 5593 26697 5627
rect 27537 5593 27571 5627
rect 28641 5593 28675 5627
rect 29561 5593 29595 5627
rect 29777 5593 29811 5627
rect 32505 5593 32539 5627
rect 32597 5593 32631 5627
rect 42073 5593 42107 5627
rect 43085 5593 43119 5627
rect 43177 5593 43211 5627
rect 46213 5593 46247 5627
rect 46397 5593 46431 5627
rect 52285 5593 52319 5627
rect 3249 5525 3283 5559
rect 9045 5525 9079 5559
rect 9689 5525 9723 5559
rect 10057 5525 10091 5559
rect 21649 5525 21683 5559
rect 25053 5525 25087 5559
rect 26157 5525 26191 5559
rect 27261 5525 27295 5559
rect 28365 5525 28399 5559
rect 29929 5525 29963 5559
rect 35909 5525 35943 5559
rect 41245 5525 41279 5559
rect 41705 5525 41739 5559
rect 42809 5525 42843 5559
rect 54401 5525 54435 5559
rect 4721 5321 4755 5355
rect 8769 5321 8803 5355
rect 10793 5321 10827 5355
rect 22385 5321 22419 5355
rect 32873 5321 32907 5355
rect 36093 5321 36127 5355
rect 36553 5321 36587 5355
rect 38761 5321 38795 5355
rect 40693 5321 40727 5355
rect 43085 5321 43119 5355
rect 50997 5321 51031 5355
rect 1869 5253 1903 5287
rect 31309 5253 31343 5287
rect 32597 5253 32631 5287
rect 34980 5253 35014 5287
rect 40325 5253 40359 5287
rect 42717 5253 42751 5287
rect 42917 5253 42951 5287
rect 45385 5253 45419 5287
rect 2697 5185 2731 5219
rect 3617 5185 3651 5219
rect 4261 5185 4295 5219
rect 4905 5185 4939 5219
rect 7645 5185 7679 5219
rect 10977 5185 11011 5219
rect 14841 5185 14875 5219
rect 15025 5185 15059 5219
rect 15117 5185 15151 5219
rect 18429 5185 18463 5219
rect 19073 5185 19107 5219
rect 19257 5185 19291 5219
rect 22017 5185 22051 5219
rect 22109 5185 22143 5219
rect 22201 5185 22235 5219
rect 25697 5185 25731 5219
rect 25881 5185 25915 5219
rect 27813 5185 27847 5219
rect 27997 5185 28031 5219
rect 28089 5185 28123 5219
rect 28825 5185 28859 5219
rect 29009 5185 29043 5219
rect 29101 5185 29135 5219
rect 32321 5185 32355 5219
rect 32505 5185 32539 5219
rect 32689 5185 32723 5219
rect 36737 5185 36771 5219
rect 38669 5185 38703 5219
rect 40141 5185 40175 5219
rect 40417 5185 40451 5219
rect 40533 5185 40567 5219
rect 46213 5185 46247 5219
rect 49873 5185 49907 5219
rect 7389 5117 7423 5151
rect 21833 5117 21867 5151
rect 25973 5117 26007 5151
rect 29929 5117 29963 5151
rect 30205 5117 30239 5151
rect 34713 5117 34747 5151
rect 37289 5117 37323 5151
rect 37565 5117 37599 5151
rect 46489 5117 46523 5151
rect 49617 5117 49651 5151
rect 46397 5049 46431 5083
rect 2145 4981 2179 5015
rect 2881 4981 2915 5015
rect 3433 4981 3467 5015
rect 4077 4981 4111 5015
rect 14657 4981 14691 5015
rect 18521 4981 18555 5015
rect 19441 4981 19475 5015
rect 25513 4981 25547 5015
rect 27629 4981 27663 5015
rect 28641 4981 28675 5015
rect 31401 4981 31435 5015
rect 42901 4981 42935 5015
rect 45477 4981 45511 5015
rect 46029 4981 46063 5015
rect 2053 4777 2087 4811
rect 7297 4777 7331 4811
rect 10333 4777 10367 4811
rect 15485 4777 15519 4811
rect 21281 4777 21315 4811
rect 24777 4777 24811 4811
rect 25697 4777 25731 4811
rect 26525 4777 26559 4811
rect 27353 4777 27387 4811
rect 27537 4777 27571 4811
rect 42533 4777 42567 4811
rect 43453 4777 43487 4811
rect 46489 4777 46523 4811
rect 2329 4709 2363 4743
rect 5273 4709 5307 4743
rect 47317 4709 47351 4743
rect 7113 4641 7147 4675
rect 11621 4641 11655 4675
rect 14105 4641 14139 4675
rect 15945 4641 15979 4675
rect 19441 4641 19475 4675
rect 19533 4641 19567 4675
rect 20361 4641 20395 4675
rect 21465 4641 21499 4675
rect 21649 4641 21683 4675
rect 40877 4641 40911 4675
rect 1409 4573 1443 4607
rect 2145 4573 2179 4607
rect 2881 4573 2915 4607
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 5457 4573 5491 4607
rect 6101 4573 6135 4607
rect 7573 4573 7607 4607
rect 8953 4573 8987 4607
rect 11805 4573 11839 4607
rect 14372 4573 14406 4607
rect 16221 4573 16255 4607
rect 18521 4573 18555 4607
rect 19625 4573 19659 4607
rect 19717 4573 19751 4607
rect 20269 4573 20303 4607
rect 20453 4573 20487 4607
rect 21557 4573 21591 4607
rect 21741 4573 21775 4607
rect 24593 4573 24627 4607
rect 24869 4573 24903 4607
rect 25513 4573 25547 4607
rect 25789 4573 25823 4607
rect 32045 4573 32079 4607
rect 32321 4573 32355 4607
rect 32413 4573 32447 4607
rect 35633 4573 35667 4607
rect 35726 4573 35760 4607
rect 36001 4573 36035 4607
rect 36139 4573 36173 4607
rect 36829 4573 36863 4607
rect 37013 4573 37047 4607
rect 38209 4573 38243 4607
rect 42349 4573 42383 4607
rect 42625 4573 42659 4607
rect 43269 4573 43303 4607
rect 43545 4573 43579 4607
rect 45937 4573 45971 4607
rect 46121 4573 46155 4607
rect 46305 4573 46339 4607
rect 47133 4573 47167 4607
rect 47409 4573 47443 4607
rect 48237 4573 48271 4607
rect 9198 4505 9232 4539
rect 18337 4505 18371 4539
rect 26341 4505 26375 4539
rect 26557 4505 26591 4539
rect 27169 4505 27203 4539
rect 32229 4505 32263 4539
rect 35909 4505 35943 4539
rect 40693 4505 40727 4539
rect 46213 4505 46247 4539
rect 46949 4505 46983 4539
rect 48482 4505 48516 4539
rect 1593 4437 1627 4471
rect 3065 4437 3099 4471
rect 4629 4437 4663 4471
rect 5917 4437 5951 4471
rect 7481 4437 7515 4471
rect 11989 4437 12023 4471
rect 18705 4437 18739 4471
rect 19257 4437 19291 4471
rect 24409 4437 24443 4471
rect 25329 4437 25363 4471
rect 26709 4437 26743 4471
rect 27369 4437 27403 4471
rect 32597 4437 32631 4471
rect 36277 4437 36311 4471
rect 38301 4437 38335 4471
rect 42165 4437 42199 4471
rect 43085 4437 43119 4471
rect 49617 4437 49651 4471
rect 42825 4233 42859 4267
rect 42993 4233 43027 4267
rect 43821 4233 43855 4267
rect 28540 4165 28574 4199
rect 36001 4165 36035 4199
rect 42625 4165 42659 4199
rect 43453 4165 43487 4199
rect 46121 4165 46155 4199
rect 43683 4131 43717 4165
rect 1409 4097 1443 4131
rect 2145 4097 2179 4131
rect 2412 4097 2446 4131
rect 3985 4097 4019 4131
rect 4169 4097 4203 4131
rect 4813 4097 4847 4131
rect 5641 4097 5675 4131
rect 6561 4097 6595 4131
rect 8079 4097 8113 4131
rect 8217 4097 8251 4131
rect 8330 4097 8364 4131
rect 8493 4097 8527 4131
rect 10701 4097 10735 4131
rect 11529 4097 11563 4131
rect 16681 4097 16715 4131
rect 18245 4097 18279 4131
rect 18429 4097 18463 4131
rect 19165 4097 19199 4131
rect 22017 4097 22051 4131
rect 34529 4097 34563 4131
rect 34713 4097 34747 4131
rect 34897 4097 34931 4131
rect 35081 4097 35115 4131
rect 35725 4097 35759 4131
rect 35818 4097 35852 4131
rect 36093 4097 36127 4131
rect 36190 4097 36224 4131
rect 38485 4097 38519 4131
rect 38578 4097 38612 4131
rect 38761 4097 38795 4131
rect 38853 4097 38887 4131
rect 38991 4097 39025 4131
rect 40049 4097 40083 4131
rect 41245 4097 41279 4131
rect 45937 4097 45971 4131
rect 46213 4097 46247 4131
rect 46305 4097 46339 4131
rect 7849 4029 7883 4063
rect 11805 4029 11839 4063
rect 15025 4029 15059 4063
rect 15301 4029 15335 4063
rect 16957 4029 16991 4063
rect 18337 4029 18371 4063
rect 19073 4029 19107 4063
rect 19257 4029 19291 4063
rect 19349 4029 19383 4063
rect 28273 4029 28307 4063
rect 34805 4029 34839 4063
rect 6377 3961 6411 3995
rect 46489 3961 46523 3995
rect 1593 3893 1627 3927
rect 3525 3893 3559 3927
rect 4077 3893 4111 3927
rect 5457 3893 5491 3927
rect 10517 3893 10551 3927
rect 18889 3893 18923 3927
rect 21833 3893 21867 3927
rect 29653 3893 29687 3927
rect 35265 3893 35299 3927
rect 36369 3893 36403 3927
rect 39129 3893 39163 3927
rect 39865 3893 39899 3927
rect 41429 3893 41463 3927
rect 42809 3893 42843 3927
rect 43637 3893 43671 3927
rect 35127 3689 35161 3723
rect 40233 3689 40267 3723
rect 7941 3621 7975 3655
rect 13369 3621 13403 3655
rect 15577 3621 15611 3655
rect 23673 3621 23707 3655
rect 25789 3621 25823 3655
rect 43545 3621 43579 3655
rect 4445 3553 4479 3587
rect 4813 3553 4847 3587
rect 5273 3553 5307 3587
rect 7113 3553 7147 3587
rect 31493 3553 31527 3587
rect 33701 3553 33735 3587
rect 33793 3553 33827 3587
rect 37381 3553 37415 3587
rect 46489 3553 46523 3587
rect 1869 3485 1903 3519
rect 2697 3485 2731 3519
rect 3985 3485 4019 3519
rect 4629 3485 4663 3519
rect 7297 3485 7331 3519
rect 7481 3485 7515 3519
rect 8125 3485 8159 3519
rect 10057 3485 10091 3519
rect 10333 3485 10367 3519
rect 10517 3485 10551 3519
rect 10977 3485 11011 3519
rect 11161 3485 11195 3519
rect 11805 3485 11839 3519
rect 11989 3485 12023 3519
rect 13553 3485 13587 3519
rect 14933 3485 14967 3519
rect 15026 3485 15060 3519
rect 15301 3485 15335 3519
rect 15439 3485 15473 3519
rect 16037 3485 16071 3519
rect 16185 3485 16219 3519
rect 16502 3485 16536 3519
rect 17325 3485 17359 3519
rect 19441 3485 19475 3519
rect 20269 3485 20303 3519
rect 21373 3485 21407 3519
rect 23857 3485 23891 3519
rect 24409 3485 24443 3519
rect 24676 3485 24710 3519
rect 26249 3485 26283 3519
rect 26505 3485 26539 3519
rect 28273 3485 28307 3519
rect 30665 3485 30699 3519
rect 31125 3485 31159 3519
rect 31309 3485 31343 3519
rect 33425 3485 33459 3519
rect 33613 3485 33647 3519
rect 33977 3485 34011 3519
rect 34897 3485 34931 3519
rect 36185 3485 36219 3519
rect 37105 3485 37139 3519
rect 37289 3485 37323 3519
rect 37473 3485 37507 3519
rect 37657 3485 37691 3519
rect 38301 3485 38335 3519
rect 39865 3485 39899 3519
rect 40049 3485 40083 3519
rect 41429 3485 41463 3519
rect 42165 3485 42199 3519
rect 42421 3485 42455 3519
rect 45569 3485 45603 3519
rect 57713 3485 57747 3519
rect 2237 3417 2271 3451
rect 5540 3417 5574 3451
rect 12633 3417 12667 3451
rect 15209 3417 15243 3451
rect 16313 3417 16347 3451
rect 16405 3417 16439 3451
rect 46756 3417 46790 3451
rect 57989 3417 58023 3451
rect 2881 3349 2915 3383
rect 3801 3349 3835 3383
rect 6653 3349 6687 3383
rect 9873 3349 9907 3383
rect 11345 3349 11379 3383
rect 12173 3349 12207 3383
rect 14105 3349 14139 3383
rect 16681 3349 16715 3383
rect 17141 3349 17175 3383
rect 19257 3349 19291 3383
rect 20453 3349 20487 3383
rect 21189 3349 21223 3383
rect 27629 3349 27663 3383
rect 28089 3349 28123 3383
rect 30481 3349 30515 3383
rect 34161 3349 34195 3383
rect 36369 3349 36403 3383
rect 37841 3349 37875 3383
rect 38485 3349 38519 3383
rect 41613 3349 41647 3383
rect 45753 3349 45787 3383
rect 47869 3349 47903 3383
rect 1593 3145 1627 3179
rect 3893 3145 3927 3179
rect 4721 3145 4755 3179
rect 6377 3145 6411 3179
rect 33517 3145 33551 3179
rect 38761 3145 38795 3179
rect 41153 3145 41187 3179
rect 47777 3145 47811 3179
rect 9864 3077 9898 3111
rect 14933 3077 14967 3111
rect 18972 3077 19006 3111
rect 22100 3077 22134 3111
rect 23940 3077 23974 3111
rect 27620 3077 27654 3111
rect 30472 3077 30506 3111
rect 32404 3077 32438 3111
rect 34704 3077 34738 3111
rect 37648 3077 37682 3111
rect 40018 3077 40052 3111
rect 43812 3077 43846 3111
rect 45814 3077 45848 3111
rect 57161 3077 57195 3111
rect 1409 3009 1443 3043
rect 2697 3009 2731 3043
rect 3709 3009 3743 3043
rect 4261 3009 4295 3043
rect 4537 3009 4571 3043
rect 5273 3009 5307 3043
rect 6561 3009 6595 3043
rect 7297 3009 7331 3043
rect 8309 3009 8343 3043
rect 11713 3009 11747 3043
rect 12817 3009 12851 3043
rect 13461 3009 13495 3043
rect 13921 3009 13955 3043
rect 14664 3009 14698 3043
rect 14777 3009 14811 3043
rect 15025 3009 15059 3043
rect 15163 3009 15197 3043
rect 15761 3009 15795 3043
rect 16688 3009 16722 3043
rect 16774 3009 16808 3043
rect 16957 3009 16991 3043
rect 17049 3009 17083 3043
rect 17146 3009 17180 3043
rect 17785 3009 17819 3043
rect 20637 3009 20671 3043
rect 23673 3009 23707 3043
rect 26249 3009 26283 3043
rect 30205 3009 30239 3043
rect 32137 3009 32171 3043
rect 34437 3009 34471 3043
rect 36277 3009 36311 3043
rect 37381 3009 37415 3043
rect 39773 3009 39807 3043
rect 42717 3009 42751 3043
rect 47593 3009 47627 3043
rect 48329 3009 48363 3043
rect 49985 3009 50019 3043
rect 51457 3009 51491 3043
rect 52929 3009 52963 3043
rect 54401 3009 54435 3043
rect 55873 3009 55907 3043
rect 56885 3009 56919 3043
rect 57897 3009 57931 3043
rect 3525 2941 3559 2975
rect 6837 2941 6871 2975
rect 8769 2941 8803 2975
rect 9597 2941 9631 2975
rect 18705 2941 18739 2975
rect 21833 2941 21867 2975
rect 27353 2941 27387 2975
rect 43545 2941 43579 2975
rect 45569 2941 45603 2975
rect 5457 2873 5491 2907
rect 7481 2873 7515 2907
rect 10977 2873 11011 2907
rect 12633 2873 12667 2907
rect 13277 2873 13311 2907
rect 15945 2873 15979 2907
rect 17325 2873 17359 2907
rect 25053 2873 25087 2907
rect 26065 2873 26099 2907
rect 28733 2873 28767 2907
rect 36461 2873 36495 2907
rect 44925 2873 44959 2907
rect 48513 2873 48547 2907
rect 2881 2805 2915 2839
rect 6745 2805 6779 2839
rect 8125 2805 8159 2839
rect 11529 2805 11563 2839
rect 14105 2805 14139 2839
rect 15301 2805 15335 2839
rect 17969 2805 18003 2839
rect 20085 2805 20119 2839
rect 20821 2805 20855 2839
rect 23213 2805 23247 2839
rect 31585 2805 31619 2839
rect 35817 2805 35851 2839
rect 42901 2805 42935 2839
rect 46949 2805 46983 2839
rect 50169 2805 50203 2839
rect 51641 2805 51675 2839
rect 53113 2805 53147 2839
rect 54585 2805 54619 2839
rect 56057 2805 56091 2839
rect 58081 2805 58115 2839
rect 2789 2601 2823 2635
rect 15301 2601 15335 2635
rect 28825 2601 28859 2635
rect 30297 2601 30331 2635
rect 38025 2601 38059 2635
rect 38761 2601 38795 2635
rect 7297 2533 7331 2567
rect 10609 2533 10643 2567
rect 13185 2533 13219 2567
rect 26065 2533 26099 2567
rect 43085 2533 43119 2567
rect 19257 2465 19291 2499
rect 32413 2465 32447 2499
rect 34713 2465 34747 2499
rect 34989 2465 35023 2499
rect 40509 2465 40543 2499
rect 3801 2397 3835 2431
rect 4629 2397 4663 2431
rect 4905 2397 4939 2431
rect 6377 2397 6411 2431
rect 7113 2397 7147 2431
rect 8953 2397 8987 2431
rect 9505 2397 9539 2431
rect 10149 2397 10183 2431
rect 10425 2397 10459 2431
rect 11529 2397 11563 2431
rect 12081 2397 12115 2431
rect 12725 2397 12759 2431
rect 13001 2397 13035 2431
rect 14657 2397 14691 2431
rect 14805 2397 14839 2431
rect 14933 2397 14967 2431
rect 15025 2397 15059 2431
rect 15163 2397 15197 2431
rect 15761 2397 15795 2431
rect 16865 2397 16899 2431
rect 17601 2397 17635 2431
rect 18429 2397 18463 2431
rect 19524 2397 19558 2431
rect 21833 2397 21867 2431
rect 22569 2397 22603 2431
rect 23305 2397 23339 2431
rect 24409 2397 24443 2431
rect 25145 2397 25179 2431
rect 25881 2397 25915 2431
rect 26985 2397 27019 2431
rect 28089 2397 28123 2431
rect 29009 2397 29043 2431
rect 29561 2397 29595 2431
rect 30481 2397 30515 2431
rect 30941 2397 30975 2431
rect 32137 2397 32171 2431
rect 33425 2397 33459 2431
rect 38577 2397 38611 2431
rect 48789 2397 48823 2431
rect 52745 2397 52779 2431
rect 53941 2397 53975 2431
rect 55321 2397 55355 2431
rect 56793 2397 56827 2431
rect 57897 2397 57931 2431
rect 1501 2329 1535 2363
rect 7849 2329 7883 2363
rect 36461 2329 36495 2363
rect 37933 2329 37967 2363
rect 40325 2329 40359 2363
rect 41061 2329 41095 2363
rect 42901 2329 42935 2363
rect 43729 2329 43763 2363
rect 45477 2329 45511 2363
rect 46673 2329 46707 2363
rect 48145 2329 48179 2363
rect 50629 2329 50663 2363
rect 51549 2329 51583 2363
rect 53021 2329 53055 2363
rect 54217 2329 54251 2363
rect 55597 2329 55631 2363
rect 57069 2329 57103 2363
rect 3985 2261 4019 2295
rect 6561 2261 6595 2295
rect 9137 2261 9171 2295
rect 9689 2261 9723 2295
rect 11713 2261 11747 2295
rect 12265 2261 12299 2295
rect 15945 2261 15979 2295
rect 17049 2261 17083 2295
rect 17785 2261 17819 2295
rect 18613 2261 18647 2295
rect 20637 2261 20671 2295
rect 22017 2261 22051 2295
rect 22753 2261 22787 2295
rect 23489 2261 23523 2295
rect 24593 2261 24627 2295
rect 25329 2261 25363 2295
rect 27169 2261 27203 2295
rect 28273 2261 28307 2295
rect 29745 2261 29779 2295
rect 31125 2261 31159 2295
rect 33609 2261 33643 2295
rect 36553 2261 36587 2295
rect 41153 2261 41187 2295
rect 43821 2261 43855 2295
rect 45569 2261 45603 2295
rect 46765 2261 46799 2295
rect 48237 2261 48271 2295
rect 48973 2261 49007 2295
rect 50721 2261 50755 2295
rect 51641 2261 51675 2295
rect 58081 2261 58115 2295
<< metal1 >>
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 2317 39627 2375 39633
rect 2317 39593 2329 39627
rect 2363 39624 2375 39627
rect 2774 39624 2780 39636
rect 2363 39596 2780 39624
rect 2363 39593 2375 39596
rect 2317 39587 2375 39593
rect 2774 39584 2780 39596
rect 2832 39584 2838 39636
rect 3050 39624 3056 39636
rect 3011 39596 3056 39624
rect 3050 39584 3056 39596
rect 3108 39584 3114 39636
rect 3694 39584 3700 39636
rect 3752 39624 3758 39636
rect 3973 39627 4031 39633
rect 3973 39624 3985 39627
rect 3752 39596 3985 39624
rect 3752 39584 3758 39596
rect 3973 39593 3985 39596
rect 4019 39593 4031 39627
rect 3973 39587 4031 39593
rect 26234 39584 26240 39636
rect 26292 39624 26298 39636
rect 27157 39627 27215 39633
rect 27157 39624 27169 39627
rect 26292 39596 27169 39624
rect 26292 39584 26298 39596
rect 27157 39593 27169 39596
rect 27203 39593 27215 39627
rect 41414 39624 41420 39636
rect 41375 39596 41420 39624
rect 27157 39587 27215 39593
rect 41414 39584 41420 39596
rect 41472 39584 41478 39636
rect 48682 39584 48688 39636
rect 48740 39624 48746 39636
rect 48961 39627 49019 39633
rect 48961 39624 48973 39627
rect 48740 39596 48973 39624
rect 48740 39584 48746 39596
rect 48961 39593 48973 39596
rect 49007 39593 49019 39627
rect 48961 39587 49019 39593
rect 56134 39584 56140 39636
rect 56192 39624 56198 39636
rect 56413 39627 56471 39633
rect 56413 39624 56425 39627
rect 56192 39596 56425 39624
rect 56192 39584 56198 39596
rect 56413 39593 56425 39596
rect 56459 39593 56471 39627
rect 56413 39587 56471 39593
rect 8846 39488 8852 39500
rect 2148 39460 8852 39488
rect 1397 39423 1455 39429
rect 1397 39389 1409 39423
rect 1443 39420 1455 39423
rect 1486 39420 1492 39432
rect 1443 39392 1492 39420
rect 1443 39389 1455 39392
rect 1397 39383 1455 39389
rect 1486 39380 1492 39392
rect 1544 39380 1550 39432
rect 2148 39429 2176 39460
rect 8846 39448 8852 39460
rect 8904 39448 8910 39500
rect 18690 39448 18696 39500
rect 18748 39488 18754 39500
rect 19245 39491 19303 39497
rect 19245 39488 19257 39491
rect 18748 39460 19257 39488
rect 18748 39448 18754 39460
rect 19245 39457 19257 39460
rect 19291 39457 19303 39491
rect 19245 39451 19303 39457
rect 2133 39423 2191 39429
rect 2133 39389 2145 39423
rect 2179 39389 2191 39423
rect 2133 39383 2191 39389
rect 2869 39423 2927 39429
rect 2869 39389 2881 39423
rect 2915 39420 2927 39423
rect 3234 39420 3240 39432
rect 2915 39392 3240 39420
rect 2915 39389 2927 39392
rect 2869 39383 2927 39389
rect 3234 39380 3240 39392
rect 3292 39380 3298 39432
rect 3789 39423 3847 39429
rect 3789 39389 3801 39423
rect 3835 39420 3847 39423
rect 26970 39420 26976 39432
rect 3835 39392 4476 39420
rect 26931 39392 26976 39420
rect 3835 39389 3847 39392
rect 3789 39383 3847 39389
rect 4448 39296 4476 39392
rect 26970 39380 26976 39392
rect 27028 39380 27034 39432
rect 33686 39380 33692 39432
rect 33744 39420 33750 39432
rect 33781 39423 33839 39429
rect 33781 39420 33793 39423
rect 33744 39392 33793 39420
rect 33744 39380 33750 39392
rect 33781 39389 33793 39392
rect 33827 39389 33839 39423
rect 33781 39383 33839 39389
rect 55398 39380 55404 39432
rect 55456 39420 55462 39432
rect 56229 39423 56287 39429
rect 56229 39420 56241 39423
rect 55456 39392 56241 39420
rect 55456 39380 55462 39392
rect 56229 39389 56241 39392
rect 56275 39389 56287 39423
rect 56229 39383 56287 39389
rect 1578 39284 1584 39296
rect 1539 39256 1584 39284
rect 1578 39244 1584 39256
rect 1636 39244 1642 39296
rect 4430 39284 4436 39296
rect 4391 39256 4436 39284
rect 4430 39244 4436 39256
rect 4488 39244 4494 39296
rect 33965 39287 34023 39293
rect 33965 39253 33977 39287
rect 34011 39284 34023 39287
rect 34238 39284 34244 39296
rect 34011 39256 34244 39284
rect 34011 39253 34023 39256
rect 33965 39247 34023 39253
rect 34238 39244 34244 39256
rect 34296 39244 34302 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 4430 39040 4436 39092
rect 4488 39080 4494 39092
rect 4488 39052 26234 39080
rect 4488 39040 4494 39052
rect 26206 39012 26234 39052
rect 26970 39040 26976 39092
rect 27028 39080 27034 39092
rect 35069 39083 35127 39089
rect 35069 39080 35081 39083
rect 27028 39052 35081 39080
rect 27028 39040 27034 39052
rect 35069 39049 35081 39052
rect 35115 39049 35127 39083
rect 35069 39043 35127 39049
rect 35802 39012 35808 39024
rect 26206 38984 35808 39012
rect 35802 38972 35808 38984
rect 35860 38972 35866 39024
rect 1397 38947 1455 38953
rect 1397 38913 1409 38947
rect 1443 38944 1455 38947
rect 7190 38944 7196 38956
rect 1443 38916 7196 38944
rect 1443 38913 1455 38916
rect 1397 38907 1455 38913
rect 7190 38904 7196 38916
rect 7248 38904 7254 38956
rect 35253 38947 35311 38953
rect 35253 38913 35265 38947
rect 35299 38944 35311 38947
rect 35710 38944 35716 38956
rect 35299 38916 35716 38944
rect 35299 38913 35311 38916
rect 35253 38907 35311 38913
rect 35710 38904 35716 38916
rect 35768 38904 35774 38956
rect 1578 38740 1584 38752
rect 1539 38712 1584 38740
rect 1578 38700 1584 38712
rect 1636 38700 1642 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1581 38539 1639 38545
rect 1581 38505 1593 38539
rect 1627 38536 1639 38539
rect 2866 38536 2872 38548
rect 1627 38508 2872 38536
rect 1627 38505 1639 38508
rect 1581 38499 1639 38505
rect 2866 38496 2872 38508
rect 2924 38496 2930 38548
rect 1397 38335 1455 38341
rect 1397 38301 1409 38335
rect 1443 38332 1455 38335
rect 2406 38332 2412 38344
rect 1443 38304 2412 38332
rect 1443 38301 1455 38304
rect 1397 38295 1455 38301
rect 2406 38292 2412 38304
rect 2464 38292 2470 38344
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1397 37859 1455 37865
rect 1397 37825 1409 37859
rect 1443 37856 1455 37859
rect 1762 37856 1768 37868
rect 1443 37828 1768 37856
rect 1443 37825 1455 37828
rect 1397 37819 1455 37825
rect 1762 37816 1768 37828
rect 1820 37816 1826 37868
rect 1578 37652 1584 37664
rect 1539 37624 1584 37652
rect 1578 37612 1584 37624
rect 1636 37612 1642 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1397 36771 1455 36777
rect 1397 36737 1409 36771
rect 1443 36768 1455 36771
rect 1670 36768 1676 36780
rect 1443 36740 1676 36768
rect 1443 36737 1455 36740
rect 1397 36731 1455 36737
rect 1670 36728 1676 36740
rect 1728 36728 1734 36780
rect 1578 36632 1584 36644
rect 1539 36604 1584 36632
rect 1578 36592 1584 36604
rect 1636 36592 1642 36644
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1397 36159 1455 36165
rect 1397 36125 1409 36159
rect 1443 36156 1455 36159
rect 12802 36156 12808 36168
rect 1443 36128 12808 36156
rect 1443 36125 1455 36128
rect 1397 36119 1455 36125
rect 12802 36116 12808 36128
rect 12860 36116 12866 36168
rect 1578 36020 1584 36032
rect 1539 35992 1584 36020
rect 1578 35980 1584 35992
rect 1636 35980 1642 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1854 35000 1860 35012
rect 1815 34972 1860 35000
rect 1854 34960 1860 34972
rect 1912 34960 1918 35012
rect 1946 34932 1952 34944
rect 1907 34904 1952 34932
rect 1946 34892 1952 34904
rect 2004 34892 2010 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1578 34728 1584 34740
rect 1539 34700 1584 34728
rect 1578 34688 1584 34700
rect 1636 34688 1642 34740
rect 2133 34731 2191 34737
rect 2133 34697 2145 34731
rect 2179 34728 2191 34731
rect 5626 34728 5632 34740
rect 2179 34700 5632 34728
rect 2179 34697 2191 34700
rect 2133 34691 2191 34697
rect 5626 34688 5632 34700
rect 5684 34688 5690 34740
rect 1397 34595 1455 34601
rect 1397 34561 1409 34595
rect 1443 34561 1455 34595
rect 2314 34592 2320 34604
rect 2275 34564 2320 34592
rect 1397 34555 1455 34561
rect 1412 34524 1440 34555
rect 2314 34552 2320 34564
rect 2372 34552 2378 34604
rect 5718 34524 5724 34536
rect 1412 34496 5724 34524
rect 5718 34484 5724 34496
rect 5776 34484 5782 34536
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1397 33983 1455 33989
rect 1397 33949 1409 33983
rect 1443 33980 1455 33983
rect 13814 33980 13820 33992
rect 1443 33952 13820 33980
rect 1443 33949 1455 33952
rect 1397 33943 1455 33949
rect 13814 33940 13820 33952
rect 13872 33940 13878 33992
rect 1578 33844 1584 33856
rect 1539 33816 1584 33844
rect 1578 33804 1584 33816
rect 1636 33804 1642 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1854 33504 1860 33516
rect 1815 33476 1860 33504
rect 1854 33464 1860 33476
rect 1912 33464 1918 33516
rect 2866 33504 2872 33516
rect 2827 33476 2872 33504
rect 2866 33464 2872 33476
rect 2924 33464 2930 33516
rect 2038 33368 2044 33380
rect 1999 33340 2044 33368
rect 2038 33328 2044 33340
rect 2096 33328 2102 33380
rect 2685 33303 2743 33309
rect 2685 33269 2697 33303
rect 2731 33300 2743 33303
rect 5534 33300 5540 33312
rect 2731 33272 5540 33300
rect 2731 33269 2743 33272
rect 2685 33263 2743 33269
rect 5534 33260 5540 33272
rect 5592 33260 5598 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1397 32895 1455 32901
rect 1397 32861 1409 32895
rect 1443 32892 1455 32895
rect 10870 32892 10876 32904
rect 1443 32864 10876 32892
rect 1443 32861 1455 32864
rect 1397 32855 1455 32861
rect 10870 32852 10876 32864
rect 10928 32852 10934 32904
rect 1578 32756 1584 32768
rect 1539 32728 1584 32756
rect 1578 32716 1584 32728
rect 1636 32716 1642 32768
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1394 32416 1400 32428
rect 1355 32388 1400 32416
rect 1394 32376 1400 32388
rect 1452 32376 1458 32428
rect 1581 32215 1639 32221
rect 1581 32181 1593 32215
rect 1627 32212 1639 32215
rect 2222 32212 2228 32224
rect 1627 32184 2228 32212
rect 1627 32181 1639 32184
rect 1581 32175 1639 32181
rect 2222 32172 2228 32184
rect 2280 32172 2286 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 1397 31943 1455 31949
rect 1397 31909 1409 31943
rect 1443 31940 1455 31943
rect 4982 31940 4988 31952
rect 1443 31912 4988 31940
rect 1443 31909 1455 31912
rect 1397 31903 1455 31909
rect 4982 31900 4988 31912
rect 5040 31900 5046 31952
rect 1578 31804 1584 31816
rect 1539 31776 1584 31804
rect 1578 31764 1584 31776
rect 1636 31764 1642 31816
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 1854 31328 1860 31340
rect 1815 31300 1860 31328
rect 1854 31288 1860 31300
rect 1912 31288 1918 31340
rect 1670 31152 1676 31204
rect 1728 31192 1734 31204
rect 2314 31192 2320 31204
rect 1728 31164 2320 31192
rect 1728 31152 1734 31164
rect 2314 31152 2320 31164
rect 2372 31152 2378 31204
rect 2133 31127 2191 31133
rect 2133 31093 2145 31127
rect 2179 31124 2191 31127
rect 25314 31124 25320 31136
rect 2179 31096 25320 31124
rect 2179 31093 2191 31096
rect 2133 31087 2191 31093
rect 25314 31084 25320 31096
rect 25372 31084 25378 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 1578 30920 1584 30932
rect 1539 30892 1584 30920
rect 1578 30880 1584 30892
rect 1636 30880 1642 30932
rect 2133 30855 2191 30861
rect 2133 30821 2145 30855
rect 2179 30852 2191 30855
rect 4890 30852 4896 30864
rect 2179 30824 4896 30852
rect 2179 30821 2191 30824
rect 2133 30815 2191 30821
rect 4890 30812 4896 30824
rect 4948 30812 4954 30864
rect 1397 30719 1455 30725
rect 1397 30685 1409 30719
rect 1443 30716 1455 30719
rect 1486 30716 1492 30728
rect 1443 30688 1492 30716
rect 1443 30685 1455 30688
rect 1397 30679 1455 30685
rect 1486 30676 1492 30688
rect 1544 30676 1550 30728
rect 2317 30719 2375 30725
rect 2317 30685 2329 30719
rect 2363 30716 2375 30719
rect 2958 30716 2964 30728
rect 2363 30688 2774 30716
rect 2919 30688 2964 30716
rect 2363 30685 2375 30688
rect 2317 30679 2375 30685
rect 2746 30648 2774 30688
rect 2958 30676 2964 30688
rect 3016 30676 3022 30728
rect 4798 30716 4804 30728
rect 4759 30688 4804 30716
rect 4798 30676 4804 30688
rect 4856 30676 4862 30728
rect 2866 30648 2872 30660
rect 2746 30620 2872 30648
rect 2866 30608 2872 30620
rect 2924 30608 2930 30660
rect 2774 30540 2780 30592
rect 2832 30580 2838 30592
rect 4617 30583 4675 30589
rect 2832 30552 2877 30580
rect 2832 30540 2838 30552
rect 4617 30549 4629 30583
rect 4663 30580 4675 30583
rect 4706 30580 4712 30592
rect 4663 30552 4712 30580
rect 4663 30549 4675 30552
rect 4617 30543 4675 30549
rect 4706 30540 4712 30552
rect 4764 30540 4770 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 2774 30336 2780 30388
rect 2832 30376 2838 30388
rect 2832 30348 2877 30376
rect 2832 30336 2838 30348
rect 1394 30240 1400 30252
rect 1355 30212 1400 30240
rect 1394 30200 1400 30212
rect 1452 30200 1458 30252
rect 2682 30240 2688 30252
rect 2643 30212 2688 30240
rect 2682 30200 2688 30212
rect 2740 30200 2746 30252
rect 4706 30249 4712 30252
rect 4700 30240 4712 30249
rect 4667 30212 4712 30240
rect 4700 30203 4712 30212
rect 4706 30200 4712 30203
rect 4764 30200 4770 30252
rect 2958 30172 2964 30184
rect 2919 30144 2964 30172
rect 2958 30132 2964 30144
rect 3016 30132 3022 30184
rect 4062 30132 4068 30184
rect 4120 30172 4126 30184
rect 4433 30175 4491 30181
rect 4433 30172 4445 30175
rect 4120 30144 4445 30172
rect 4120 30132 4126 30144
rect 4433 30141 4445 30144
rect 4479 30141 4491 30175
rect 4433 30135 4491 30141
rect 1578 30036 1584 30048
rect 1539 30008 1584 30036
rect 1578 29996 1584 30008
rect 1636 29996 1642 30048
rect 2317 30039 2375 30045
rect 2317 30005 2329 30039
rect 2363 30036 2375 30039
rect 3602 30036 3608 30048
rect 2363 30008 3608 30036
rect 2363 30005 2375 30008
rect 2317 29999 2375 30005
rect 3602 29996 3608 30008
rect 3660 29996 3666 30048
rect 4614 29996 4620 30048
rect 4672 30036 4678 30048
rect 5813 30039 5871 30045
rect 5813 30036 5825 30039
rect 4672 30008 5825 30036
rect 4672 29996 4678 30008
rect 5813 30005 5825 30008
rect 5859 30005 5871 30039
rect 5813 29999 5871 30005
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 1394 29792 1400 29844
rect 1452 29832 1458 29844
rect 6822 29832 6828 29844
rect 1452 29804 6684 29832
rect 6783 29804 6828 29832
rect 1452 29792 1458 29804
rect 4249 29767 4307 29773
rect 4249 29733 4261 29767
rect 4295 29764 4307 29767
rect 4706 29764 4712 29776
rect 4295 29736 4712 29764
rect 4295 29733 4307 29736
rect 4249 29727 4307 29733
rect 4706 29724 4712 29736
rect 4764 29724 4770 29776
rect 6656 29764 6684 29804
rect 6822 29792 6828 29804
rect 6880 29792 6886 29844
rect 7193 29835 7251 29841
rect 7193 29801 7205 29835
rect 7239 29832 7251 29835
rect 7466 29832 7472 29844
rect 7239 29804 7472 29832
rect 7239 29801 7251 29804
rect 7193 29795 7251 29801
rect 7466 29792 7472 29804
rect 7524 29792 7530 29844
rect 6656 29736 12434 29764
rect 2958 29656 2964 29708
rect 3016 29696 3022 29708
rect 4798 29696 4804 29708
rect 3016 29668 4804 29696
rect 3016 29656 3022 29668
rect 4798 29656 4804 29668
rect 4856 29656 4862 29708
rect 12406 29696 12434 29736
rect 15102 29696 15108 29708
rect 12406 29668 15108 29696
rect 15102 29656 15108 29668
rect 15160 29656 15166 29708
rect 1857 29631 1915 29637
rect 1857 29597 1869 29631
rect 1903 29628 1915 29631
rect 4154 29628 4160 29640
rect 1903 29600 4160 29628
rect 1903 29597 1915 29600
rect 1857 29591 1915 29597
rect 4154 29588 4160 29600
rect 4212 29588 4218 29640
rect 4614 29628 4620 29640
rect 4575 29600 4620 29628
rect 4614 29588 4620 29600
rect 4672 29588 4678 29640
rect 4709 29631 4767 29637
rect 4709 29597 4721 29631
rect 4755 29628 4767 29631
rect 4982 29628 4988 29640
rect 4755 29600 4988 29628
rect 4755 29597 4767 29600
rect 4709 29591 4767 29597
rect 4982 29588 4988 29600
rect 5040 29588 5046 29640
rect 6917 29631 6975 29637
rect 6917 29628 6929 29631
rect 5736 29600 6929 29628
rect 2124 29563 2182 29569
rect 2124 29529 2136 29563
rect 2170 29560 2182 29563
rect 3418 29560 3424 29572
rect 2170 29532 3424 29560
rect 2170 29529 2182 29532
rect 2124 29523 2182 29529
rect 3418 29520 3424 29532
rect 3476 29520 3482 29572
rect 4632 29560 4660 29588
rect 5736 29560 5764 29600
rect 6917 29597 6929 29600
rect 6963 29597 6975 29631
rect 6917 29591 6975 29597
rect 7006 29588 7012 29640
rect 7064 29628 7070 29640
rect 7926 29628 7932 29640
rect 7064 29600 7109 29628
rect 7887 29600 7932 29628
rect 7064 29588 7070 29600
rect 7926 29588 7932 29600
rect 7984 29588 7990 29640
rect 4632 29532 5764 29560
rect 6733 29563 6791 29569
rect 6733 29529 6745 29563
rect 6779 29560 6791 29563
rect 7282 29560 7288 29572
rect 6779 29532 7288 29560
rect 6779 29529 6791 29532
rect 6733 29523 6791 29529
rect 7282 29520 7288 29532
rect 7340 29520 7346 29572
rect 2682 29452 2688 29504
rect 2740 29492 2746 29504
rect 3237 29495 3295 29501
rect 3237 29492 3249 29495
rect 2740 29464 3249 29492
rect 2740 29452 2746 29464
rect 3237 29461 3249 29464
rect 3283 29492 3295 29495
rect 6822 29492 6828 29504
rect 3283 29464 6828 29492
rect 3283 29461 3295 29464
rect 3237 29455 3295 29461
rect 6822 29452 6828 29464
rect 6880 29452 6886 29504
rect 7374 29452 7380 29504
rect 7432 29492 7438 29504
rect 7745 29495 7803 29501
rect 7745 29492 7757 29495
rect 7432 29464 7757 29492
rect 7432 29452 7438 29464
rect 7745 29461 7757 29464
rect 7791 29461 7803 29495
rect 7745 29455 7803 29461
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 3418 29288 3424 29300
rect 2700 29260 3280 29288
rect 3379 29260 3424 29288
rect 1854 29220 1860 29232
rect 1815 29192 1860 29220
rect 1854 29180 1860 29192
rect 1912 29180 1918 29232
rect 2700 29161 2728 29260
rect 3252 29220 3280 29260
rect 3418 29248 3424 29260
rect 3476 29248 3482 29300
rect 7282 29248 7288 29300
rect 7340 29288 7346 29300
rect 8205 29291 8263 29297
rect 8205 29288 8217 29291
rect 7340 29260 8217 29288
rect 7340 29248 7346 29260
rect 8205 29257 8217 29260
rect 8251 29257 8263 29291
rect 8205 29251 8263 29257
rect 17402 29220 17408 29232
rect 3252 29192 17408 29220
rect 17402 29180 17408 29192
rect 17460 29180 17466 29232
rect 2685 29155 2743 29161
rect 2685 29121 2697 29155
rect 2731 29121 2743 29155
rect 3602 29152 3608 29164
rect 3563 29124 3608 29152
rect 2685 29115 2743 29121
rect 3602 29112 3608 29124
rect 3660 29112 3666 29164
rect 4154 29112 4160 29164
rect 4212 29152 4218 29164
rect 4249 29155 4307 29161
rect 4249 29152 4261 29155
rect 4212 29124 4261 29152
rect 4212 29112 4218 29124
rect 4249 29121 4261 29124
rect 4295 29121 4307 29155
rect 4249 29115 4307 29121
rect 7092 29155 7150 29161
rect 7092 29121 7104 29155
rect 7138 29152 7150 29155
rect 7374 29152 7380 29164
rect 7138 29124 7380 29152
rect 7138 29121 7150 29124
rect 7092 29115 7150 29121
rect 7374 29112 7380 29124
rect 7432 29112 7438 29164
rect 3970 29044 3976 29096
rect 4028 29084 4034 29096
rect 5442 29084 5448 29096
rect 4028 29056 5448 29084
rect 4028 29044 4034 29056
rect 5442 29044 5448 29056
rect 5500 29084 5506 29096
rect 6825 29087 6883 29093
rect 6825 29084 6837 29087
rect 5500 29056 6837 29084
rect 5500 29044 5506 29056
rect 6825 29053 6837 29056
rect 6871 29053 6883 29087
rect 6825 29047 6883 29053
rect 2133 29019 2191 29025
rect 2133 28985 2145 29019
rect 2179 29016 2191 29019
rect 2590 29016 2596 29028
rect 2179 28988 2596 29016
rect 2179 28985 2191 28988
rect 2133 28979 2191 28985
rect 2590 28976 2596 28988
rect 2648 28976 2654 29028
rect 2866 29016 2872 29028
rect 2827 28988 2872 29016
rect 2866 28976 2872 28988
rect 2924 28976 2930 29028
rect 4065 29019 4123 29025
rect 4065 28985 4077 29019
rect 4111 29016 4123 29019
rect 4614 29016 4620 29028
rect 4111 28988 4620 29016
rect 4111 28985 4123 28988
rect 4065 28979 4123 28985
rect 4614 28976 4620 28988
rect 4672 28976 4678 29028
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 3881 28747 3939 28753
rect 3881 28713 3893 28747
rect 3927 28744 3939 28747
rect 4062 28744 4068 28756
rect 3927 28716 4068 28744
rect 3927 28713 3939 28716
rect 3881 28707 3939 28713
rect 4062 28704 4068 28716
rect 4120 28704 4126 28756
rect 6917 28747 6975 28753
rect 6917 28713 6929 28747
rect 6963 28744 6975 28747
rect 7926 28744 7932 28756
rect 6963 28716 7932 28744
rect 6963 28713 6975 28716
rect 6917 28707 6975 28713
rect 7926 28704 7932 28716
rect 7984 28704 7990 28756
rect 15102 28704 15108 28756
rect 15160 28744 15166 28756
rect 15473 28747 15531 28753
rect 15473 28744 15485 28747
rect 15160 28716 15485 28744
rect 15160 28704 15166 28716
rect 15473 28713 15485 28716
rect 15519 28713 15531 28747
rect 15473 28707 15531 28713
rect 4525 28611 4583 28617
rect 4525 28577 4537 28611
rect 4571 28608 4583 28611
rect 4798 28608 4804 28620
rect 4571 28580 4804 28608
rect 4571 28577 4583 28580
rect 4525 28571 4583 28577
rect 4798 28568 4804 28580
rect 4856 28568 4862 28620
rect 5534 28568 5540 28620
rect 5592 28608 5598 28620
rect 7377 28611 7435 28617
rect 7377 28608 7389 28611
rect 5592 28580 7389 28608
rect 5592 28568 5598 28580
rect 7377 28577 7389 28580
rect 7423 28577 7435 28611
rect 7558 28608 7564 28620
rect 7519 28580 7564 28608
rect 7377 28571 7435 28577
rect 7558 28568 7564 28580
rect 7616 28568 7622 28620
rect 4341 28543 4399 28549
rect 4341 28509 4353 28543
rect 4387 28540 4399 28543
rect 4890 28540 4896 28552
rect 4387 28512 4896 28540
rect 4387 28509 4399 28512
rect 4341 28503 4399 28509
rect 4890 28500 4896 28512
rect 4948 28500 4954 28552
rect 7282 28540 7288 28552
rect 7243 28512 7288 28540
rect 7282 28500 7288 28512
rect 7340 28500 7346 28552
rect 10689 28543 10747 28549
rect 10689 28509 10701 28543
rect 10735 28509 10747 28543
rect 10870 28540 10876 28552
rect 10831 28512 10876 28540
rect 10689 28503 10747 28509
rect 1854 28472 1860 28484
rect 1815 28444 1860 28472
rect 1854 28432 1860 28444
rect 1912 28432 1918 28484
rect 10704 28472 10732 28503
rect 10870 28500 10876 28512
rect 10928 28500 10934 28552
rect 10962 28500 10968 28552
rect 11020 28540 11026 28552
rect 11020 28512 11065 28540
rect 11020 28500 11026 28512
rect 12526 28500 12532 28552
rect 12584 28540 12590 28552
rect 14093 28543 14151 28549
rect 14093 28540 14105 28543
rect 12584 28512 14105 28540
rect 12584 28500 12590 28512
rect 14093 28509 14105 28512
rect 14139 28540 14151 28543
rect 16669 28543 16727 28549
rect 16669 28540 16681 28543
rect 14139 28512 16681 28540
rect 14139 28509 14151 28512
rect 14093 28503 14151 28509
rect 16669 28509 16681 28512
rect 16715 28509 16727 28543
rect 16669 28503 16727 28509
rect 13446 28472 13452 28484
rect 10704 28444 13452 28472
rect 13446 28432 13452 28444
rect 13504 28432 13510 28484
rect 14360 28475 14418 28481
rect 14360 28441 14372 28475
rect 14406 28472 14418 28475
rect 14642 28472 14648 28484
rect 14406 28444 14648 28472
rect 14406 28441 14418 28444
rect 14360 28435 14418 28441
rect 14642 28432 14648 28444
rect 14700 28432 14706 28484
rect 16936 28475 16994 28481
rect 16936 28441 16948 28475
rect 16982 28472 16994 28475
rect 17034 28472 17040 28484
rect 16982 28444 17040 28472
rect 16982 28441 16994 28444
rect 16936 28435 16994 28441
rect 17034 28432 17040 28444
rect 17092 28432 17098 28484
rect 2130 28404 2136 28416
rect 2091 28376 2136 28404
rect 2130 28364 2136 28376
rect 2188 28364 2194 28416
rect 4249 28407 4307 28413
rect 4249 28373 4261 28407
rect 4295 28404 4307 28407
rect 7006 28404 7012 28416
rect 4295 28376 7012 28404
rect 4295 28373 4307 28376
rect 4249 28367 4307 28373
rect 7006 28364 7012 28376
rect 7064 28364 7070 28416
rect 10502 28404 10508 28416
rect 10463 28376 10508 28404
rect 10502 28364 10508 28376
rect 10560 28364 10566 28416
rect 17402 28364 17408 28416
rect 17460 28404 17466 28416
rect 18049 28407 18107 28413
rect 18049 28404 18061 28407
rect 17460 28376 18061 28404
rect 17460 28364 17466 28376
rect 18049 28373 18061 28376
rect 18095 28373 18107 28407
rect 18049 28367 18107 28373
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 2130 28160 2136 28212
rect 2188 28200 2194 28212
rect 13814 28200 13820 28212
rect 2188 28172 12434 28200
rect 13775 28172 13820 28200
rect 2188 28160 2194 28172
rect 4424 28135 4482 28141
rect 1412 28104 4384 28132
rect 1412 28073 1440 28104
rect 1397 28067 1455 28073
rect 1397 28033 1409 28067
rect 1443 28033 1455 28067
rect 2406 28064 2412 28076
rect 2367 28036 2412 28064
rect 1397 28027 1455 28033
rect 2406 28024 2412 28036
rect 2464 28024 2470 28076
rect 3050 28064 3056 28076
rect 3011 28036 3056 28064
rect 3050 28024 3056 28036
rect 3108 28024 3114 28076
rect 3970 28024 3976 28076
rect 4028 28064 4034 28076
rect 4157 28067 4215 28073
rect 4157 28064 4169 28067
rect 4028 28036 4169 28064
rect 4028 28024 4034 28036
rect 4157 28033 4169 28036
rect 4203 28033 4215 28067
rect 4356 28064 4384 28104
rect 4424 28101 4436 28135
rect 4470 28132 4482 28135
rect 4614 28132 4620 28144
rect 4470 28104 4620 28132
rect 4470 28101 4482 28104
rect 4424 28095 4482 28101
rect 4614 28092 4620 28104
rect 4672 28092 4678 28144
rect 9852 28135 9910 28141
rect 9852 28101 9864 28135
rect 9898 28132 9910 28135
rect 10502 28132 10508 28144
rect 9898 28104 10508 28132
rect 9898 28101 9910 28104
rect 9852 28095 9910 28101
rect 10502 28092 10508 28104
rect 10560 28092 10566 28144
rect 12406 28132 12434 28172
rect 13814 28160 13820 28172
rect 13872 28160 13878 28212
rect 14642 28200 14648 28212
rect 14603 28172 14648 28200
rect 14642 28160 14648 28172
rect 14700 28160 14706 28212
rect 15013 28203 15071 28209
rect 15013 28169 15025 28203
rect 15059 28200 15071 28203
rect 15102 28200 15108 28212
rect 15059 28172 15108 28200
rect 15059 28169 15071 28172
rect 15013 28163 15071 28169
rect 15102 28160 15108 28172
rect 15160 28160 15166 28212
rect 17034 28200 17040 28212
rect 16995 28172 17040 28200
rect 17034 28160 17040 28172
rect 17092 28160 17098 28212
rect 17402 28200 17408 28212
rect 17363 28172 17408 28200
rect 17402 28160 17408 28172
rect 17460 28160 17466 28212
rect 12406 28104 22094 28132
rect 6822 28064 6828 28076
rect 4356 28036 5212 28064
rect 6783 28036 6828 28064
rect 4157 28027 4215 28033
rect 5184 27996 5212 28036
rect 6822 28024 6828 28036
rect 6880 28024 6886 28076
rect 9585 28067 9643 28073
rect 9585 28033 9597 28067
rect 9631 28064 9643 28067
rect 9674 28064 9680 28076
rect 9631 28036 9680 28064
rect 9631 28033 9643 28036
rect 9585 28027 9643 28033
rect 9674 28024 9680 28036
rect 9732 28024 9738 28076
rect 12437 28067 12495 28073
rect 12437 28033 12449 28067
rect 12483 28064 12495 28067
rect 12526 28064 12532 28076
rect 12483 28036 12532 28064
rect 12483 28033 12495 28036
rect 12437 28027 12495 28033
rect 12526 28024 12532 28036
rect 12584 28024 12590 28076
rect 12710 28073 12716 28076
rect 12704 28027 12716 28073
rect 12768 28064 12774 28076
rect 14829 28067 14887 28073
rect 12768 28036 12804 28064
rect 12710 28024 12716 28027
rect 12768 28024 12774 28036
rect 14829 28033 14841 28067
rect 14875 28033 14887 28067
rect 14829 28027 14887 28033
rect 15105 28067 15163 28073
rect 15105 28033 15117 28067
rect 15151 28064 15163 28067
rect 16942 28064 16948 28076
rect 15151 28036 16948 28064
rect 15151 28033 15163 28036
rect 15105 28027 15163 28033
rect 14844 27996 14872 28027
rect 16942 28024 16948 28036
rect 17000 28024 17006 28076
rect 17218 28064 17224 28076
rect 17179 28036 17224 28064
rect 17218 28024 17224 28036
rect 17276 28024 17282 28076
rect 17497 28067 17555 28073
rect 17497 28033 17509 28067
rect 17543 28033 17555 28067
rect 17497 28027 17555 28033
rect 16758 27996 16764 28008
rect 5184 27968 7788 27996
rect 14844 27968 16764 27996
rect 5537 27931 5595 27937
rect 5537 27897 5549 27931
rect 5583 27928 5595 27931
rect 7006 27928 7012 27940
rect 5583 27900 7012 27928
rect 5583 27897 5595 27900
rect 5537 27891 5595 27897
rect 7006 27888 7012 27900
rect 7064 27928 7070 27940
rect 7650 27928 7656 27940
rect 7064 27900 7656 27928
rect 7064 27888 7070 27900
rect 7650 27888 7656 27900
rect 7708 27888 7714 27940
rect 1578 27860 1584 27872
rect 1539 27832 1584 27860
rect 1578 27820 1584 27832
rect 1636 27820 1642 27872
rect 2130 27820 2136 27872
rect 2188 27860 2194 27872
rect 2225 27863 2283 27869
rect 2225 27860 2237 27863
rect 2188 27832 2237 27860
rect 2188 27820 2194 27832
rect 2225 27829 2237 27832
rect 2271 27829 2283 27863
rect 2866 27860 2872 27872
rect 2827 27832 2872 27860
rect 2225 27823 2283 27829
rect 2866 27820 2872 27832
rect 2924 27820 2930 27872
rect 6638 27860 6644 27872
rect 6599 27832 6644 27860
rect 6638 27820 6644 27832
rect 6696 27820 6702 27872
rect 7760 27860 7788 27968
rect 16758 27956 16764 27968
rect 16816 27956 16822 28008
rect 16960 27996 16988 28024
rect 17512 27996 17540 28027
rect 16960 27968 17540 27996
rect 22066 27996 22094 28104
rect 25498 27996 25504 28008
rect 22066 27968 25504 27996
rect 25498 27956 25504 27968
rect 25556 27956 25562 28008
rect 10870 27888 10876 27940
rect 10928 27928 10934 27940
rect 10965 27931 11023 27937
rect 10965 27928 10977 27931
rect 10928 27900 10977 27928
rect 10928 27888 10934 27900
rect 10965 27897 10977 27900
rect 11011 27897 11023 27931
rect 10965 27891 11023 27897
rect 17954 27860 17960 27872
rect 7760 27832 17960 27860
rect 17954 27820 17960 27832
rect 18012 27820 18018 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 6733 27659 6791 27665
rect 6733 27625 6745 27659
rect 6779 27656 6791 27659
rect 6822 27656 6828 27668
rect 6779 27628 6828 27656
rect 6779 27625 6791 27628
rect 6733 27619 6791 27625
rect 6822 27616 6828 27628
rect 6880 27616 6886 27668
rect 9674 27616 9680 27668
rect 9732 27656 9738 27668
rect 12618 27656 12624 27668
rect 9732 27628 12624 27656
rect 9732 27616 9738 27628
rect 12618 27616 12624 27628
rect 12676 27616 12682 27668
rect 12710 27616 12716 27668
rect 12768 27656 12774 27668
rect 12897 27659 12955 27665
rect 12897 27656 12909 27659
rect 12768 27628 12909 27656
rect 12768 27616 12774 27628
rect 12897 27625 12909 27628
rect 12943 27625 12955 27659
rect 12897 27619 12955 27625
rect 5626 27480 5632 27532
rect 5684 27520 5690 27532
rect 7193 27523 7251 27529
rect 7193 27520 7205 27523
rect 5684 27492 7205 27520
rect 5684 27480 5690 27492
rect 7193 27489 7205 27492
rect 7239 27489 7251 27523
rect 7193 27483 7251 27489
rect 7377 27523 7435 27529
rect 7377 27489 7389 27523
rect 7423 27520 7435 27523
rect 7558 27520 7564 27532
rect 7423 27492 7564 27520
rect 7423 27489 7435 27492
rect 7377 27483 7435 27489
rect 7558 27480 7564 27492
rect 7616 27520 7622 27532
rect 8110 27520 8116 27532
rect 7616 27492 8116 27520
rect 7616 27480 7622 27492
rect 8110 27480 8116 27492
rect 8168 27480 8174 27532
rect 9674 27520 9680 27532
rect 9635 27492 9680 27520
rect 9674 27480 9680 27492
rect 9732 27480 9738 27532
rect 13906 27520 13912 27532
rect 13096 27492 13912 27520
rect 1854 27452 1860 27464
rect 1815 27424 1860 27452
rect 1854 27412 1860 27424
rect 1912 27412 1918 27464
rect 2130 27461 2136 27464
rect 2124 27452 2136 27461
rect 2091 27424 2136 27452
rect 2124 27415 2136 27424
rect 2130 27412 2136 27415
rect 2188 27412 2194 27464
rect 13096 27461 13124 27492
rect 13906 27480 13912 27492
rect 13964 27480 13970 27532
rect 13081 27455 13139 27461
rect 13081 27421 13093 27455
rect 13127 27421 13139 27455
rect 13357 27455 13415 27461
rect 13357 27452 13369 27455
rect 13081 27415 13139 27421
rect 13188 27424 13369 27452
rect 2958 27344 2964 27396
rect 3016 27384 3022 27396
rect 4798 27384 4804 27396
rect 3016 27356 4804 27384
rect 3016 27344 3022 27356
rect 4798 27344 4804 27356
rect 4856 27344 4862 27396
rect 5718 27344 5724 27396
rect 5776 27384 5782 27396
rect 9944 27387 10002 27393
rect 5776 27356 9444 27384
rect 5776 27344 5782 27356
rect 1486 27276 1492 27328
rect 1544 27316 1550 27328
rect 3142 27316 3148 27328
rect 1544 27288 3148 27316
rect 1544 27276 1550 27288
rect 3142 27276 3148 27288
rect 3200 27276 3206 27328
rect 3237 27319 3295 27325
rect 3237 27285 3249 27319
rect 3283 27316 3295 27319
rect 3786 27316 3792 27328
rect 3283 27288 3792 27316
rect 3283 27285 3295 27288
rect 3237 27279 3295 27285
rect 3786 27276 3792 27288
rect 3844 27276 3850 27328
rect 7006 27276 7012 27328
rect 7064 27316 7070 27328
rect 7101 27319 7159 27325
rect 7101 27316 7113 27319
rect 7064 27288 7113 27316
rect 7064 27276 7070 27288
rect 7101 27285 7113 27288
rect 7147 27285 7159 27319
rect 9416 27316 9444 27356
rect 9944 27353 9956 27387
rect 9990 27384 10002 27387
rect 10502 27384 10508 27396
rect 9990 27356 10508 27384
rect 9990 27353 10002 27356
rect 9944 27347 10002 27353
rect 10502 27344 10508 27356
rect 10560 27344 10566 27396
rect 10962 27344 10968 27396
rect 11020 27384 11026 27396
rect 12894 27384 12900 27396
rect 11020 27356 12900 27384
rect 11020 27344 11026 27356
rect 12894 27344 12900 27356
rect 12952 27384 12958 27396
rect 13188 27384 13216 27424
rect 13357 27421 13369 27424
rect 13403 27421 13415 27455
rect 13357 27415 13415 27421
rect 12952 27356 13216 27384
rect 13265 27387 13323 27393
rect 12952 27344 12958 27356
rect 13265 27353 13277 27387
rect 13311 27384 13323 27387
rect 13814 27384 13820 27396
rect 13311 27356 13820 27384
rect 13311 27353 13323 27356
rect 13265 27347 13323 27353
rect 13814 27344 13820 27356
rect 13872 27344 13878 27396
rect 10870 27316 10876 27328
rect 9416 27288 10876 27316
rect 7101 27279 7159 27285
rect 10870 27276 10876 27288
rect 10928 27316 10934 27328
rect 11057 27319 11115 27325
rect 11057 27316 11069 27319
rect 10928 27288 11069 27316
rect 10928 27276 10934 27288
rect 11057 27285 11069 27288
rect 11103 27285 11115 27319
rect 11057 27279 11115 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 2317 27115 2375 27121
rect 2317 27081 2329 27115
rect 2363 27112 2375 27115
rect 2406 27112 2412 27124
rect 2363 27084 2412 27112
rect 2363 27081 2375 27084
rect 2317 27075 2375 27081
rect 2406 27072 2412 27084
rect 2464 27072 2470 27124
rect 2777 27115 2835 27121
rect 2777 27081 2789 27115
rect 2823 27112 2835 27115
rect 2866 27112 2872 27124
rect 2823 27084 2872 27112
rect 2823 27081 2835 27084
rect 2777 27075 2835 27081
rect 2866 27072 2872 27084
rect 2924 27072 2930 27124
rect 3142 27072 3148 27124
rect 3200 27112 3206 27124
rect 3200 27084 6776 27112
rect 3200 27072 3206 27084
rect 1486 27044 1492 27056
rect 1447 27016 1492 27044
rect 1486 27004 1492 27016
rect 1544 27004 1550 27056
rect 2685 27047 2743 27053
rect 2685 27013 2697 27047
rect 2731 27044 2743 27047
rect 3786 27044 3792 27056
rect 2731 27016 3792 27044
rect 2731 27013 2743 27016
rect 2685 27007 2743 27013
rect 3786 27004 3792 27016
rect 3844 27004 3850 27056
rect 6638 27053 6644 27056
rect 6632 27044 6644 27053
rect 6599 27016 6644 27044
rect 6632 27007 6644 27016
rect 6638 27004 6644 27007
rect 6696 27004 6702 27056
rect 6748 27044 6776 27084
rect 7006 27072 7012 27124
rect 7064 27112 7070 27124
rect 7745 27115 7803 27121
rect 7745 27112 7757 27115
rect 7064 27084 7757 27112
rect 7064 27072 7070 27084
rect 7745 27081 7757 27084
rect 7791 27081 7803 27115
rect 10502 27112 10508 27124
rect 10463 27084 10508 27112
rect 7745 27075 7803 27081
rect 10502 27072 10508 27084
rect 10560 27072 10566 27124
rect 10870 27112 10876 27124
rect 10831 27084 10876 27112
rect 10870 27072 10876 27084
rect 10928 27072 10934 27124
rect 16574 27044 16580 27056
rect 6748 27016 16580 27044
rect 16574 27004 16580 27016
rect 16632 27044 16638 27056
rect 17037 27047 17095 27053
rect 17037 27044 17049 27047
rect 16632 27016 17049 27044
rect 16632 27004 16638 27016
rect 17037 27013 17049 27016
rect 17083 27013 17095 27047
rect 17037 27007 17095 27013
rect 3694 26976 3700 26988
rect 3655 26948 3700 26976
rect 3694 26936 3700 26948
rect 3752 26936 3758 26988
rect 10686 26976 10692 26988
rect 3804 26948 7420 26976
rect 10647 26948 10692 26976
rect 2958 26908 2964 26920
rect 2919 26880 2964 26908
rect 2958 26868 2964 26880
rect 3016 26868 3022 26920
rect 3050 26868 3056 26920
rect 3108 26908 3114 26920
rect 3804 26908 3832 26948
rect 3108 26880 3832 26908
rect 3108 26868 3114 26880
rect 5442 26868 5448 26920
rect 5500 26908 5506 26920
rect 5902 26908 5908 26920
rect 5500 26880 5908 26908
rect 5500 26868 5506 26880
rect 5902 26868 5908 26880
rect 5960 26908 5966 26920
rect 6365 26911 6423 26917
rect 6365 26908 6377 26911
rect 5960 26880 6377 26908
rect 5960 26868 5966 26880
rect 6365 26877 6377 26880
rect 6411 26877 6423 26911
rect 7392 26908 7420 26948
rect 10686 26936 10692 26948
rect 10744 26936 10750 26988
rect 10962 26936 10968 26988
rect 11020 26976 11026 26988
rect 11020 26948 11065 26976
rect 11020 26936 11026 26948
rect 15838 26936 15844 26988
rect 15896 26976 15902 26988
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 15896 26948 16865 26976
rect 15896 26936 15902 26948
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 16942 26936 16948 26988
rect 17000 26976 17006 26988
rect 17129 26979 17187 26985
rect 17129 26976 17141 26979
rect 17000 26948 17141 26976
rect 17000 26936 17006 26948
rect 17129 26945 17141 26948
rect 17175 26976 17187 26979
rect 17770 26976 17776 26988
rect 17175 26948 17776 26976
rect 17175 26945 17187 26948
rect 17129 26939 17187 26945
rect 17770 26936 17776 26948
rect 17828 26936 17834 26988
rect 17310 26908 17316 26920
rect 7392 26880 17316 26908
rect 6365 26871 6423 26877
rect 17310 26868 17316 26880
rect 17368 26868 17374 26920
rect 1765 26843 1823 26849
rect 1765 26809 1777 26843
rect 1811 26840 1823 26843
rect 24486 26840 24492 26852
rect 1811 26812 6408 26840
rect 1811 26809 1823 26812
rect 1765 26803 1823 26809
rect 3510 26772 3516 26784
rect 3471 26744 3516 26772
rect 3510 26732 3516 26744
rect 3568 26732 3574 26784
rect 6380 26772 6408 26812
rect 7300 26812 24492 26840
rect 7300 26772 7328 26812
rect 24486 26800 24492 26812
rect 24544 26800 24550 26852
rect 6380 26744 7328 26772
rect 10686 26732 10692 26784
rect 10744 26772 10750 26784
rect 13722 26772 13728 26784
rect 10744 26744 13728 26772
rect 10744 26732 10750 26744
rect 13722 26732 13728 26744
rect 13780 26732 13786 26784
rect 16666 26772 16672 26784
rect 16627 26744 16672 26772
rect 16666 26732 16672 26744
rect 16724 26732 16730 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 1412 26540 3372 26568
rect 1412 26373 1440 26540
rect 3053 26503 3111 26509
rect 3053 26469 3065 26503
rect 3099 26469 3111 26503
rect 3344 26500 3372 26540
rect 3418 26528 3424 26580
rect 3476 26568 3482 26580
rect 5169 26571 5227 26577
rect 5169 26568 5181 26571
rect 3476 26540 5181 26568
rect 3476 26528 3482 26540
rect 5169 26537 5181 26540
rect 5215 26537 5227 26571
rect 5169 26531 5227 26537
rect 16574 26528 16580 26580
rect 16632 26568 16638 26580
rect 16669 26571 16727 26577
rect 16669 26568 16681 26571
rect 16632 26540 16681 26568
rect 16632 26528 16638 26540
rect 16669 26537 16681 26540
rect 16715 26537 16727 26571
rect 16669 26531 16727 26537
rect 18046 26528 18052 26580
rect 18104 26568 18110 26580
rect 18509 26571 18567 26577
rect 18509 26568 18521 26571
rect 18104 26540 18521 26568
rect 18104 26528 18110 26540
rect 18509 26537 18521 26540
rect 18555 26537 18567 26571
rect 18509 26531 18567 26537
rect 3694 26500 3700 26512
rect 3344 26472 3700 26500
rect 3053 26463 3111 26469
rect 3068 26432 3096 26463
rect 3694 26460 3700 26472
rect 3752 26460 3758 26512
rect 3068 26404 3924 26432
rect 1397 26367 1455 26373
rect 1397 26333 1409 26367
rect 1443 26333 1455 26367
rect 1397 26327 1455 26333
rect 2133 26367 2191 26373
rect 2133 26333 2145 26367
rect 2179 26364 2191 26367
rect 3050 26364 3056 26376
rect 2179 26336 3056 26364
rect 2179 26333 2191 26336
rect 2133 26327 2191 26333
rect 3050 26324 3056 26336
rect 3108 26324 3114 26376
rect 3234 26364 3240 26376
rect 3195 26336 3240 26364
rect 3234 26324 3240 26336
rect 3292 26324 3298 26376
rect 3789 26367 3847 26373
rect 3789 26333 3801 26367
rect 3835 26333 3847 26367
rect 3896 26364 3924 26404
rect 4045 26367 4103 26373
rect 4045 26364 4057 26367
rect 3896 26336 4057 26364
rect 3789 26327 3847 26333
rect 4045 26333 4057 26336
rect 4091 26333 4103 26367
rect 15289 26367 15347 26373
rect 15289 26364 15301 26367
rect 4045 26327 4103 26333
rect 15212 26336 15301 26364
rect 1854 26256 1860 26308
rect 1912 26296 1918 26308
rect 3804 26296 3832 26327
rect 15102 26296 15108 26308
rect 1912 26268 3832 26296
rect 3896 26268 15108 26296
rect 1912 26256 1918 26268
rect 1578 26228 1584 26240
rect 1539 26200 1584 26228
rect 1578 26188 1584 26200
rect 1636 26188 1642 26240
rect 2314 26228 2320 26240
rect 2275 26200 2320 26228
rect 2314 26188 2320 26200
rect 2372 26188 2378 26240
rect 3694 26188 3700 26240
rect 3752 26228 3758 26240
rect 3896 26228 3924 26268
rect 15102 26256 15108 26268
rect 15160 26256 15166 26308
rect 15212 26296 15240 26336
rect 15289 26333 15301 26336
rect 15335 26333 15347 26367
rect 15289 26327 15347 26333
rect 15556 26367 15614 26373
rect 15556 26333 15568 26367
rect 15602 26364 15614 26367
rect 16666 26364 16672 26376
rect 15602 26336 16672 26364
rect 15602 26333 15614 26336
rect 15556 26327 15614 26333
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 17129 26367 17187 26373
rect 17129 26333 17141 26367
rect 17175 26333 17187 26367
rect 17129 26327 17187 26333
rect 17144 26296 17172 26327
rect 17402 26305 17408 26308
rect 15212 26268 17172 26296
rect 3752 26200 3924 26228
rect 3752 26188 3758 26200
rect 13630 26188 13636 26240
rect 13688 26228 13694 26240
rect 15212 26228 15240 26268
rect 17396 26259 17408 26305
rect 17460 26296 17466 26308
rect 17460 26268 17496 26296
rect 17402 26256 17408 26259
rect 17460 26256 17466 26268
rect 13688 26200 15240 26228
rect 13688 26188 13694 26200
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 3053 26027 3111 26033
rect 3053 25993 3065 26027
rect 3099 26024 3111 26027
rect 3234 26024 3240 26036
rect 3099 25996 3240 26024
rect 3099 25993 3111 25996
rect 3053 25987 3111 25993
rect 3234 25984 3240 25996
rect 3292 25984 3298 26036
rect 3510 26024 3516 26036
rect 3471 25996 3516 26024
rect 3510 25984 3516 25996
rect 3568 25984 3574 26036
rect 8757 26027 8815 26033
rect 8757 26024 8769 26027
rect 4356 25996 8769 26024
rect 1670 25916 1676 25968
rect 1728 25956 1734 25968
rect 3418 25956 3424 25968
rect 1728 25928 2774 25956
rect 3379 25928 3424 25956
rect 1728 25916 1734 25928
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25848 1458 25900
rect 2314 25888 2320 25900
rect 2275 25860 2320 25888
rect 2314 25848 2320 25860
rect 2372 25848 2378 25900
rect 2746 25888 2774 25928
rect 3418 25916 3424 25928
rect 3476 25916 3482 25968
rect 4356 25888 4384 25996
rect 8757 25993 8769 25996
rect 8803 26024 8815 26027
rect 9306 26024 9312 26036
rect 8803 25996 9312 26024
rect 8803 25993 8815 25996
rect 8757 25987 8815 25993
rect 9306 25984 9312 25996
rect 9364 25984 9370 26036
rect 12802 25984 12808 26036
rect 12860 26024 12866 26036
rect 13909 26027 13967 26033
rect 13909 26024 13921 26027
rect 12860 25996 13921 26024
rect 12860 25984 12866 25996
rect 13909 25993 13921 25996
rect 13955 25993 13967 26027
rect 13909 25987 13967 25993
rect 17313 26027 17371 26033
rect 17313 25993 17325 26027
rect 17359 26024 17371 26027
rect 17402 26024 17408 26036
rect 17359 25996 17408 26024
rect 17359 25993 17371 25996
rect 17313 25987 17371 25993
rect 17402 25984 17408 25996
rect 17460 25984 17466 26036
rect 17681 26027 17739 26033
rect 17681 25993 17693 26027
rect 17727 26024 17739 26027
rect 17954 26024 17960 26036
rect 17727 25996 17960 26024
rect 17727 25993 17739 25996
rect 17681 25987 17739 25993
rect 17954 25984 17960 25996
rect 18012 25984 18018 26036
rect 4617 25959 4675 25965
rect 4617 25925 4629 25959
rect 4663 25956 4675 25959
rect 4798 25956 4804 25968
rect 4663 25928 4804 25956
rect 4663 25925 4675 25928
rect 4617 25919 4675 25925
rect 4798 25916 4804 25928
rect 4856 25916 4862 25968
rect 9674 25956 9680 25968
rect 7392 25928 9680 25956
rect 2746 25860 4384 25888
rect 4433 25891 4491 25897
rect 4433 25857 4445 25891
rect 4479 25888 4491 25891
rect 5534 25888 5540 25900
rect 4479 25860 5540 25888
rect 4479 25857 4491 25860
rect 4433 25851 4491 25857
rect 5534 25848 5540 25860
rect 5592 25848 5598 25900
rect 5902 25848 5908 25900
rect 5960 25888 5966 25900
rect 7392 25897 7420 25928
rect 7377 25891 7435 25897
rect 7377 25888 7389 25891
rect 5960 25860 7389 25888
rect 5960 25848 5966 25860
rect 7377 25857 7389 25860
rect 7423 25857 7435 25891
rect 7377 25851 7435 25857
rect 7644 25891 7702 25897
rect 7644 25857 7656 25891
rect 7690 25888 7702 25891
rect 9490 25888 9496 25900
rect 7690 25860 9496 25888
rect 7690 25857 7702 25860
rect 7644 25851 7702 25857
rect 9490 25848 9496 25860
rect 9548 25848 9554 25900
rect 9600 25897 9628 25928
rect 9674 25916 9680 25928
rect 9732 25916 9738 25968
rect 13630 25956 13636 25968
rect 12636 25928 13636 25956
rect 12636 25900 12664 25928
rect 13630 25916 13636 25928
rect 13688 25956 13694 25968
rect 13688 25928 13768 25956
rect 13688 25916 13694 25928
rect 9585 25891 9643 25897
rect 9585 25857 9597 25891
rect 9631 25857 9643 25891
rect 9585 25851 9643 25857
rect 9852 25891 9910 25897
rect 9852 25857 9864 25891
rect 9898 25888 9910 25891
rect 10870 25888 10876 25900
rect 9898 25860 10876 25888
rect 9898 25857 9910 25860
rect 9852 25851 9910 25857
rect 10870 25848 10876 25860
rect 10928 25848 10934 25900
rect 12529 25891 12587 25897
rect 12529 25857 12541 25891
rect 12575 25888 12587 25891
rect 12618 25888 12624 25900
rect 12575 25860 12624 25888
rect 12575 25857 12587 25860
rect 12529 25851 12587 25857
rect 12618 25848 12624 25860
rect 12676 25848 12682 25900
rect 12796 25891 12854 25897
rect 12796 25857 12808 25891
rect 12842 25888 12854 25891
rect 13078 25888 13084 25900
rect 12842 25860 13084 25888
rect 12842 25857 12854 25860
rect 12796 25851 12854 25857
rect 13078 25848 13084 25860
rect 13136 25848 13142 25900
rect 3697 25823 3755 25829
rect 3697 25789 3709 25823
rect 3743 25820 3755 25823
rect 4798 25820 4804 25832
rect 3743 25792 4804 25820
rect 3743 25789 3755 25792
rect 3697 25783 3755 25789
rect 4798 25780 4804 25792
rect 4856 25780 4862 25832
rect 13740 25820 13768 25928
rect 13814 25848 13820 25900
rect 13872 25888 13878 25900
rect 14625 25891 14683 25897
rect 14625 25888 14637 25891
rect 13872 25860 14637 25888
rect 13872 25848 13878 25860
rect 14625 25857 14637 25860
rect 14671 25857 14683 25891
rect 14625 25851 14683 25857
rect 17497 25891 17555 25897
rect 17497 25857 17509 25891
rect 17543 25857 17555 25891
rect 17770 25888 17776 25900
rect 17731 25860 17776 25888
rect 17497 25851 17555 25857
rect 14369 25823 14427 25829
rect 14369 25820 14381 25823
rect 13740 25792 14381 25820
rect 14369 25789 14381 25792
rect 14415 25789 14427 25823
rect 17512 25820 17540 25851
rect 17770 25848 17776 25860
rect 17828 25848 17834 25900
rect 19242 25820 19248 25832
rect 17512 25792 19248 25820
rect 14369 25783 14427 25789
rect 19242 25780 19248 25792
rect 19300 25780 19306 25832
rect 1581 25755 1639 25761
rect 1581 25721 1593 25755
rect 1627 25752 1639 25755
rect 7282 25752 7288 25764
rect 1627 25724 7288 25752
rect 1627 25721 1639 25724
rect 1581 25715 1639 25721
rect 7282 25712 7288 25724
rect 7340 25712 7346 25764
rect 2133 25687 2191 25693
rect 2133 25653 2145 25687
rect 2179 25684 2191 25687
rect 2866 25684 2872 25696
rect 2179 25656 2872 25684
rect 2179 25653 2191 25656
rect 2133 25647 2191 25653
rect 2866 25644 2872 25656
rect 2924 25644 2930 25696
rect 10962 25684 10968 25696
rect 10923 25656 10968 25684
rect 10962 25644 10968 25656
rect 11020 25644 11026 25696
rect 15746 25684 15752 25696
rect 15707 25656 15752 25684
rect 15746 25644 15752 25656
rect 15804 25644 15810 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 1762 25440 1768 25492
rect 1820 25480 1826 25492
rect 1820 25452 9444 25480
rect 1820 25440 1826 25452
rect 7190 25372 7196 25424
rect 7248 25412 7254 25424
rect 7285 25415 7343 25421
rect 7285 25412 7297 25415
rect 7248 25384 7297 25412
rect 7248 25372 7254 25384
rect 7285 25381 7297 25384
rect 7331 25381 7343 25415
rect 9416 25412 9444 25452
rect 9490 25440 9496 25492
rect 9548 25480 9554 25492
rect 9585 25483 9643 25489
rect 9585 25480 9597 25483
rect 9548 25452 9597 25480
rect 9548 25440 9554 25452
rect 9585 25449 9597 25452
rect 9631 25449 9643 25483
rect 10870 25480 10876 25492
rect 10831 25452 10876 25480
rect 9585 25443 9643 25449
rect 10870 25440 10876 25452
rect 10928 25440 10934 25492
rect 13078 25480 13084 25492
rect 13039 25452 13084 25480
rect 13078 25440 13084 25452
rect 13136 25440 13142 25492
rect 10962 25412 10968 25424
rect 9416 25384 10968 25412
rect 7285 25375 7343 25381
rect 1854 25344 1860 25356
rect 1815 25316 1860 25344
rect 1854 25304 1860 25316
rect 1912 25304 1918 25356
rect 5902 25344 5908 25356
rect 5863 25316 5908 25344
rect 5902 25304 5908 25316
rect 5960 25304 5966 25356
rect 10152 25316 10548 25344
rect 1872 25276 1900 25304
rect 3878 25276 3884 25288
rect 1872 25248 3884 25276
rect 3878 25236 3884 25248
rect 3936 25236 3942 25288
rect 8570 25236 8576 25288
rect 8628 25276 8634 25288
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8628 25248 8953 25276
rect 8628 25236 8634 25248
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 9034 25279 9092 25285
rect 9034 25245 9046 25279
rect 9080 25245 9092 25279
rect 9306 25276 9312 25288
rect 9267 25248 9312 25276
rect 9034 25239 9092 25245
rect 2124 25211 2182 25217
rect 2124 25177 2136 25211
rect 2170 25208 2182 25211
rect 2314 25208 2320 25220
rect 2170 25180 2320 25208
rect 2170 25177 2182 25180
rect 2124 25171 2182 25177
rect 2314 25168 2320 25180
rect 2372 25168 2378 25220
rect 6172 25211 6230 25217
rect 6172 25177 6184 25211
rect 6218 25208 6230 25211
rect 7742 25208 7748 25220
rect 6218 25180 7748 25208
rect 6218 25177 6230 25180
rect 6172 25171 6230 25177
rect 7742 25168 7748 25180
rect 7800 25168 7806 25220
rect 7837 25211 7895 25217
rect 7837 25177 7849 25211
rect 7883 25177 7895 25211
rect 7837 25171 7895 25177
rect 3234 25140 3240 25152
rect 3195 25112 3240 25140
rect 3234 25100 3240 25112
rect 3292 25100 3298 25152
rect 5534 25100 5540 25152
rect 5592 25140 5598 25152
rect 7852 25140 7880 25171
rect 8662 25168 8668 25220
rect 8720 25208 8726 25220
rect 9048 25208 9076 25239
rect 9306 25236 9312 25248
rect 9364 25236 9370 25288
rect 9447 25279 9505 25285
rect 9447 25245 9459 25279
rect 9493 25276 9505 25279
rect 9674 25276 9680 25288
rect 9493 25248 9680 25276
rect 9493 25245 9505 25248
rect 9447 25239 9505 25245
rect 9674 25236 9680 25248
rect 9732 25236 9738 25288
rect 8720 25180 9076 25208
rect 9217 25211 9275 25217
rect 8720 25168 8726 25180
rect 9217 25177 9229 25211
rect 9263 25177 9275 25211
rect 9217 25171 9275 25177
rect 8110 25140 8116 25152
rect 5592 25112 7880 25140
rect 8071 25112 8116 25140
rect 5592 25100 5598 25112
rect 8110 25100 8116 25112
rect 8168 25100 8174 25152
rect 9030 25100 9036 25152
rect 9088 25140 9094 25152
rect 9232 25140 9260 25171
rect 10152 25140 10180 25316
rect 10410 25285 10416 25288
rect 10229 25279 10287 25285
rect 10229 25245 10241 25279
rect 10275 25245 10287 25279
rect 10229 25239 10287 25245
rect 10377 25279 10416 25285
rect 10377 25245 10389 25279
rect 10377 25239 10416 25245
rect 10244 25208 10272 25239
rect 10410 25236 10416 25239
rect 10468 25236 10474 25288
rect 10520 25285 10548 25316
rect 10612 25285 10640 25384
rect 10962 25372 10968 25384
rect 11020 25372 11026 25424
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25245 10563 25279
rect 10505 25239 10563 25245
rect 10597 25279 10655 25285
rect 10597 25245 10609 25279
rect 10643 25245 10655 25279
rect 10597 25239 10655 25245
rect 10686 25236 10692 25288
rect 10744 25285 10750 25288
rect 10744 25276 10752 25285
rect 10744 25248 10789 25276
rect 10744 25239 10752 25248
rect 10744 25236 10750 25239
rect 12066 25236 12072 25288
rect 12124 25276 12130 25288
rect 12437 25279 12495 25285
rect 12437 25276 12449 25279
rect 12124 25248 12449 25276
rect 12124 25236 12130 25248
rect 12437 25245 12449 25248
rect 12483 25245 12495 25279
rect 12437 25239 12495 25245
rect 12526 25236 12532 25288
rect 12584 25276 12590 25288
rect 12802 25276 12808 25288
rect 12584 25248 12678 25276
rect 12763 25248 12808 25276
rect 12584 25236 12590 25248
rect 12084 25208 12112 25236
rect 10244 25180 12112 25208
rect 12161 25211 12219 25217
rect 12161 25177 12173 25211
rect 12207 25208 12219 25211
rect 12636 25208 12664 25248
rect 12802 25236 12808 25248
rect 12860 25236 12866 25288
rect 12894 25236 12900 25288
rect 12952 25285 12958 25288
rect 12952 25276 12960 25285
rect 13170 25276 13176 25288
rect 12952 25248 13176 25276
rect 12952 25239 12960 25248
rect 12952 25236 12958 25239
rect 13170 25236 13176 25248
rect 13228 25236 13234 25288
rect 17126 25276 17132 25288
rect 17087 25248 17132 25276
rect 17126 25236 17132 25248
rect 17184 25236 17190 25288
rect 17402 25276 17408 25288
rect 17363 25248 17408 25276
rect 17402 25236 17408 25248
rect 17460 25276 17466 25288
rect 17770 25276 17776 25288
rect 17460 25248 17776 25276
rect 17460 25236 17466 25248
rect 17770 25236 17776 25248
rect 17828 25236 17834 25288
rect 12207 25180 12664 25208
rect 12713 25211 12771 25217
rect 12207 25177 12219 25180
rect 12161 25171 12219 25177
rect 12713 25177 12725 25211
rect 12759 25177 12771 25211
rect 17310 25208 17316 25220
rect 17271 25180 17316 25208
rect 12713 25171 12771 25177
rect 12728 25140 12756 25171
rect 17310 25168 17316 25180
rect 17368 25168 17374 25220
rect 12894 25140 12900 25152
rect 9088 25112 12900 25140
rect 9088 25100 9094 25112
rect 12894 25100 12900 25112
rect 12952 25100 12958 25152
rect 16942 25140 16948 25152
rect 16903 25112 16948 25140
rect 16942 25100 16948 25112
rect 17000 25100 17006 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 2314 24936 2320 24948
rect 2275 24908 2320 24936
rect 2314 24896 2320 24908
rect 2372 24896 2378 24948
rect 7282 24896 7288 24948
rect 7340 24936 7346 24948
rect 21634 24936 21640 24948
rect 7340 24908 21640 24936
rect 7340 24896 7346 24908
rect 21634 24896 21640 24908
rect 21692 24896 21698 24948
rect 1673 24871 1731 24877
rect 1673 24837 1685 24871
rect 1719 24868 1731 24871
rect 5626 24868 5632 24880
rect 1719 24840 5632 24868
rect 1719 24837 1731 24840
rect 1673 24831 1731 24837
rect 5626 24828 5632 24840
rect 5684 24828 5690 24880
rect 9030 24868 9036 24880
rect 8991 24840 9036 24868
rect 9030 24828 9036 24840
rect 9088 24828 9094 24880
rect 13170 24868 13176 24880
rect 12406 24840 13176 24868
rect 1394 24800 1400 24812
rect 1355 24772 1400 24800
rect 1394 24760 1400 24772
rect 1452 24760 1458 24812
rect 2222 24760 2228 24812
rect 2280 24800 2286 24812
rect 2501 24803 2559 24809
rect 2501 24800 2513 24803
rect 2280 24772 2513 24800
rect 2280 24760 2286 24772
rect 2501 24769 2513 24772
rect 2547 24769 2559 24803
rect 3142 24800 3148 24812
rect 3103 24772 3148 24800
rect 2501 24763 2559 24769
rect 3142 24760 3148 24772
rect 3200 24760 3206 24812
rect 3786 24800 3792 24812
rect 3747 24772 3792 24800
rect 3786 24760 3792 24772
rect 3844 24760 3850 24812
rect 4062 24800 4068 24812
rect 4023 24772 4068 24800
rect 4062 24760 4068 24772
rect 4120 24760 4126 24812
rect 8570 24760 8576 24812
rect 8628 24800 8634 24812
rect 8757 24803 8815 24809
rect 8757 24800 8769 24803
rect 8628 24772 8769 24800
rect 8628 24760 8634 24772
rect 8757 24769 8769 24772
rect 8803 24769 8815 24803
rect 8757 24763 8815 24769
rect 8846 24760 8852 24812
rect 8904 24800 8910 24812
rect 9125 24803 9183 24809
rect 8904 24772 8949 24800
rect 8904 24760 8910 24772
rect 9125 24769 9137 24803
rect 9171 24769 9183 24803
rect 9125 24763 9183 24769
rect 9263 24803 9321 24809
rect 9263 24769 9275 24803
rect 9309 24800 9321 24803
rect 9674 24800 9680 24812
rect 9309 24772 9680 24800
rect 9309 24769 9321 24772
rect 9263 24763 9321 24769
rect 3418 24692 3424 24744
rect 3476 24732 3482 24744
rect 3881 24735 3939 24741
rect 3881 24732 3893 24735
rect 3476 24704 3893 24732
rect 3476 24692 3482 24704
rect 3881 24701 3893 24704
rect 3927 24701 3939 24735
rect 3881 24695 3939 24701
rect 7190 24692 7196 24744
rect 7248 24732 7254 24744
rect 9140 24732 9168 24763
rect 9674 24760 9680 24772
rect 9732 24800 9738 24812
rect 10686 24800 10692 24812
rect 9732 24772 10692 24800
rect 9732 24760 9738 24772
rect 10686 24760 10692 24772
rect 10744 24760 10750 24812
rect 10778 24760 10784 24812
rect 10836 24800 10842 24812
rect 11793 24803 11851 24809
rect 11793 24800 11805 24803
rect 10836 24772 11805 24800
rect 10836 24760 10842 24772
rect 11793 24769 11805 24772
rect 11839 24769 11851 24803
rect 11793 24763 11851 24769
rect 11977 24803 12035 24809
rect 11977 24769 11989 24803
rect 12023 24800 12035 24803
rect 12406 24800 12434 24840
rect 13170 24828 13176 24840
rect 13228 24828 13234 24880
rect 16942 24877 16948 24880
rect 16936 24868 16948 24877
rect 16903 24840 16948 24868
rect 16936 24831 16948 24840
rect 16942 24828 16948 24831
rect 17000 24828 17006 24880
rect 12023 24772 12434 24800
rect 12621 24803 12679 24809
rect 12023 24769 12035 24772
rect 11977 24763 12035 24769
rect 12621 24769 12633 24803
rect 12667 24769 12679 24803
rect 12621 24763 12679 24769
rect 7248 24704 9168 24732
rect 12345 24735 12403 24741
rect 7248 24692 7254 24704
rect 12345 24701 12357 24735
rect 12391 24732 12403 24735
rect 12526 24732 12532 24744
rect 12391 24704 12532 24732
rect 12391 24701 12403 24704
rect 12345 24695 12403 24701
rect 12526 24692 12532 24704
rect 12584 24692 12590 24744
rect 2406 24624 2412 24676
rect 2464 24664 2470 24676
rect 2464 24636 9536 24664
rect 2464 24624 2470 24636
rect 2682 24556 2688 24608
rect 2740 24596 2746 24608
rect 2961 24599 3019 24605
rect 2961 24596 2973 24599
rect 2740 24568 2973 24596
rect 2740 24556 2746 24568
rect 2961 24565 2973 24568
rect 3007 24565 3019 24599
rect 2961 24559 3019 24565
rect 3234 24556 3240 24608
rect 3292 24596 3298 24608
rect 3789 24599 3847 24605
rect 3789 24596 3801 24599
rect 3292 24568 3801 24596
rect 3292 24556 3298 24568
rect 3789 24565 3801 24568
rect 3835 24565 3847 24599
rect 3789 24559 3847 24565
rect 4249 24599 4307 24605
rect 4249 24565 4261 24599
rect 4295 24596 4307 24599
rect 6178 24596 6184 24608
rect 4295 24568 6184 24596
rect 4295 24565 4307 24568
rect 4249 24559 4307 24565
rect 6178 24556 6184 24568
rect 6236 24556 6242 24608
rect 7742 24556 7748 24608
rect 7800 24596 7806 24608
rect 9401 24599 9459 24605
rect 9401 24596 9413 24599
rect 7800 24568 9413 24596
rect 7800 24556 7806 24568
rect 9401 24565 9413 24568
rect 9447 24565 9459 24599
rect 9508 24596 9536 24636
rect 12066 24624 12072 24676
rect 12124 24664 12130 24676
rect 12636 24664 12664 24763
rect 12710 24760 12716 24812
rect 12768 24800 12774 24812
rect 12894 24800 12900 24812
rect 12768 24772 12813 24800
rect 12855 24772 12900 24800
rect 12768 24760 12774 24772
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 13086 24803 13144 24809
rect 13086 24769 13098 24803
rect 13132 24800 13144 24803
rect 13188 24800 13216 24828
rect 13132 24772 13216 24800
rect 13132 24769 13144 24772
rect 13086 24763 13144 24769
rect 12124 24636 12664 24664
rect 13004 24732 13032 24763
rect 15746 24732 15752 24744
rect 13004 24704 15752 24732
rect 12124 24624 12130 24636
rect 13004 24596 13032 24704
rect 15746 24692 15752 24704
rect 15804 24692 15810 24744
rect 16669 24735 16727 24741
rect 16669 24701 16681 24735
rect 16715 24701 16727 24735
rect 16669 24695 16727 24701
rect 13265 24667 13323 24673
rect 13265 24633 13277 24667
rect 13311 24664 13323 24667
rect 13814 24664 13820 24676
rect 13311 24636 13820 24664
rect 13311 24633 13323 24636
rect 13265 24627 13323 24633
rect 13814 24624 13820 24636
rect 13872 24624 13878 24676
rect 15194 24624 15200 24676
rect 15252 24664 15258 24676
rect 16684 24664 16712 24695
rect 15252 24636 16712 24664
rect 15252 24624 15258 24636
rect 9508 24568 13032 24596
rect 9401 24559 9459 24565
rect 17310 24556 17316 24608
rect 17368 24596 17374 24608
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 17368 24568 18061 24596
rect 17368 24556 17374 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 2222 24392 2228 24404
rect 2183 24364 2228 24392
rect 2222 24352 2228 24364
rect 2280 24352 2286 24404
rect 4062 24352 4068 24404
rect 4120 24392 4126 24404
rect 5169 24395 5227 24401
rect 5169 24392 5181 24395
rect 4120 24364 5181 24392
rect 4120 24352 4126 24364
rect 5169 24361 5181 24364
rect 5215 24361 5227 24395
rect 24578 24392 24584 24404
rect 5169 24355 5227 24361
rect 12406 24364 24584 24392
rect 2682 24256 2688 24268
rect 2643 24228 2688 24256
rect 2682 24216 2688 24228
rect 2740 24216 2746 24268
rect 2869 24259 2927 24265
rect 2869 24225 2881 24259
rect 2915 24256 2927 24259
rect 3050 24256 3056 24268
rect 2915 24228 3056 24256
rect 2915 24225 2927 24228
rect 2869 24219 2927 24225
rect 3050 24216 3056 24228
rect 3108 24216 3114 24268
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24148 1458 24200
rect 2593 24191 2651 24197
rect 2593 24157 2605 24191
rect 2639 24188 2651 24191
rect 3234 24188 3240 24200
rect 2639 24160 3240 24188
rect 2639 24157 2651 24160
rect 2593 24151 2651 24157
rect 3234 24148 3240 24160
rect 3292 24148 3298 24200
rect 3796 24191 3854 24197
rect 3796 24157 3808 24191
rect 3842 24188 3854 24191
rect 3842 24160 3924 24188
rect 3842 24157 3854 24160
rect 3796 24151 3854 24157
rect 3896 24064 3924 24160
rect 5626 24148 5632 24200
rect 5684 24188 5690 24200
rect 12406 24188 12434 24364
rect 24578 24352 24584 24364
rect 24636 24352 24642 24404
rect 12805 24259 12863 24265
rect 12805 24225 12817 24259
rect 12851 24256 12863 24259
rect 12894 24256 12900 24268
rect 12851 24228 12900 24256
rect 12851 24225 12863 24228
rect 12805 24219 12863 24225
rect 12894 24216 12900 24228
rect 12952 24216 12958 24268
rect 12526 24188 12532 24200
rect 5684 24160 12434 24188
rect 12487 24160 12532 24188
rect 5684 24148 5690 24160
rect 12526 24148 12532 24160
rect 12584 24148 12590 24200
rect 15194 24148 15200 24200
rect 15252 24188 15258 24200
rect 15473 24191 15531 24197
rect 15473 24188 15485 24191
rect 15252 24160 15485 24188
rect 15252 24148 15258 24160
rect 15473 24157 15485 24160
rect 15519 24157 15531 24191
rect 17402 24188 17408 24200
rect 15473 24151 15531 24157
rect 15672 24160 17408 24188
rect 4056 24123 4114 24129
rect 4056 24089 4068 24123
rect 4102 24120 4114 24123
rect 4154 24120 4160 24132
rect 4102 24092 4160 24120
rect 4102 24089 4114 24092
rect 4056 24083 4114 24089
rect 4154 24080 4160 24092
rect 4212 24080 4218 24132
rect 13814 24080 13820 24132
rect 13872 24120 13878 24132
rect 14553 24123 14611 24129
rect 14553 24120 14565 24123
rect 13872 24092 14565 24120
rect 13872 24080 13878 24092
rect 14553 24089 14565 24092
rect 14599 24089 14611 24123
rect 14553 24083 14611 24089
rect 14737 24123 14795 24129
rect 14737 24089 14749 24123
rect 14783 24120 14795 24123
rect 15672 24120 15700 24160
rect 17402 24148 17408 24160
rect 17460 24148 17466 24200
rect 15746 24129 15752 24132
rect 14783 24092 15700 24120
rect 14783 24089 14795 24092
rect 14737 24083 14795 24089
rect 15740 24083 15752 24129
rect 15804 24120 15810 24132
rect 15804 24092 15840 24120
rect 15746 24080 15752 24083
rect 15804 24080 15810 24092
rect 1578 24052 1584 24064
rect 1539 24024 1584 24052
rect 1578 24012 1584 24024
rect 1636 24012 1642 24064
rect 3878 24012 3884 24064
rect 3936 24012 3942 24064
rect 5442 24012 5448 24064
rect 5500 24052 5506 24064
rect 11882 24052 11888 24064
rect 5500 24024 11888 24052
rect 5500 24012 5506 24024
rect 11882 24012 11888 24024
rect 11940 24012 11946 24064
rect 16022 24012 16028 24064
rect 16080 24052 16086 24064
rect 16853 24055 16911 24061
rect 16853 24052 16865 24055
rect 16080 24024 16865 24052
rect 16080 24012 16086 24024
rect 16853 24021 16865 24024
rect 16899 24021 16911 24055
rect 16853 24015 16911 24021
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 2409 23851 2467 23857
rect 2409 23817 2421 23851
rect 2455 23817 2467 23851
rect 2409 23811 2467 23817
rect 3421 23851 3479 23857
rect 3421 23817 3433 23851
rect 3467 23848 3479 23851
rect 4062 23848 4068 23860
rect 3467 23820 4068 23848
rect 3467 23817 3479 23820
rect 3421 23811 3479 23817
rect 2424 23780 2452 23811
rect 4062 23808 4068 23820
rect 4120 23808 4126 23860
rect 8849 23851 8907 23857
rect 8849 23817 8861 23851
rect 8895 23848 8907 23851
rect 8938 23848 8944 23860
rect 8895 23820 8944 23848
rect 8895 23817 8907 23820
rect 8849 23811 8907 23817
rect 8938 23808 8944 23820
rect 8996 23808 9002 23860
rect 9953 23851 10011 23857
rect 9953 23817 9965 23851
rect 9999 23817 10011 23851
rect 12710 23848 12716 23860
rect 9953 23811 10011 23817
rect 11532 23820 12716 23848
rect 4154 23780 4160 23792
rect 2424 23752 4160 23780
rect 4154 23740 4160 23752
rect 4212 23740 4218 23792
rect 7736 23783 7794 23789
rect 7736 23749 7748 23783
rect 7782 23780 7794 23783
rect 9968 23780 9996 23811
rect 10778 23780 10784 23792
rect 7782 23752 9996 23780
rect 10739 23752 10784 23780
rect 7782 23749 7794 23752
rect 7736 23743 7794 23749
rect 10778 23740 10784 23752
rect 10836 23740 10842 23792
rect 1394 23712 1400 23724
rect 1355 23684 1400 23712
rect 1394 23672 1400 23684
rect 1452 23672 1458 23724
rect 2593 23715 2651 23721
rect 2593 23681 2605 23715
rect 2639 23712 2651 23715
rect 4341 23715 4399 23721
rect 2639 23684 2774 23712
rect 2639 23681 2651 23684
rect 2593 23675 2651 23681
rect 2746 23576 2774 23684
rect 4341 23681 4353 23715
rect 4387 23712 4399 23715
rect 5534 23712 5540 23724
rect 4387 23684 5540 23712
rect 4387 23681 4399 23684
rect 4341 23675 4399 23681
rect 5534 23672 5540 23684
rect 5592 23712 5598 23724
rect 6454 23712 6460 23724
rect 5592 23684 6460 23712
rect 5592 23672 5598 23684
rect 6454 23672 6460 23684
rect 6512 23672 6518 23724
rect 9306 23712 9312 23724
rect 9267 23684 9312 23712
rect 9306 23672 9312 23684
rect 9364 23672 9370 23724
rect 9398 23672 9404 23724
rect 9456 23712 9462 23724
rect 9582 23712 9588 23724
rect 9456 23684 9501 23712
rect 9543 23684 9588 23712
rect 9456 23672 9462 23684
rect 9582 23672 9588 23684
rect 9640 23672 9646 23724
rect 9677 23715 9735 23721
rect 9677 23681 9689 23715
rect 9723 23681 9735 23715
rect 9677 23675 9735 23681
rect 9815 23715 9873 23721
rect 9815 23681 9827 23715
rect 9861 23712 9873 23715
rect 10686 23712 10692 23724
rect 9861 23684 10692 23712
rect 9861 23681 9873 23684
rect 9815 23675 9873 23681
rect 3510 23644 3516 23656
rect 3471 23616 3516 23644
rect 3510 23604 3516 23616
rect 3568 23604 3574 23656
rect 3605 23647 3663 23653
rect 3605 23613 3617 23647
rect 3651 23613 3663 23647
rect 3605 23607 3663 23613
rect 3053 23579 3111 23585
rect 3053 23576 3065 23579
rect 2746 23548 3065 23576
rect 3053 23545 3065 23548
rect 3099 23545 3111 23579
rect 3053 23539 3111 23545
rect 3142 23536 3148 23588
rect 3200 23576 3206 23588
rect 3620 23576 3648 23607
rect 7098 23604 7104 23656
rect 7156 23644 7162 23656
rect 7469 23647 7527 23653
rect 7469 23644 7481 23647
rect 7156 23616 7481 23644
rect 7156 23604 7162 23616
rect 7469 23613 7481 23616
rect 7515 23613 7527 23647
rect 7469 23607 7527 23613
rect 8938 23604 8944 23656
rect 8996 23644 9002 23656
rect 9692 23644 9720 23675
rect 10686 23672 10692 23684
rect 10744 23712 10750 23724
rect 11532 23721 11560 23820
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 15657 23851 15715 23857
rect 15657 23817 15669 23851
rect 15703 23848 15715 23851
rect 15746 23848 15752 23860
rect 15703 23820 15752 23848
rect 15703 23817 15715 23820
rect 15657 23811 15715 23817
rect 15746 23808 15752 23820
rect 15804 23808 15810 23860
rect 16114 23808 16120 23860
rect 16172 23808 16178 23860
rect 15102 23740 15108 23792
rect 15160 23780 15166 23792
rect 16022 23780 16028 23792
rect 15160 23752 16028 23780
rect 15160 23740 15166 23752
rect 16022 23740 16028 23752
rect 16080 23740 16086 23792
rect 11790 23721 11796 23724
rect 11517 23715 11575 23721
rect 10744 23684 11008 23712
rect 10744 23672 10750 23684
rect 8996 23616 9720 23644
rect 8996 23604 9002 23616
rect 10980 23588 11008 23684
rect 11517 23681 11529 23715
rect 11563 23681 11575 23715
rect 11517 23675 11575 23681
rect 11784 23675 11796 23721
rect 11848 23712 11854 23724
rect 16132 23721 16160 23808
rect 15841 23715 15899 23721
rect 11848 23684 11884 23712
rect 11790 23672 11796 23675
rect 11848 23672 11854 23684
rect 15841 23681 15853 23715
rect 15887 23681 15899 23715
rect 15841 23675 15899 23681
rect 16117 23715 16175 23721
rect 16117 23681 16129 23715
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 15856 23644 15884 23675
rect 17402 23644 17408 23656
rect 15856 23616 17408 23644
rect 17402 23604 17408 23616
rect 17460 23604 17466 23656
rect 4525 23579 4583 23585
rect 4525 23576 4537 23579
rect 3200 23548 4537 23576
rect 3200 23536 3206 23548
rect 4525 23545 4537 23548
rect 4571 23545 4583 23579
rect 10962 23576 10968 23588
rect 10923 23548 10968 23576
rect 4525 23539 4583 23545
rect 10962 23536 10968 23548
rect 11020 23536 11026 23588
rect 1578 23508 1584 23520
rect 1539 23480 1584 23508
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 3602 23468 3608 23520
rect 3660 23508 3666 23520
rect 11698 23508 11704 23520
rect 3660 23480 11704 23508
rect 3660 23468 3666 23480
rect 11698 23468 11704 23480
rect 11756 23508 11762 23520
rect 12897 23511 12955 23517
rect 12897 23508 12909 23511
rect 11756 23480 12909 23508
rect 11756 23468 11762 23480
rect 12897 23477 12909 23480
rect 12943 23477 12955 23511
rect 12897 23471 12955 23477
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 2041 23307 2099 23313
rect 2041 23273 2053 23307
rect 2087 23304 2099 23307
rect 3510 23304 3516 23316
rect 2087 23276 3516 23304
rect 2087 23273 2099 23276
rect 2041 23267 2099 23273
rect 3510 23264 3516 23276
rect 3568 23264 3574 23316
rect 8389 23307 8447 23313
rect 8389 23304 8401 23307
rect 6748 23276 8401 23304
rect 2498 23196 2504 23248
rect 2556 23236 2562 23248
rect 6748 23236 6776 23276
rect 8389 23273 8401 23276
rect 8435 23304 8447 23307
rect 9030 23304 9036 23316
rect 8435 23276 9036 23304
rect 8435 23273 8447 23276
rect 8389 23267 8447 23273
rect 9030 23264 9036 23276
rect 9088 23264 9094 23316
rect 11790 23264 11796 23316
rect 11848 23304 11854 23316
rect 11885 23307 11943 23313
rect 11885 23304 11897 23307
rect 11848 23276 11897 23304
rect 11848 23264 11854 23276
rect 11885 23273 11897 23276
rect 11931 23273 11943 23307
rect 15194 23304 15200 23316
rect 11885 23267 11943 23273
rect 14108 23276 15200 23304
rect 2556 23208 6776 23236
rect 2556 23196 2562 23208
rect 8570 23128 8576 23180
rect 8628 23168 8634 23180
rect 9306 23168 9312 23180
rect 8628 23140 9312 23168
rect 8628 23128 8634 23140
rect 9306 23128 9312 23140
rect 9364 23168 9370 23180
rect 9364 23140 10916 23168
rect 9364 23128 9370 23140
rect 1394 23060 1400 23112
rect 1452 23100 1458 23112
rect 1581 23103 1639 23109
rect 1581 23100 1593 23103
rect 1452 23072 1593 23100
rect 1452 23060 1458 23072
rect 1581 23069 1593 23072
rect 1627 23069 1639 23103
rect 2222 23100 2228 23112
rect 2183 23072 2228 23100
rect 1581 23063 1639 23069
rect 2222 23060 2228 23072
rect 2280 23060 2286 23112
rect 7009 23103 7067 23109
rect 7009 23069 7021 23103
rect 7055 23100 7067 23103
rect 7098 23100 7104 23112
rect 7055 23072 7104 23100
rect 7055 23069 7067 23072
rect 7009 23063 7067 23069
rect 7098 23060 7104 23072
rect 7156 23060 7162 23112
rect 10505 23103 10563 23109
rect 10505 23069 10517 23103
rect 10551 23100 10563 23103
rect 10778 23100 10784 23112
rect 10551 23072 10784 23100
rect 10551 23069 10563 23072
rect 10505 23063 10563 23069
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 10888 23100 10916 23140
rect 10962 23128 10968 23180
rect 11020 23168 11026 23180
rect 11020 23140 11744 23168
rect 11020 23128 11026 23140
rect 11238 23100 11244 23112
rect 10888 23072 11244 23100
rect 11238 23060 11244 23072
rect 11296 23060 11302 23112
rect 11330 23060 11336 23112
rect 11388 23100 11394 23112
rect 11606 23100 11612 23112
rect 11388 23072 11433 23100
rect 11567 23072 11612 23100
rect 11388 23060 11394 23072
rect 11606 23060 11612 23072
rect 11664 23060 11670 23112
rect 11716 23109 11744 23140
rect 12710 23128 12716 23180
rect 12768 23168 12774 23180
rect 14108 23177 14136 23276
rect 15194 23264 15200 23276
rect 15252 23264 15258 23316
rect 14093 23171 14151 23177
rect 14093 23168 14105 23171
rect 12768 23140 14105 23168
rect 12768 23128 12774 23140
rect 14093 23137 14105 23140
rect 14139 23137 14151 23171
rect 14093 23131 14151 23137
rect 15746 23128 15752 23180
rect 15804 23168 15810 23180
rect 17405 23171 17463 23177
rect 17405 23168 17417 23171
rect 15804 23140 17417 23168
rect 15804 23128 15810 23140
rect 17405 23137 17417 23140
rect 17451 23137 17463 23171
rect 17405 23131 17463 23137
rect 17497 23171 17555 23177
rect 17497 23137 17509 23171
rect 17543 23168 17555 23171
rect 17543 23140 20116 23168
rect 17543 23137 17555 23140
rect 17497 23131 17555 23137
rect 11706 23103 11764 23109
rect 11706 23069 11718 23103
rect 11752 23069 11764 23103
rect 11706 23063 11764 23069
rect 11882 23060 11888 23112
rect 11940 23100 11946 23112
rect 17310 23100 17316 23112
rect 11940 23072 14044 23100
rect 17271 23072 17316 23100
rect 11940 23060 11946 23072
rect 7276 23035 7334 23041
rect 7276 23001 7288 23035
rect 7322 23032 7334 23035
rect 9306 23032 9312 23044
rect 7322 23004 9312 23032
rect 7322 23001 7334 23004
rect 7276 22995 7334 23001
rect 9306 22992 9312 23004
rect 9364 22992 9370 23044
rect 9582 22992 9588 23044
rect 9640 23032 9646 23044
rect 11517 23035 11575 23041
rect 11517 23032 11529 23035
rect 9640 23004 11529 23032
rect 9640 22992 9646 23004
rect 11517 23001 11529 23004
rect 11563 23032 11575 23035
rect 12526 23032 12532 23044
rect 11563 23004 12532 23032
rect 11563 23001 11575 23004
rect 11517 22995 11575 23001
rect 12526 22992 12532 23004
rect 12584 23032 12590 23044
rect 13262 23032 13268 23044
rect 12584 23004 13268 23032
rect 12584 22992 12590 23004
rect 13262 22992 13268 23004
rect 13320 22992 13326 23044
rect 1397 22967 1455 22973
rect 1397 22933 1409 22967
rect 1443 22964 1455 22967
rect 2958 22964 2964 22976
rect 1443 22936 2964 22964
rect 1443 22933 1455 22936
rect 1397 22927 1455 22933
rect 2958 22924 2964 22936
rect 3016 22924 3022 22976
rect 5626 22924 5632 22976
rect 5684 22964 5690 22976
rect 9214 22964 9220 22976
rect 5684 22936 9220 22964
rect 5684 22924 5690 22936
rect 9214 22924 9220 22936
rect 9272 22964 9278 22976
rect 10689 22967 10747 22973
rect 10689 22964 10701 22967
rect 9272 22936 10701 22964
rect 9272 22924 9278 22936
rect 10689 22933 10701 22936
rect 10735 22964 10747 22967
rect 11422 22964 11428 22976
rect 10735 22936 11428 22964
rect 10735 22933 10747 22936
rect 10689 22927 10747 22933
rect 11422 22924 11428 22936
rect 11480 22924 11486 22976
rect 11790 22924 11796 22976
rect 11848 22964 11854 22976
rect 13814 22964 13820 22976
rect 11848 22936 13820 22964
rect 11848 22924 11854 22936
rect 13814 22924 13820 22936
rect 13872 22924 13878 22976
rect 14016 22964 14044 23072
rect 17310 23060 17316 23072
rect 17368 23060 17374 23112
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23069 17647 23103
rect 19978 23100 19984 23112
rect 19939 23072 19984 23100
rect 17589 23063 17647 23069
rect 14182 22992 14188 23044
rect 14240 23032 14246 23044
rect 14338 23035 14396 23041
rect 14338 23032 14350 23035
rect 14240 23004 14350 23032
rect 14240 22992 14246 23004
rect 14338 23001 14350 23004
rect 14384 23001 14396 23035
rect 14338 22995 14396 23001
rect 17494 22992 17500 23044
rect 17552 23032 17558 23044
rect 17604 23032 17632 23063
rect 19978 23060 19984 23072
rect 20036 23060 20042 23112
rect 20088 23100 20116 23140
rect 22462 23128 22468 23180
rect 22520 23168 22526 23180
rect 22520 23140 24440 23168
rect 22520 23128 22526 23140
rect 24412 23109 24440 23140
rect 24397 23103 24455 23109
rect 20088 23072 24256 23100
rect 17552 23004 17632 23032
rect 20248 23035 20306 23041
rect 17552 22992 17558 23004
rect 20248 23001 20260 23035
rect 20294 23032 20306 23035
rect 20806 23032 20812 23044
rect 20294 23004 20812 23032
rect 20294 23001 20306 23004
rect 20248 22995 20306 23001
rect 20806 22992 20812 23004
rect 20864 22992 20870 23044
rect 14458 22964 14464 22976
rect 14016 22936 14464 22964
rect 14458 22924 14464 22936
rect 14516 22964 14522 22976
rect 15473 22967 15531 22973
rect 15473 22964 15485 22967
rect 14516 22936 15485 22964
rect 14516 22924 14522 22936
rect 15473 22933 15485 22936
rect 15519 22933 15531 22967
rect 15473 22927 15531 22933
rect 15930 22924 15936 22976
rect 15988 22964 15994 22976
rect 17129 22967 17187 22973
rect 17129 22964 17141 22967
rect 15988 22936 17141 22964
rect 15988 22924 15994 22936
rect 17129 22933 17141 22936
rect 17175 22933 17187 22967
rect 17129 22927 17187 22933
rect 20346 22924 20352 22976
rect 20404 22964 20410 22976
rect 21361 22967 21419 22973
rect 21361 22964 21373 22967
rect 20404 22936 21373 22964
rect 20404 22924 20410 22936
rect 21361 22933 21373 22936
rect 21407 22933 21419 22967
rect 24228 22964 24256 23072
rect 24397 23069 24409 23103
rect 24443 23100 24455 23103
rect 27614 23100 27620 23112
rect 24443 23072 27620 23100
rect 24443 23069 24455 23072
rect 24397 23063 24455 23069
rect 27614 23060 27620 23072
rect 27672 23060 27678 23112
rect 29730 23060 29736 23112
rect 29788 23100 29794 23112
rect 33229 23103 33287 23109
rect 33229 23100 33241 23103
rect 29788 23072 33241 23100
rect 29788 23060 29794 23072
rect 33229 23069 33241 23072
rect 33275 23069 33287 23103
rect 33502 23100 33508 23112
rect 33463 23072 33508 23100
rect 33229 23063 33287 23069
rect 33502 23060 33508 23072
rect 33560 23060 33566 23112
rect 24670 23041 24676 23044
rect 24664 22995 24676 23041
rect 24728 23032 24734 23044
rect 27884 23035 27942 23041
rect 24728 23004 24764 23032
rect 24670 22992 24676 22995
rect 24728 22992 24734 23004
rect 27884 23001 27896 23035
rect 27930 23032 27942 23035
rect 27982 23032 27988 23044
rect 27930 23004 27988 23032
rect 27930 23001 27942 23004
rect 27884 22995 27942 23001
rect 27982 22992 27988 23004
rect 28040 22992 28046 23044
rect 25038 22964 25044 22976
rect 24228 22936 25044 22964
rect 21361 22927 21419 22933
rect 25038 22924 25044 22936
rect 25096 22964 25102 22976
rect 25777 22967 25835 22973
rect 25777 22964 25789 22967
rect 25096 22936 25789 22964
rect 25096 22924 25102 22936
rect 25777 22933 25789 22936
rect 25823 22933 25835 22967
rect 25777 22927 25835 22933
rect 28997 22967 29055 22973
rect 28997 22933 29009 22967
rect 29043 22964 29055 22967
rect 29546 22964 29552 22976
rect 29043 22936 29552 22964
rect 29043 22933 29055 22936
rect 28997 22927 29055 22933
rect 29546 22924 29552 22936
rect 29604 22924 29610 22976
rect 33042 22964 33048 22976
rect 33003 22936 33048 22964
rect 33042 22924 33048 22936
rect 33100 22924 33106 22976
rect 33410 22964 33416 22976
rect 33371 22936 33416 22964
rect 33410 22924 33416 22936
rect 33468 22924 33474 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1578 22720 1584 22772
rect 1636 22760 1642 22772
rect 2961 22763 3019 22769
rect 1636 22732 2774 22760
rect 1636 22720 1642 22732
rect 2746 22692 2774 22732
rect 2961 22729 2973 22763
rect 3007 22760 3019 22763
rect 4890 22760 4896 22772
rect 3007 22732 4896 22760
rect 3007 22729 3019 22732
rect 2961 22723 3019 22729
rect 4890 22720 4896 22732
rect 4948 22760 4954 22772
rect 5169 22763 5227 22769
rect 5169 22760 5181 22763
rect 4948 22732 5181 22760
rect 4948 22720 4954 22732
rect 5169 22729 5181 22732
rect 5215 22729 5227 22763
rect 9306 22760 9312 22772
rect 9267 22732 9312 22760
rect 5169 22723 5227 22729
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 12434 22720 12440 22772
rect 12492 22760 12498 22772
rect 12710 22760 12716 22772
rect 12492 22732 12716 22760
rect 12492 22720 12498 22732
rect 12710 22720 12716 22732
rect 12768 22720 12774 22772
rect 14093 22763 14151 22769
rect 14093 22729 14105 22763
rect 14139 22760 14151 22763
rect 14182 22760 14188 22772
rect 14139 22732 14188 22760
rect 14139 22729 14151 22732
rect 14093 22723 14151 22729
rect 14182 22720 14188 22732
rect 14240 22720 14246 22772
rect 14458 22760 14464 22772
rect 14419 22732 14464 22760
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 17589 22763 17647 22769
rect 17589 22760 17601 22763
rect 17276 22732 17601 22760
rect 17276 22720 17282 22732
rect 17589 22729 17601 22732
rect 17635 22729 17647 22763
rect 20806 22760 20812 22772
rect 20767 22732 20812 22760
rect 17589 22723 17647 22729
rect 20806 22720 20812 22732
rect 20864 22720 20870 22772
rect 24670 22760 24676 22772
rect 24631 22732 24676 22760
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 25038 22760 25044 22772
rect 24999 22732 25044 22760
rect 25038 22720 25044 22732
rect 25096 22720 25102 22772
rect 27982 22760 27988 22772
rect 27943 22732 27988 22760
rect 27982 22720 27988 22732
rect 28040 22720 28046 22772
rect 28166 22720 28172 22772
rect 28224 22760 28230 22772
rect 28353 22763 28411 22769
rect 28353 22760 28365 22763
rect 28224 22732 28365 22760
rect 28224 22720 28230 22732
rect 28353 22729 28365 22732
rect 28399 22760 28411 22763
rect 33410 22760 33416 22772
rect 28399 22732 33416 22760
rect 28399 22729 28411 22732
rect 28353 22723 28411 22729
rect 33410 22720 33416 22732
rect 33468 22720 33474 22772
rect 13449 22695 13507 22701
rect 2746 22664 10272 22692
rect 1397 22627 1455 22633
rect 1397 22593 1409 22627
rect 1443 22624 1455 22627
rect 2774 22624 2780 22636
rect 1443 22596 2780 22624
rect 1443 22593 1455 22596
rect 1397 22587 1455 22593
rect 2774 22584 2780 22596
rect 2832 22584 2838 22636
rect 2866 22584 2872 22636
rect 2924 22624 2930 22636
rect 3053 22627 3111 22633
rect 3053 22624 3065 22627
rect 2924 22596 3065 22624
rect 2924 22584 2930 22596
rect 3053 22593 3065 22596
rect 3099 22593 3111 22627
rect 3786 22624 3792 22636
rect 3747 22596 3792 22624
rect 3053 22587 3111 22593
rect 3786 22584 3792 22596
rect 3844 22584 3850 22636
rect 3878 22584 3884 22636
rect 3936 22624 3942 22636
rect 4045 22627 4103 22633
rect 4045 22624 4057 22627
rect 3936 22596 4057 22624
rect 3936 22584 3942 22596
rect 4045 22593 4057 22596
rect 4091 22593 4103 22627
rect 4045 22587 4103 22593
rect 8570 22584 8576 22636
rect 8628 22624 8634 22636
rect 8846 22633 8852 22636
rect 8665 22627 8723 22633
rect 8665 22624 8677 22627
rect 8628 22596 8677 22624
rect 8628 22584 8634 22596
rect 8665 22593 8677 22596
rect 8711 22593 8723 22627
rect 8665 22587 8723 22593
rect 8813 22627 8852 22633
rect 8813 22593 8825 22627
rect 8813 22587 8852 22593
rect 8846 22584 8852 22587
rect 8904 22584 8910 22636
rect 8941 22627 8999 22633
rect 8941 22593 8953 22627
rect 8987 22593 8999 22627
rect 8941 22587 8999 22593
rect 3142 22516 3148 22568
rect 3200 22556 3206 22568
rect 8956 22556 8984 22587
rect 9030 22584 9036 22636
rect 9088 22624 9094 22636
rect 9214 22633 9220 22636
rect 9171 22627 9220 22633
rect 9088 22596 9133 22624
rect 9088 22584 9094 22596
rect 9171 22593 9183 22627
rect 9217 22593 9220 22627
rect 9171 22587 9220 22593
rect 9214 22584 9220 22587
rect 9272 22584 9278 22636
rect 9582 22556 9588 22568
rect 3200 22528 3245 22556
rect 8956 22528 9588 22556
rect 3200 22516 3206 22528
rect 9582 22516 9588 22528
rect 9640 22516 9646 22568
rect 10244 22556 10272 22664
rect 13449 22661 13461 22695
rect 13495 22692 13507 22695
rect 13814 22692 13820 22704
rect 13495 22664 13820 22692
rect 13495 22661 13507 22664
rect 13449 22655 13507 22661
rect 13814 22652 13820 22664
rect 13872 22652 13878 22704
rect 13924 22664 14596 22692
rect 13630 22624 13636 22636
rect 13543 22596 13636 22624
rect 13630 22584 13636 22596
rect 13688 22624 13694 22636
rect 13924 22624 13952 22664
rect 14568 22633 14596 22664
rect 17604 22664 18092 22692
rect 17604 22636 17632 22664
rect 13688 22596 13952 22624
rect 14277 22627 14335 22633
rect 13688 22584 13694 22596
rect 14277 22593 14289 22627
rect 14323 22593 14335 22627
rect 14277 22587 14335 22593
rect 14553 22627 14611 22633
rect 14553 22593 14565 22627
rect 14599 22624 14611 22627
rect 16114 22624 16120 22636
rect 14599 22596 16120 22624
rect 14599 22593 14611 22596
rect 14553 22587 14611 22593
rect 14292 22556 14320 22587
rect 16114 22584 16120 22596
rect 16172 22584 16178 22636
rect 17586 22584 17592 22636
rect 17644 22584 17650 22636
rect 17678 22584 17684 22636
rect 17736 22624 17742 22636
rect 18064 22633 18092 22664
rect 20346 22652 20352 22704
rect 20404 22692 20410 22704
rect 21177 22695 21235 22701
rect 21177 22692 21189 22695
rect 20404 22664 21189 22692
rect 20404 22652 20410 22664
rect 21177 22661 21189 22664
rect 21223 22661 21235 22695
rect 25682 22692 25688 22704
rect 21177 22655 21235 22661
rect 24780 22664 25688 22692
rect 17865 22627 17923 22633
rect 17865 22624 17877 22627
rect 17736 22596 17877 22624
rect 17736 22584 17742 22596
rect 17865 22593 17877 22596
rect 17911 22593 17923 22627
rect 17865 22587 17923 22593
rect 18049 22627 18107 22633
rect 18049 22593 18061 22627
rect 18095 22593 18107 22627
rect 18049 22587 18107 22593
rect 20993 22627 21051 22633
rect 20993 22593 21005 22627
rect 21039 22593 21051 22627
rect 21266 22624 21272 22636
rect 21227 22596 21272 22624
rect 20993 22587 21051 22593
rect 16022 22556 16028 22568
rect 10244 22528 13860 22556
rect 14292 22528 16028 22556
rect 13832 22488 13860 22528
rect 16022 22516 16028 22528
rect 16080 22516 16086 22568
rect 17770 22556 17776 22568
rect 17731 22528 17776 22556
rect 17770 22516 17776 22528
rect 17828 22516 17834 22568
rect 17954 22516 17960 22568
rect 18012 22556 18018 22568
rect 21008 22556 21036 22587
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 24780 22556 24808 22664
rect 25682 22652 25688 22664
rect 25740 22692 25746 22704
rect 25740 22664 26234 22692
rect 25740 22652 25746 22664
rect 24857 22627 24915 22633
rect 24857 22593 24869 22627
rect 24903 22593 24915 22627
rect 24857 22587 24915 22593
rect 18012 22528 18057 22556
rect 21008 22528 24808 22556
rect 24872 22556 24900 22587
rect 25038 22584 25044 22636
rect 25096 22624 25102 22636
rect 25133 22627 25191 22633
rect 25133 22624 25145 22627
rect 25096 22596 25145 22624
rect 25096 22584 25102 22596
rect 25133 22593 25145 22596
rect 25179 22593 25191 22627
rect 26206 22624 26234 22664
rect 33042 22652 33048 22704
rect 33100 22692 33106 22704
rect 33290 22695 33348 22701
rect 33290 22692 33302 22695
rect 33100 22664 33302 22692
rect 33100 22652 33106 22664
rect 33290 22661 33302 22664
rect 33336 22661 33348 22695
rect 33290 22655 33348 22661
rect 28169 22627 28227 22633
rect 28169 22624 28181 22627
rect 26206 22596 28181 22624
rect 25133 22587 25191 22593
rect 28169 22593 28181 22596
rect 28215 22593 28227 22627
rect 28169 22587 28227 22593
rect 28445 22627 28503 22633
rect 28445 22593 28457 22627
rect 28491 22624 28503 22627
rect 29638 22624 29644 22636
rect 28491 22596 29644 22624
rect 28491 22593 28503 22596
rect 28445 22587 28503 22593
rect 29638 22584 29644 22596
rect 29696 22584 29702 22636
rect 30460 22627 30518 22633
rect 30460 22593 30472 22627
rect 30506 22624 30518 22627
rect 30834 22624 30840 22636
rect 30506 22596 30840 22624
rect 30506 22593 30518 22596
rect 30460 22587 30518 22593
rect 30834 22584 30840 22596
rect 30892 22584 30898 22636
rect 25774 22556 25780 22568
rect 24872 22528 25780 22556
rect 18012 22516 18018 22528
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 30193 22559 30251 22565
rect 30193 22525 30205 22559
rect 30239 22525 30251 22559
rect 30193 22519 30251 22525
rect 33045 22559 33103 22565
rect 33045 22525 33057 22559
rect 33091 22525 33103 22559
rect 33045 22519 33103 22525
rect 28258 22488 28264 22500
rect 13832 22460 28264 22488
rect 28258 22448 28264 22460
rect 28316 22448 28322 22500
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 2593 22423 2651 22429
rect 2593 22389 2605 22423
rect 2639 22420 2651 22423
rect 3970 22420 3976 22432
rect 2639 22392 3976 22420
rect 2639 22389 2651 22392
rect 2593 22383 2651 22389
rect 3970 22380 3976 22392
rect 4028 22380 4034 22432
rect 17218 22380 17224 22432
rect 17276 22420 17282 22432
rect 17494 22420 17500 22432
rect 17276 22392 17500 22420
rect 17276 22380 17282 22392
rect 17494 22380 17500 22392
rect 17552 22420 17558 22432
rect 18230 22420 18236 22432
rect 17552 22392 18236 22420
rect 17552 22380 17558 22392
rect 18230 22380 18236 22392
rect 18288 22380 18294 22432
rect 27614 22380 27620 22432
rect 27672 22420 27678 22432
rect 30208 22420 30236 22519
rect 33060 22488 33088 22519
rect 31128 22460 33088 22488
rect 31128 22420 31156 22460
rect 27672 22392 31156 22420
rect 31573 22423 31631 22429
rect 27672 22380 27678 22392
rect 31573 22389 31585 22423
rect 31619 22420 31631 22423
rect 32030 22420 32036 22432
rect 31619 22392 32036 22420
rect 31619 22389 31631 22392
rect 31573 22383 31631 22389
rect 32030 22380 32036 22392
rect 32088 22380 32094 22432
rect 33060 22420 33088 22460
rect 33686 22420 33692 22432
rect 33060 22392 33692 22420
rect 33686 22380 33692 22392
rect 33744 22380 33750 22432
rect 34422 22420 34428 22432
rect 34383 22392 34428 22420
rect 34422 22380 34428 22392
rect 34480 22380 34486 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 3789 22219 3847 22225
rect 3789 22185 3801 22219
rect 3835 22216 3847 22219
rect 3878 22216 3884 22228
rect 3835 22188 3884 22216
rect 3835 22185 3847 22188
rect 3789 22179 3847 22185
rect 3878 22176 3884 22188
rect 3936 22176 3942 22228
rect 17310 22216 17316 22228
rect 16951 22188 17316 22216
rect 2774 22108 2780 22160
rect 2832 22148 2838 22160
rect 10870 22148 10876 22160
rect 2832 22120 10876 22148
rect 2832 22108 2838 22120
rect 10870 22108 10876 22120
rect 10928 22108 10934 22160
rect 16298 22108 16304 22160
rect 16356 22148 16362 22160
rect 16951 22148 16979 22188
rect 17310 22176 17316 22188
rect 17368 22216 17374 22228
rect 17770 22216 17776 22228
rect 17368 22188 17632 22216
rect 17731 22188 17776 22216
rect 17368 22176 17374 22188
rect 16356 22120 16979 22148
rect 17604 22148 17632 22188
rect 17770 22176 17776 22188
rect 17828 22176 17834 22228
rect 25498 22216 25504 22228
rect 20456 22188 22094 22216
rect 25459 22188 25504 22216
rect 17604 22120 18000 22148
rect 16356 22108 16362 22120
rect 2041 22083 2099 22089
rect 2041 22049 2053 22083
rect 2087 22080 2099 22083
rect 15654 22080 15660 22092
rect 2087 22052 15660 22080
rect 2087 22049 2099 22052
rect 2041 22043 2099 22049
rect 15654 22040 15660 22052
rect 15712 22040 15718 22092
rect 15749 22083 15807 22089
rect 15749 22049 15761 22083
rect 15795 22080 15807 22083
rect 15838 22080 15844 22092
rect 15795 22052 15844 22080
rect 15795 22049 15807 22052
rect 15749 22043 15807 22049
rect 15838 22040 15844 22052
rect 15896 22040 15902 22092
rect 15930 22040 15936 22092
rect 15988 22080 15994 22092
rect 16117 22083 16175 22089
rect 15988 22052 16033 22080
rect 15988 22040 15994 22052
rect 16117 22049 16129 22083
rect 16163 22080 16175 22083
rect 16574 22080 16580 22092
rect 16163 22052 16580 22080
rect 16163 22049 16175 22052
rect 16117 22043 16175 22049
rect 16574 22040 16580 22052
rect 16632 22040 16638 22092
rect 16951 22089 16979 22120
rect 16946 22083 17004 22089
rect 16946 22049 16958 22083
rect 16992 22049 17004 22083
rect 17218 22080 17224 22092
rect 17179 22052 17224 22080
rect 16946 22043 17004 22049
rect 17218 22040 17224 22052
rect 17276 22040 17282 22092
rect 17972 22089 18000 22120
rect 19978 22108 19984 22160
rect 20036 22148 20042 22160
rect 20456 22148 20484 22188
rect 20036 22120 20484 22148
rect 22066 22148 22094 22188
rect 25498 22176 25504 22188
rect 25556 22176 25562 22228
rect 25682 22216 25688 22228
rect 25643 22188 25688 22216
rect 25682 22176 25688 22188
rect 25740 22176 25746 22228
rect 25774 22176 25780 22228
rect 25832 22216 25838 22228
rect 26142 22216 26148 22228
rect 25832 22188 26148 22216
rect 25832 22176 25838 22188
rect 26142 22176 26148 22188
rect 26200 22216 26206 22228
rect 29730 22216 29736 22228
rect 26200 22188 29736 22216
rect 26200 22176 26206 22188
rect 29730 22176 29736 22188
rect 29788 22176 29794 22228
rect 30834 22216 30840 22228
rect 30795 22188 30840 22216
rect 30834 22176 30840 22188
rect 30892 22176 30898 22228
rect 33229 22219 33287 22225
rect 33229 22185 33241 22219
rect 33275 22216 33287 22219
rect 33502 22216 33508 22228
rect 33275 22188 33508 22216
rect 33275 22185 33287 22188
rect 33229 22179 33287 22185
rect 33502 22176 33508 22188
rect 33560 22176 33566 22228
rect 22066 22120 22508 22148
rect 20036 22108 20042 22120
rect 18156 22089 18276 22094
rect 17957 22083 18015 22089
rect 17957 22049 17969 22083
rect 18003 22049 18015 22083
rect 17957 22043 18015 22049
rect 18141 22083 18276 22089
rect 18141 22049 18153 22083
rect 18187 22080 18276 22083
rect 20346 22080 20352 22092
rect 18187 22066 20352 22080
rect 18187 22049 18199 22066
rect 18248 22052 20352 22066
rect 18141 22043 18199 22049
rect 20346 22040 20352 22052
rect 20404 22040 20410 22092
rect 20456 22089 20484 22120
rect 20441 22083 20499 22089
rect 20441 22049 20453 22083
rect 20487 22049 20499 22083
rect 22480 22080 22508 22120
rect 29638 22080 29644 22092
rect 22480 22052 22600 22080
rect 29599 22052 29644 22080
rect 20441 22043 20499 22049
rect 1854 22012 1860 22024
rect 1815 21984 1860 22012
rect 1854 21972 1860 21984
rect 1912 21972 1918 22024
rect 2498 21972 2504 22024
rect 2556 22012 2562 22024
rect 2869 22015 2927 22021
rect 2869 22012 2881 22015
rect 2556 21984 2881 22012
rect 2556 21972 2562 21984
rect 2869 21981 2881 21984
rect 2915 21981 2927 22015
rect 3970 22012 3976 22024
rect 3931 21984 3976 22012
rect 2869 21975 2927 21981
rect 3970 21972 3976 21984
rect 4028 21972 4034 22024
rect 11333 22015 11391 22021
rect 11333 21981 11345 22015
rect 11379 22012 11391 22015
rect 11514 22012 11520 22024
rect 11379 21984 11520 22012
rect 11379 21981 11391 21984
rect 11333 21975 11391 21981
rect 11514 21972 11520 21984
rect 11572 21972 11578 22024
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 21981 11667 22015
rect 16025 22015 16083 22021
rect 16025 22012 16037 22015
rect 11609 21975 11667 21981
rect 15948 21984 16037 22012
rect 11238 21904 11244 21956
rect 11296 21944 11302 21956
rect 11624 21944 11652 21975
rect 15948 21956 15976 21984
rect 16025 21981 16037 21984
rect 16071 21981 16083 22015
rect 16025 21975 16083 21981
rect 16206 21972 16212 22024
rect 16264 22012 16270 22024
rect 17034 22012 17040 22024
rect 16264 21984 16309 22012
rect 16995 21984 17040 22012
rect 16264 21972 16270 21984
rect 17034 21972 17040 21984
rect 17092 21972 17098 22024
rect 17129 22015 17187 22021
rect 17129 21981 17141 22015
rect 17175 21981 17187 22015
rect 18046 22012 18052 22024
rect 18007 21984 18052 22012
rect 17129 21975 17187 21981
rect 11296 21916 11652 21944
rect 11296 21904 11302 21916
rect 15930 21904 15936 21956
rect 15988 21904 15994 21956
rect 17144 21944 17172 21975
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 18230 22012 18236 22024
rect 18191 21984 18236 22012
rect 18230 21972 18236 21984
rect 18288 22012 18294 22024
rect 18598 22012 18604 22024
rect 18288 21984 18604 22012
rect 18288 21972 18294 21984
rect 18598 21972 18604 21984
rect 18656 21972 18662 22024
rect 18690 21972 18696 22024
rect 18748 22012 18754 22024
rect 22462 22012 22468 22024
rect 18748 21984 22094 22012
rect 22375 21984 22468 22012
rect 18748 21972 18754 21984
rect 20708 21947 20766 21953
rect 17144 21916 20392 21944
rect 2682 21876 2688 21888
rect 2643 21848 2688 21876
rect 2682 21836 2688 21848
rect 2740 21836 2746 21888
rect 16761 21879 16819 21885
rect 16761 21845 16773 21879
rect 16807 21876 16819 21879
rect 17218 21876 17224 21888
rect 16807 21848 17224 21876
rect 16807 21845 16819 21848
rect 16761 21839 16819 21845
rect 17218 21836 17224 21848
rect 17276 21836 17282 21888
rect 20364 21876 20392 21916
rect 20708 21913 20720 21947
rect 20754 21944 20766 21947
rect 21726 21944 21732 21956
rect 20754 21916 21732 21944
rect 20754 21913 20766 21916
rect 20708 21907 20766 21913
rect 21726 21904 21732 21916
rect 21784 21904 21790 21956
rect 22066 21944 22094 21984
rect 22462 21972 22468 21984
rect 22520 22012 22526 22024
rect 22572 22012 22600 22052
rect 29638 22040 29644 22052
rect 29696 22040 29702 22092
rect 31113 22083 31171 22089
rect 31113 22049 31125 22083
rect 31159 22080 31171 22083
rect 32217 22083 32275 22089
rect 32217 22080 32229 22083
rect 31159 22052 32229 22080
rect 31159 22049 31171 22052
rect 31113 22043 31171 22049
rect 32217 22049 32229 22052
rect 32263 22049 32275 22083
rect 32217 22043 32275 22049
rect 32490 22040 32496 22092
rect 32548 22080 32554 22092
rect 32861 22083 32919 22089
rect 32861 22080 32873 22083
rect 32548 22052 32873 22080
rect 32548 22040 32554 22052
rect 32861 22049 32873 22052
rect 32907 22049 32919 22083
rect 32861 22043 32919 22049
rect 23106 22012 23112 22024
rect 22520 21984 23112 22012
rect 22520 21972 22526 21984
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 22732 21947 22790 21953
rect 22066 21916 22692 21944
rect 21821 21879 21879 21885
rect 21821 21876 21833 21879
rect 20364 21848 21833 21876
rect 21821 21845 21833 21848
rect 21867 21876 21879 21879
rect 22186 21876 22192 21888
rect 21867 21848 22192 21876
rect 21867 21845 21879 21848
rect 21821 21839 21879 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 22664 21876 22692 21916
rect 22732 21913 22744 21947
rect 22778 21944 22790 21947
rect 24397 21947 24455 21953
rect 24397 21944 24409 21947
rect 22778 21916 24409 21944
rect 22778 21913 22790 21916
rect 22732 21907 22790 21913
rect 24397 21913 24409 21916
rect 24443 21913 24455 21947
rect 24596 21944 24624 21975
rect 24670 21972 24676 22024
rect 24728 22012 24734 22024
rect 24857 22015 24915 22021
rect 24857 22012 24869 22015
rect 24728 21984 24869 22012
rect 24728 21972 24734 21984
rect 24857 21981 24869 21984
rect 24903 22012 24915 22015
rect 25038 22012 25044 22024
rect 24903 21984 25044 22012
rect 24903 21981 24915 21984
rect 24857 21975 24915 21981
rect 25038 21972 25044 21984
rect 25096 21972 25102 22024
rect 29549 22015 29607 22021
rect 29549 21981 29561 22015
rect 29595 21981 29607 22015
rect 29730 22012 29736 22024
rect 29691 21984 29736 22012
rect 29549 21975 29607 21981
rect 25130 21944 25136 21956
rect 24596 21916 25136 21944
rect 24397 21907 24455 21913
rect 25130 21904 25136 21916
rect 25188 21904 25194 21956
rect 25317 21947 25375 21953
rect 25317 21913 25329 21947
rect 25363 21913 25375 21947
rect 29564 21944 29592 21975
rect 29730 21972 29736 21984
rect 29788 21972 29794 22024
rect 31018 22012 31024 22024
rect 30979 21984 31024 22012
rect 31018 21972 31024 21984
rect 31076 21972 31082 22024
rect 31202 22012 31208 22024
rect 31163 21984 31208 22012
rect 31202 21972 31208 21984
rect 31260 21972 31266 22024
rect 31294 21972 31300 22024
rect 31352 22012 31358 22024
rect 32953 22015 33011 22021
rect 31352 21984 31397 22012
rect 31352 21972 31358 21984
rect 32953 21981 32965 22015
rect 32999 22012 33011 22015
rect 33502 22012 33508 22024
rect 32999 21984 33508 22012
rect 32999 21981 33011 21984
rect 32953 21975 33011 21981
rect 33502 21972 33508 21984
rect 33560 22012 33566 22024
rect 34422 22012 34428 22024
rect 33560 21984 34428 22012
rect 33560 21972 33566 21984
rect 34422 21972 34428 21984
rect 34480 21972 34486 22024
rect 30098 21944 30104 21956
rect 29564 21916 30104 21944
rect 25317 21907 25375 21913
rect 23845 21879 23903 21885
rect 23845 21876 23857 21879
rect 22664 21848 23857 21876
rect 23845 21845 23857 21848
rect 23891 21876 23903 21879
rect 24765 21879 24823 21885
rect 24765 21876 24777 21879
rect 23891 21848 24777 21876
rect 23891 21845 23903 21848
rect 23845 21839 23903 21845
rect 24765 21845 24777 21848
rect 24811 21845 24823 21879
rect 24765 21839 24823 21845
rect 25038 21836 25044 21888
rect 25096 21876 25102 21888
rect 25332 21876 25360 21907
rect 30098 21904 30104 21916
rect 30156 21944 30162 21956
rect 31846 21944 31852 21956
rect 30156 21916 31852 21944
rect 30156 21904 30162 21916
rect 31846 21904 31852 21916
rect 31904 21904 31910 21956
rect 31938 21904 31944 21956
rect 31996 21944 32002 21956
rect 32033 21947 32091 21953
rect 32033 21944 32045 21947
rect 31996 21916 32045 21944
rect 31996 21904 32002 21916
rect 32033 21913 32045 21916
rect 32079 21913 32091 21947
rect 32033 21907 32091 21913
rect 25096 21848 25360 21876
rect 25096 21836 25102 21848
rect 25406 21836 25412 21888
rect 25464 21876 25470 21888
rect 25517 21879 25575 21885
rect 25517 21876 25529 21879
rect 25464 21848 25529 21876
rect 25464 21836 25470 21848
rect 25517 21845 25529 21848
rect 25563 21845 25575 21879
rect 25517 21839 25575 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 7650 21672 7656 21684
rect 3988 21644 7656 21672
rect 2682 21564 2688 21616
rect 2740 21604 2746 21616
rect 2930 21607 2988 21613
rect 2930 21604 2942 21607
rect 2740 21576 2942 21604
rect 2740 21564 2746 21576
rect 2930 21573 2942 21576
rect 2976 21573 2988 21607
rect 2930 21567 2988 21573
rect 1397 21539 1455 21545
rect 1397 21505 1409 21539
rect 1443 21536 1455 21539
rect 3988 21536 4016 21644
rect 7650 21632 7656 21644
rect 7708 21632 7714 21684
rect 10870 21672 10876 21684
rect 10831 21644 10876 21672
rect 10870 21632 10876 21644
rect 10928 21632 10934 21684
rect 16850 21632 16856 21684
rect 16908 21672 16914 21684
rect 17129 21675 17187 21681
rect 17129 21672 17141 21675
rect 16908 21644 17141 21672
rect 16908 21632 16914 21644
rect 17129 21641 17141 21644
rect 17175 21641 17187 21675
rect 17129 21635 17187 21641
rect 21726 21632 21732 21684
rect 21784 21672 21790 21684
rect 21821 21675 21879 21681
rect 21821 21672 21833 21675
rect 21784 21644 21833 21672
rect 21784 21632 21790 21644
rect 21821 21641 21833 21644
rect 21867 21641 21879 21675
rect 22186 21672 22192 21684
rect 22147 21644 22192 21672
rect 21821 21635 21879 21641
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 26142 21672 26148 21684
rect 22293 21644 25912 21672
rect 26103 21644 26148 21672
rect 4890 21604 4896 21616
rect 4851 21576 4896 21604
rect 4890 21564 4896 21576
rect 4948 21564 4954 21616
rect 8294 21604 8300 21616
rect 7760 21576 8300 21604
rect 7760 21545 7788 21576
rect 8294 21564 8300 21576
rect 8352 21604 8358 21616
rect 10594 21604 10600 21616
rect 8352 21576 10600 21604
rect 8352 21564 8358 21576
rect 10594 21564 10600 21576
rect 10652 21564 10658 21616
rect 15654 21564 15660 21616
rect 15712 21604 15718 21616
rect 18046 21604 18052 21616
rect 15712 21576 18052 21604
rect 15712 21564 15718 21576
rect 18046 21564 18052 21576
rect 18104 21564 18110 21616
rect 18874 21604 18880 21616
rect 18432 21576 18880 21604
rect 5077 21539 5135 21545
rect 5077 21536 5089 21539
rect 1443 21508 4016 21536
rect 4080 21508 5089 21536
rect 1443 21505 1455 21508
rect 1397 21499 1455 21505
rect 2685 21471 2743 21477
rect 2685 21437 2697 21471
rect 2731 21437 2743 21471
rect 2685 21431 2743 21437
rect 2700 21344 2728 21431
rect 4080 21344 4108 21508
rect 5077 21505 5089 21508
rect 5123 21505 5135 21539
rect 5077 21499 5135 21505
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21505 7803 21539
rect 7745 21499 7803 21505
rect 9760 21539 9818 21545
rect 9760 21505 9772 21539
rect 9806 21536 9818 21539
rect 10134 21536 10140 21548
rect 9806 21508 10140 21536
rect 9806 21505 9818 21508
rect 9760 21499 9818 21505
rect 7484 21468 7512 21499
rect 10134 21496 10140 21508
rect 10192 21496 10198 21548
rect 13814 21496 13820 21548
rect 13872 21536 13878 21548
rect 14093 21539 14151 21545
rect 14093 21536 14105 21539
rect 13872 21508 14105 21536
rect 13872 21496 13878 21508
rect 14093 21505 14105 21508
rect 14139 21536 14151 21539
rect 14366 21536 14372 21548
rect 14139 21508 14372 21536
rect 14139 21505 14151 21508
rect 14093 21499 14151 21505
rect 14366 21496 14372 21508
rect 14424 21536 14430 21548
rect 15746 21536 15752 21548
rect 14424 21508 15752 21536
rect 14424 21496 14430 21508
rect 15746 21496 15752 21508
rect 15804 21496 15810 21548
rect 17218 21496 17224 21548
rect 17276 21536 17282 21548
rect 17313 21539 17371 21545
rect 17313 21536 17325 21539
rect 17276 21508 17325 21536
rect 17276 21496 17282 21508
rect 17313 21505 17325 21508
rect 17359 21505 17371 21539
rect 17313 21499 17371 21505
rect 17405 21539 17463 21545
rect 17405 21505 17417 21539
rect 17451 21536 17463 21539
rect 17954 21536 17960 21548
rect 17451 21508 17960 21536
rect 17451 21505 17463 21508
rect 17405 21499 17463 21505
rect 17954 21496 17960 21508
rect 18012 21496 18018 21548
rect 18138 21496 18144 21548
rect 18196 21536 18202 21548
rect 18432 21545 18460 21576
rect 18874 21564 18880 21576
rect 18932 21564 18938 21616
rect 22094 21604 22100 21616
rect 22007 21576 22100 21604
rect 18417 21539 18475 21545
rect 18417 21536 18429 21539
rect 18196 21508 18429 21536
rect 18196 21496 18202 21508
rect 18417 21505 18429 21508
rect 18463 21505 18475 21539
rect 18417 21499 18475 21505
rect 18506 21496 18512 21548
rect 18564 21536 18570 21548
rect 22020 21545 22048 21576
rect 22094 21564 22100 21576
rect 22152 21604 22158 21616
rect 22293 21604 22321 21644
rect 22152 21576 22321 21604
rect 24765 21607 24823 21613
rect 22152 21564 22158 21576
rect 24765 21573 24777 21607
rect 24811 21573 24823 21607
rect 24946 21604 24952 21616
rect 25004 21613 25010 21616
rect 25004 21607 25039 21613
rect 24891 21576 24952 21604
rect 24765 21567 24823 21573
rect 22005 21539 22063 21545
rect 18564 21508 18609 21536
rect 18564 21496 18570 21508
rect 22005 21505 22017 21539
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 22281 21539 22339 21545
rect 22281 21505 22293 21539
rect 22327 21536 22339 21539
rect 24670 21536 24676 21548
rect 22327 21508 24676 21536
rect 22327 21505 22339 21508
rect 22281 21499 22339 21505
rect 8938 21468 8944 21480
rect 7484 21440 8944 21468
rect 8938 21428 8944 21440
rect 8996 21428 9002 21480
rect 9490 21468 9496 21480
rect 9451 21440 9496 21468
rect 9490 21428 9496 21440
rect 9548 21428 9554 21480
rect 17497 21471 17555 21477
rect 17497 21468 17509 21471
rect 17145 21440 17509 21468
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 2682 21332 2688 21344
rect 2595 21304 2688 21332
rect 2682 21292 2688 21304
rect 2740 21332 2746 21344
rect 3786 21332 3792 21344
rect 2740 21304 3792 21332
rect 2740 21292 2746 21304
rect 3786 21292 3792 21304
rect 3844 21292 3850 21344
rect 4062 21332 4068 21344
rect 4023 21304 4068 21332
rect 4062 21292 4068 21304
rect 4120 21292 4126 21344
rect 5258 21332 5264 21344
rect 5219 21304 5264 21332
rect 5258 21292 5264 21304
rect 5316 21292 5322 21344
rect 7282 21332 7288 21344
rect 7243 21304 7288 21332
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 11606 21292 11612 21344
rect 11664 21332 11670 21344
rect 14182 21332 14188 21344
rect 11664 21304 14188 21332
rect 11664 21292 11670 21304
rect 14182 21292 14188 21304
rect 14240 21292 14246 21344
rect 15930 21292 15936 21344
rect 15988 21332 15994 21344
rect 16390 21332 16396 21344
rect 15988 21304 16396 21332
rect 15988 21292 15994 21304
rect 16390 21292 16396 21304
rect 16448 21292 16454 21344
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 17145 21332 17173 21440
rect 17497 21437 17509 21440
rect 17543 21437 17555 21471
rect 17497 21431 17555 21437
rect 17586 21428 17592 21480
rect 17644 21468 17650 21480
rect 18322 21468 18328 21480
rect 17644 21440 17689 21468
rect 18283 21440 18328 21468
rect 17644 21428 17650 21440
rect 18322 21428 18328 21440
rect 18380 21428 18386 21480
rect 18598 21468 18604 21480
rect 18559 21440 18604 21468
rect 18598 21428 18604 21440
rect 18656 21428 18662 21480
rect 21174 21428 21180 21480
rect 21232 21468 21238 21480
rect 22296 21468 22324 21499
rect 24670 21496 24676 21508
rect 24728 21496 24734 21548
rect 21232 21440 22324 21468
rect 24780 21468 24808 21567
rect 24946 21564 24952 21576
rect 25027 21604 25039 21607
rect 25406 21604 25412 21616
rect 25027 21576 25412 21604
rect 25027 21573 25039 21576
rect 25004 21567 25039 21573
rect 25004 21564 25010 21567
rect 25406 21564 25412 21576
rect 25464 21564 25470 21616
rect 25777 21607 25835 21613
rect 25777 21573 25789 21607
rect 25823 21573 25835 21607
rect 25777 21567 25835 21573
rect 25038 21468 25044 21480
rect 24780 21440 25044 21468
rect 21232 21428 21238 21440
rect 25038 21428 25044 21440
rect 25096 21468 25102 21480
rect 25792 21468 25820 21567
rect 25096 21440 25820 21468
rect 25884 21468 25912 21644
rect 26142 21632 26148 21644
rect 26200 21632 26206 21684
rect 29549 21675 29607 21681
rect 29549 21641 29561 21675
rect 29595 21672 29607 21675
rect 29730 21672 29736 21684
rect 29595 21644 29736 21672
rect 29595 21641 29607 21644
rect 29549 21635 29607 21641
rect 29730 21632 29736 21644
rect 29788 21632 29794 21684
rect 31018 21632 31024 21684
rect 31076 21672 31082 21684
rect 32490 21672 32496 21684
rect 31076 21644 32496 21672
rect 31076 21632 31082 21644
rect 32490 21632 32496 21644
rect 32548 21632 32554 21684
rect 26050 21604 26056 21616
rect 25992 21573 26056 21604
rect 25992 21542 26019 21573
rect 26007 21539 26019 21542
rect 26053 21564 26056 21573
rect 26108 21564 26114 21616
rect 31294 21604 31300 21616
rect 26160 21576 31300 21604
rect 26053 21539 26065 21564
rect 26007 21533 26065 21539
rect 26160 21468 26188 21576
rect 31294 21564 31300 21576
rect 31352 21564 31358 21616
rect 31938 21564 31944 21616
rect 31996 21604 32002 21616
rect 31996 21576 32536 21604
rect 31996 21564 32002 21576
rect 27890 21545 27896 21548
rect 27884 21499 27896 21545
rect 27948 21536 27954 21548
rect 29454 21536 29460 21548
rect 27948 21508 27984 21536
rect 29415 21508 29460 21536
rect 27890 21496 27896 21499
rect 27948 21496 27954 21508
rect 29454 21496 29460 21508
rect 29512 21496 29518 21548
rect 29546 21496 29552 21548
rect 29604 21536 29610 21548
rect 29641 21539 29699 21545
rect 29641 21536 29653 21539
rect 29604 21508 29653 21536
rect 29604 21496 29610 21508
rect 29641 21505 29653 21508
rect 29687 21505 29699 21539
rect 29641 21499 29699 21505
rect 31846 21496 31852 21548
rect 31904 21536 31910 21548
rect 32508 21545 32536 21576
rect 32309 21539 32367 21545
rect 32309 21536 32321 21539
rect 31904 21508 32321 21536
rect 31904 21496 31910 21508
rect 32309 21505 32321 21508
rect 32355 21505 32367 21539
rect 32309 21499 32367 21505
rect 32493 21539 32551 21545
rect 32493 21505 32505 21539
rect 32539 21505 32551 21539
rect 32493 21499 32551 21505
rect 27614 21468 27620 21480
rect 25884 21440 26188 21468
rect 27575 21440 27620 21468
rect 25096 21428 25102 21440
rect 27614 21428 27620 21440
rect 27672 21428 27678 21480
rect 32324 21468 32352 21499
rect 34790 21496 34796 21548
rect 34848 21536 34854 21548
rect 35253 21539 35311 21545
rect 35253 21536 35265 21539
rect 34848 21508 35265 21536
rect 34848 21496 34854 21508
rect 35253 21505 35265 21508
rect 35299 21505 35311 21539
rect 35253 21499 35311 21505
rect 33318 21468 33324 21480
rect 32324 21440 33324 21468
rect 33318 21428 33324 21440
rect 33376 21428 33382 21480
rect 17218 21360 17224 21412
rect 17276 21400 17282 21412
rect 23934 21400 23940 21412
rect 17276 21372 23940 21400
rect 17276 21360 17282 21372
rect 23934 21360 23940 21372
rect 23992 21360 23998 21412
rect 25590 21400 25596 21412
rect 24964 21372 25596 21400
rect 17862 21332 17868 21344
rect 16632 21304 17868 21332
rect 16632 21292 16638 21304
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 18141 21335 18199 21341
rect 18141 21301 18153 21335
rect 18187 21332 18199 21335
rect 19426 21332 19432 21344
rect 18187 21304 19432 21332
rect 18187 21301 18199 21304
rect 18141 21295 18199 21301
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 24486 21292 24492 21344
rect 24544 21332 24550 21344
rect 24964 21341 24992 21372
rect 25590 21360 25596 21372
rect 25648 21360 25654 21412
rect 24673 21335 24731 21341
rect 24673 21332 24685 21335
rect 24544 21304 24685 21332
rect 24544 21292 24550 21304
rect 24673 21301 24685 21304
rect 24719 21332 24731 21335
rect 24949 21335 25007 21341
rect 24949 21332 24961 21335
rect 24719 21304 24961 21332
rect 24719 21301 24731 21304
rect 24673 21295 24731 21301
rect 24949 21301 24961 21304
rect 24995 21301 25007 21335
rect 25130 21332 25136 21344
rect 25091 21304 25136 21332
rect 24949 21295 25007 21301
rect 25130 21292 25136 21304
rect 25188 21292 25194 21344
rect 25314 21292 25320 21344
rect 25372 21332 25378 21344
rect 25501 21335 25559 21341
rect 25501 21332 25513 21335
rect 25372 21304 25513 21332
rect 25372 21292 25378 21304
rect 25501 21301 25513 21304
rect 25547 21332 25559 21335
rect 25866 21332 25872 21344
rect 25547 21304 25872 21332
rect 25547 21301 25559 21304
rect 25501 21295 25559 21301
rect 25866 21292 25872 21304
rect 25924 21332 25930 21344
rect 25961 21335 26019 21341
rect 25961 21332 25973 21335
rect 25924 21304 25973 21332
rect 25924 21292 25930 21304
rect 25961 21301 25973 21304
rect 26007 21301 26019 21335
rect 25961 21295 26019 21301
rect 28997 21335 29055 21341
rect 28997 21301 29009 21335
rect 29043 21332 29055 21335
rect 29178 21332 29184 21344
rect 29043 21304 29184 21332
rect 29043 21301 29055 21304
rect 28997 21295 29055 21301
rect 29178 21292 29184 21304
rect 29236 21292 29242 21344
rect 35069 21335 35127 21341
rect 35069 21301 35081 21335
rect 35115 21332 35127 21335
rect 35434 21332 35440 21344
rect 35115 21304 35440 21332
rect 35115 21301 35127 21304
rect 35069 21295 35127 21301
rect 35434 21292 35440 21304
rect 35492 21292 35498 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 2498 21128 2504 21140
rect 2459 21100 2504 21128
rect 2498 21088 2504 21100
rect 2556 21088 2562 21140
rect 7650 21128 7656 21140
rect 2746 21100 7236 21128
rect 7611 21100 7656 21128
rect 1949 21063 2007 21069
rect 1949 21029 1961 21063
rect 1995 21060 2007 21063
rect 2746 21060 2774 21100
rect 1995 21032 2774 21060
rect 7208 21060 7236 21100
rect 7650 21088 7656 21100
rect 7708 21088 7714 21140
rect 10134 21128 10140 21140
rect 10095 21100 10140 21128
rect 10134 21088 10140 21100
rect 10192 21088 10198 21140
rect 17218 21128 17224 21140
rect 12406 21100 17224 21128
rect 12406 21060 12434 21100
rect 17218 21088 17224 21100
rect 17276 21088 17282 21140
rect 17954 21088 17960 21140
rect 18012 21128 18018 21140
rect 18690 21128 18696 21140
rect 18012 21100 18696 21128
rect 18012 21088 18018 21100
rect 18690 21088 18696 21100
rect 18748 21088 18754 21140
rect 19242 21128 19248 21140
rect 19203 21100 19248 21128
rect 19242 21088 19248 21100
rect 19300 21088 19306 21140
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 27890 21128 27896 21140
rect 19392 21100 19748 21128
rect 27851 21100 27896 21128
rect 19392 21088 19398 21100
rect 7208 21032 12434 21060
rect 1995 21029 2007 21032
rect 1949 21023 2007 21029
rect 13446 21020 13452 21072
rect 13504 21060 13510 21072
rect 15105 21063 15163 21069
rect 15105 21060 15117 21063
rect 13504 21032 15117 21060
rect 13504 21020 13510 21032
rect 15105 21029 15117 21032
rect 15151 21029 15163 21063
rect 16482 21060 16488 21072
rect 15105 21023 15163 21029
rect 15396 21032 16488 21060
rect 2958 20992 2964 21004
rect 2919 20964 2964 20992
rect 2958 20952 2964 20964
rect 3016 20952 3022 21004
rect 3142 20992 3148 21004
rect 3103 20964 3148 20992
rect 3142 20952 3148 20964
rect 3200 20952 3206 21004
rect 13170 20992 13176 21004
rect 10336 20964 13176 20992
rect 2869 20927 2927 20933
rect 2869 20893 2881 20927
rect 2915 20924 2927 20927
rect 4062 20924 4068 20936
rect 2915 20896 4068 20924
rect 2915 20893 2927 20896
rect 2869 20887 2927 20893
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 6273 20927 6331 20933
rect 6273 20893 6285 20927
rect 6319 20893 6331 20927
rect 6273 20887 6331 20893
rect 6540 20927 6598 20933
rect 6540 20893 6552 20927
rect 6586 20924 6598 20927
rect 7282 20924 7288 20936
rect 6586 20896 7288 20924
rect 6586 20893 6598 20896
rect 6540 20887 6598 20893
rect 1670 20856 1676 20868
rect 1631 20828 1676 20856
rect 1670 20816 1676 20828
rect 1728 20816 1734 20868
rect 6288 20856 6316 20887
rect 7282 20884 7288 20896
rect 7340 20884 7346 20936
rect 10336 20933 10364 20964
rect 13170 20952 13176 20964
rect 13228 20952 13234 21004
rect 14461 20995 14519 21001
rect 14461 20961 14473 20995
rect 14507 20992 14519 20995
rect 14642 20992 14648 21004
rect 14507 20964 14648 20992
rect 14507 20961 14519 20964
rect 14461 20955 14519 20961
rect 14642 20952 14648 20964
rect 14700 20952 14706 21004
rect 15396 21001 15424 21032
rect 16482 21020 16488 21032
rect 16540 21020 16546 21072
rect 17126 21020 17132 21072
rect 17184 21060 17190 21072
rect 17773 21063 17831 21069
rect 17773 21060 17785 21063
rect 17184 21032 17785 21060
rect 17184 21020 17190 21032
rect 17773 21029 17785 21032
rect 17819 21029 17831 21063
rect 17773 21023 17831 21029
rect 17862 21020 17868 21072
rect 17920 21060 17926 21072
rect 17920 21032 19656 21060
rect 17920 21020 17926 21032
rect 15381 20995 15439 21001
rect 15381 20961 15393 20995
rect 15427 20961 15439 20995
rect 15381 20955 15439 20961
rect 15473 20995 15531 21001
rect 15473 20961 15485 20995
rect 15519 20992 15531 20995
rect 16574 20992 16580 21004
rect 15519 20964 16580 20992
rect 15519 20961 15531 20964
rect 15473 20955 15531 20961
rect 16574 20952 16580 20964
rect 16632 20952 16638 21004
rect 17586 20952 17592 21004
rect 17644 20992 17650 21004
rect 18141 20995 18199 21001
rect 18141 20992 18153 20995
rect 17644 20964 18153 20992
rect 17644 20952 17650 20964
rect 18141 20961 18153 20964
rect 18187 20961 18199 20995
rect 19426 20992 19432 21004
rect 19387 20964 19432 20992
rect 18141 20955 18199 20961
rect 19426 20952 19432 20964
rect 19484 20952 19490 21004
rect 19628 21001 19656 21032
rect 19720 21001 19748 21100
rect 27890 21088 27896 21100
rect 27948 21088 27954 21140
rect 36541 21131 36599 21137
rect 36541 21128 36553 21131
rect 33612 21100 36553 21128
rect 19794 21020 19800 21072
rect 19852 21060 19858 21072
rect 30190 21060 30196 21072
rect 19852 21032 30196 21060
rect 19852 21020 19858 21032
rect 30190 21020 30196 21032
rect 30248 21020 30254 21072
rect 33612 21004 33640 21100
rect 36541 21097 36553 21100
rect 36587 21097 36599 21131
rect 36541 21091 36599 21097
rect 33686 21020 33692 21072
rect 33744 21060 33750 21072
rect 33744 21032 35204 21060
rect 33744 21020 33750 21032
rect 19613 20995 19671 21001
rect 19613 20961 19625 20995
rect 19659 20961 19671 20995
rect 19613 20955 19671 20961
rect 19705 20995 19763 21001
rect 19705 20961 19717 20995
rect 19751 20961 19763 20995
rect 19705 20955 19763 20961
rect 31938 20952 31944 21004
rect 31996 20992 32002 21004
rect 33042 20992 33048 21004
rect 31996 20964 33048 20992
rect 31996 20952 32002 20964
rect 33042 20952 33048 20964
rect 33100 20992 33106 21004
rect 33413 20995 33471 21001
rect 33413 20992 33425 20995
rect 33100 20964 33425 20992
rect 33100 20952 33106 20964
rect 33413 20961 33425 20964
rect 33459 20961 33471 20995
rect 33413 20955 33471 20961
rect 33594 20952 33600 21004
rect 33652 20992 33658 21004
rect 35176 21001 35204 21032
rect 35161 20995 35219 21001
rect 33652 20964 33745 20992
rect 33652 20952 33658 20964
rect 35161 20961 35173 20995
rect 35207 20961 35219 20995
rect 35161 20955 35219 20961
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20893 10379 20927
rect 10594 20924 10600 20936
rect 10507 20896 10600 20924
rect 10321 20887 10379 20893
rect 10594 20884 10600 20896
rect 10652 20924 10658 20936
rect 10652 20896 11468 20924
rect 10652 20884 10658 20896
rect 7098 20856 7104 20868
rect 6288 20828 7104 20856
rect 7098 20816 7104 20828
rect 7156 20816 7162 20868
rect 10505 20859 10563 20865
rect 10505 20825 10517 20859
rect 10551 20856 10563 20859
rect 10870 20856 10876 20868
rect 10551 20828 10876 20856
rect 10551 20825 10563 20828
rect 10505 20819 10563 20825
rect 10870 20816 10876 20828
rect 10928 20816 10934 20868
rect 11440 20856 11468 20896
rect 11514 20884 11520 20936
rect 11572 20924 11578 20936
rect 11793 20927 11851 20933
rect 11793 20924 11805 20927
rect 11572 20896 11805 20924
rect 11572 20884 11578 20896
rect 11793 20893 11805 20896
rect 11839 20893 11851 20927
rect 11793 20887 11851 20893
rect 13265 20927 13323 20933
rect 13265 20893 13277 20927
rect 13311 20924 13323 20927
rect 13354 20924 13360 20936
rect 13311 20896 13360 20924
rect 13311 20893 13323 20896
rect 13265 20887 13323 20893
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 13538 20924 13544 20936
rect 13499 20896 13544 20924
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 14274 20924 14280 20936
rect 14235 20896 14280 20924
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 14366 20884 14372 20936
rect 14424 20924 14430 20936
rect 14553 20927 14611 20933
rect 14424 20896 14469 20924
rect 14424 20884 14430 20896
rect 14553 20893 14565 20927
rect 14599 20924 14611 20927
rect 15286 20924 15292 20936
rect 14599 20896 15148 20924
rect 15247 20896 15292 20924
rect 14599 20893 14611 20896
rect 14553 20887 14611 20893
rect 13630 20856 13636 20868
rect 11440 20828 13636 20856
rect 13630 20816 13636 20828
rect 13688 20816 13694 20868
rect 15120 20856 15148 20896
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 15562 20924 15568 20936
rect 15523 20896 15568 20924
rect 15562 20884 15568 20896
rect 15620 20884 15626 20936
rect 17954 20924 17960 20936
rect 17915 20896 17960 20924
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 18049 20927 18107 20933
rect 18049 20893 18061 20927
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 15930 20856 15936 20868
rect 15120 20828 15936 20856
rect 15930 20816 15936 20828
rect 15988 20816 15994 20868
rect 18064 20856 18092 20887
rect 18230 20884 18236 20936
rect 18288 20924 18294 20936
rect 19334 20924 19340 20936
rect 18288 20896 19340 20924
rect 18288 20884 18294 20896
rect 19334 20884 19340 20896
rect 19392 20884 19398 20936
rect 19518 20884 19524 20936
rect 19576 20924 19582 20936
rect 19576 20896 19621 20924
rect 19576 20884 19582 20896
rect 25130 20884 25136 20936
rect 25188 20924 25194 20936
rect 28077 20927 28135 20933
rect 28077 20924 28089 20927
rect 25188 20896 28089 20924
rect 25188 20884 25194 20896
rect 28077 20893 28089 20896
rect 28123 20893 28135 20927
rect 28077 20887 28135 20893
rect 28166 20884 28172 20936
rect 28224 20924 28230 20936
rect 28261 20927 28319 20933
rect 28261 20924 28273 20927
rect 28224 20896 28273 20924
rect 28224 20884 28230 20896
rect 28261 20893 28273 20896
rect 28307 20893 28319 20927
rect 28261 20887 28319 20893
rect 28353 20927 28411 20933
rect 28353 20893 28365 20927
rect 28399 20893 28411 20927
rect 28353 20887 28411 20893
rect 28368 20856 28396 20887
rect 28534 20884 28540 20936
rect 28592 20924 28598 20936
rect 28813 20927 28871 20933
rect 28813 20924 28825 20927
rect 28592 20896 28825 20924
rect 28592 20884 28598 20896
rect 28813 20893 28825 20896
rect 28859 20893 28871 20927
rect 28813 20887 28871 20893
rect 28997 20927 29055 20933
rect 28997 20893 29009 20927
rect 29043 20924 29055 20927
rect 29086 20924 29092 20936
rect 29043 20896 29092 20924
rect 29043 20893 29055 20896
rect 28997 20887 29055 20893
rect 29086 20884 29092 20896
rect 29144 20924 29150 20936
rect 29454 20924 29460 20936
rect 29144 20896 29460 20924
rect 29144 20884 29150 20896
rect 29454 20884 29460 20896
rect 29512 20884 29518 20936
rect 33318 20924 33324 20936
rect 33231 20896 33324 20924
rect 33318 20884 33324 20896
rect 33376 20884 33382 20936
rect 33502 20884 33508 20936
rect 33560 20924 33566 20936
rect 33686 20924 33692 20936
rect 33560 20896 33692 20924
rect 33560 20884 33566 20896
rect 33686 20884 33692 20896
rect 33744 20884 33750 20936
rect 28905 20859 28963 20865
rect 28905 20856 28917 20859
rect 18064 20828 26924 20856
rect 28368 20828 28917 20856
rect 11146 20748 11152 20800
rect 11204 20788 11210 20800
rect 11977 20791 12035 20797
rect 11977 20788 11989 20791
rect 11204 20760 11989 20788
rect 11204 20748 11210 20760
rect 11977 20757 11989 20760
rect 12023 20788 12035 20791
rect 12066 20788 12072 20800
rect 12023 20760 12072 20788
rect 12023 20757 12035 20760
rect 11977 20751 12035 20757
rect 12066 20748 12072 20760
rect 12124 20748 12130 20800
rect 13078 20788 13084 20800
rect 13039 20760 13084 20788
rect 13078 20748 13084 20760
rect 13136 20748 13142 20800
rect 13446 20788 13452 20800
rect 13407 20760 13452 20788
rect 13446 20748 13452 20760
rect 13504 20748 13510 20800
rect 14093 20791 14151 20797
rect 14093 20757 14105 20791
rect 14139 20788 14151 20791
rect 14182 20788 14188 20800
rect 14139 20760 14188 20788
rect 14139 20757 14151 20760
rect 14093 20751 14151 20757
rect 14182 20748 14188 20760
rect 14240 20748 14246 20800
rect 14550 20748 14556 20800
rect 14608 20788 14614 20800
rect 25682 20788 25688 20800
rect 14608 20760 25688 20788
rect 14608 20748 14614 20760
rect 25682 20748 25688 20760
rect 25740 20748 25746 20800
rect 26896 20788 26924 20828
rect 28905 20825 28917 20828
rect 28951 20825 28963 20859
rect 28905 20819 28963 20825
rect 30374 20816 30380 20868
rect 30432 20856 30438 20868
rect 31202 20856 31208 20868
rect 30432 20828 31208 20856
rect 30432 20816 30438 20828
rect 31202 20816 31208 20828
rect 31260 20816 31266 20868
rect 31662 20816 31668 20868
rect 31720 20856 31726 20868
rect 33336 20856 33364 20884
rect 33870 20856 33876 20868
rect 31720 20828 33272 20856
rect 33336 20828 33876 20856
rect 31720 20816 31726 20828
rect 32766 20788 32772 20800
rect 26896 20760 32772 20788
rect 32766 20748 32772 20760
rect 32824 20748 32830 20800
rect 33134 20788 33140 20800
rect 33095 20760 33140 20788
rect 33134 20748 33140 20760
rect 33192 20748 33198 20800
rect 33244 20788 33272 20828
rect 33870 20816 33876 20828
rect 33928 20816 33934 20868
rect 35176 20856 35204 20955
rect 35434 20933 35440 20936
rect 35428 20924 35440 20933
rect 35395 20896 35440 20924
rect 35428 20887 35440 20896
rect 35434 20884 35440 20887
rect 35492 20884 35498 20936
rect 35710 20884 35716 20936
rect 35768 20924 35774 20936
rect 37369 20927 37427 20933
rect 37369 20924 37381 20927
rect 35768 20896 37381 20924
rect 35768 20884 35774 20896
rect 37369 20893 37381 20896
rect 37415 20893 37427 20927
rect 37642 20924 37648 20936
rect 37603 20896 37648 20924
rect 37369 20887 37427 20893
rect 37642 20884 37648 20896
rect 37700 20884 37706 20936
rect 37734 20856 37740 20868
rect 35176 20828 37740 20856
rect 37734 20816 37740 20828
rect 37792 20816 37798 20868
rect 35710 20788 35716 20800
rect 33244 20760 35716 20788
rect 35710 20748 35716 20760
rect 35768 20748 35774 20800
rect 37185 20791 37243 20797
rect 37185 20757 37197 20791
rect 37231 20788 37243 20791
rect 37366 20788 37372 20800
rect 37231 20760 37372 20788
rect 37231 20757 37243 20760
rect 37185 20751 37243 20757
rect 37366 20748 37372 20760
rect 37424 20748 37430 20800
rect 37458 20748 37464 20800
rect 37516 20788 37522 20800
rect 37553 20791 37611 20797
rect 37553 20788 37565 20791
rect 37516 20760 37565 20788
rect 37516 20748 37522 20760
rect 37553 20757 37565 20760
rect 37599 20757 37611 20791
rect 37553 20751 37611 20757
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 2961 20587 3019 20593
rect 2961 20553 2973 20587
rect 3007 20584 3019 20587
rect 3697 20587 3755 20593
rect 3697 20584 3709 20587
rect 3007 20556 3709 20584
rect 3007 20553 3019 20556
rect 2961 20547 3019 20553
rect 3697 20553 3709 20556
rect 3743 20553 3755 20587
rect 3697 20547 3755 20553
rect 8481 20587 8539 20593
rect 8481 20553 8493 20587
rect 8527 20553 8539 20587
rect 8481 20547 8539 20553
rect 8202 20516 8208 20528
rect 1412 20488 8208 20516
rect 1412 20457 1440 20488
rect 8202 20476 8208 20488
rect 8260 20516 8266 20528
rect 8496 20516 8524 20547
rect 13446 20544 13452 20596
rect 13504 20584 13510 20596
rect 14093 20587 14151 20593
rect 14093 20584 14105 20587
rect 13504 20556 14105 20584
rect 13504 20544 13510 20556
rect 14093 20553 14105 20556
rect 14139 20584 14151 20587
rect 14642 20584 14648 20596
rect 14139 20556 14648 20584
rect 14139 20553 14151 20556
rect 14093 20547 14151 20553
rect 14642 20544 14648 20556
rect 14700 20544 14706 20596
rect 15286 20544 15292 20596
rect 15344 20584 15350 20596
rect 15473 20587 15531 20593
rect 15473 20584 15485 20587
rect 15344 20556 15485 20584
rect 15344 20544 15350 20556
rect 15473 20553 15485 20556
rect 15519 20553 15531 20587
rect 16298 20584 16304 20596
rect 15473 20547 15531 20553
rect 15764 20556 16304 20584
rect 8260 20488 8524 20516
rect 12980 20519 13038 20525
rect 8260 20476 8266 20488
rect 12980 20485 12992 20519
rect 13026 20516 13038 20519
rect 13078 20516 13084 20528
rect 13026 20488 13084 20516
rect 13026 20485 13038 20488
rect 12980 20479 13038 20485
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 1397 20451 1455 20457
rect 1397 20417 1409 20451
rect 1443 20417 1455 20451
rect 1397 20411 1455 20417
rect 2869 20451 2927 20457
rect 2869 20417 2881 20451
rect 2915 20448 2927 20451
rect 3694 20448 3700 20460
rect 2915 20420 3700 20448
rect 2915 20417 2927 20420
rect 2869 20411 2927 20417
rect 3694 20408 3700 20420
rect 3752 20408 3758 20460
rect 3878 20448 3884 20460
rect 3839 20420 3884 20448
rect 3878 20408 3884 20420
rect 3936 20408 3942 20460
rect 7368 20451 7426 20457
rect 7368 20417 7380 20451
rect 7414 20448 7426 20451
rect 7834 20448 7840 20460
rect 7414 20420 7840 20448
rect 7414 20417 7426 20420
rect 7368 20411 7426 20417
rect 7834 20408 7840 20420
rect 7892 20408 7898 20460
rect 12158 20408 12164 20460
rect 12216 20448 12222 20460
rect 12342 20448 12348 20460
rect 12216 20420 12348 20448
rect 12216 20408 12222 20420
rect 12342 20408 12348 20420
rect 12400 20448 12406 20460
rect 12713 20451 12771 20457
rect 12713 20448 12725 20451
rect 12400 20420 12725 20448
rect 12400 20408 12406 20420
rect 12713 20417 12725 20420
rect 12759 20417 12771 20451
rect 12713 20411 12771 20417
rect 14274 20408 14280 20460
rect 14332 20448 14338 20460
rect 15286 20448 15292 20460
rect 14332 20420 15292 20448
rect 14332 20408 14338 20420
rect 15286 20408 15292 20420
rect 15344 20448 15350 20460
rect 15657 20451 15715 20457
rect 15657 20448 15669 20451
rect 15344 20420 15669 20448
rect 15344 20408 15350 20420
rect 15657 20417 15669 20420
rect 15703 20448 15715 20451
rect 15764 20448 15792 20556
rect 16298 20544 16304 20556
rect 16356 20544 16362 20596
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18601 20587 18659 20593
rect 18601 20584 18613 20587
rect 18012 20556 18613 20584
rect 18012 20544 18018 20556
rect 18601 20553 18613 20556
rect 18647 20553 18659 20587
rect 18601 20547 18659 20553
rect 18690 20544 18696 20596
rect 18748 20584 18754 20596
rect 33045 20587 33103 20593
rect 33045 20584 33057 20587
rect 18748 20556 33057 20584
rect 18748 20544 18754 20556
rect 33045 20553 33057 20556
rect 33091 20553 33103 20587
rect 33686 20584 33692 20596
rect 33647 20556 33692 20584
rect 33045 20547 33103 20553
rect 33686 20544 33692 20556
rect 33744 20544 33750 20596
rect 33870 20584 33876 20596
rect 33831 20556 33876 20584
rect 33870 20544 33876 20556
rect 33928 20544 33934 20596
rect 34790 20544 34796 20596
rect 34848 20584 34854 20596
rect 34885 20587 34943 20593
rect 34885 20584 34897 20587
rect 34848 20556 34897 20584
rect 34848 20544 34854 20556
rect 34885 20553 34897 20556
rect 34931 20553 34943 20587
rect 34885 20547 34943 20553
rect 23750 20516 23756 20528
rect 15856 20488 23756 20516
rect 15856 20457 15884 20488
rect 23750 20476 23756 20488
rect 23808 20516 23814 20528
rect 23808 20488 24440 20516
rect 23808 20476 23814 20488
rect 15703 20420 15792 20448
rect 15841 20451 15899 20457
rect 15703 20417 15715 20420
rect 15657 20411 15715 20417
rect 15841 20417 15853 20451
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 15988 20420 16033 20448
rect 15988 20408 15994 20420
rect 17494 20408 17500 20460
rect 17552 20448 17558 20460
rect 17589 20451 17647 20457
rect 17589 20448 17601 20451
rect 17552 20420 17601 20448
rect 17552 20408 17558 20420
rect 17589 20417 17601 20420
rect 17635 20448 17647 20451
rect 18230 20448 18236 20460
rect 17635 20420 18236 20448
rect 17635 20417 17647 20420
rect 17589 20411 17647 20417
rect 18230 20408 18236 20420
rect 18288 20408 18294 20460
rect 18786 20451 18844 20457
rect 18786 20417 18798 20451
rect 18832 20417 18844 20451
rect 18786 20411 18844 20417
rect 3142 20380 3148 20392
rect 3103 20352 3148 20380
rect 3142 20340 3148 20352
rect 3200 20340 3206 20392
rect 7098 20380 7104 20392
rect 7059 20352 7104 20380
rect 7098 20340 7104 20352
rect 7156 20340 7162 20392
rect 15746 20380 15752 20392
rect 15707 20352 15752 20380
rect 15746 20340 15752 20352
rect 15804 20340 15810 20392
rect 16942 20340 16948 20392
rect 17000 20380 17006 20392
rect 17313 20383 17371 20389
rect 17313 20380 17325 20383
rect 17000 20352 17325 20380
rect 17000 20340 17006 20352
rect 17313 20349 17325 20352
rect 17359 20349 17371 20383
rect 17313 20343 17371 20349
rect 18690 20340 18696 20392
rect 18748 20380 18754 20392
rect 18800 20380 18828 20411
rect 18874 20408 18880 20460
rect 18932 20448 18938 20460
rect 19889 20451 19947 20457
rect 18932 20420 18977 20448
rect 18932 20408 18938 20420
rect 19889 20417 19901 20451
rect 19935 20448 19947 20451
rect 19978 20448 19984 20460
rect 19935 20420 19984 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 20156 20451 20214 20457
rect 20156 20417 20168 20451
rect 20202 20448 20214 20451
rect 20714 20448 20720 20460
rect 20202 20420 20720 20448
rect 20202 20417 20214 20420
rect 20156 20411 20214 20417
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 23017 20451 23075 20457
rect 23017 20417 23029 20451
rect 23063 20448 23075 20451
rect 23106 20448 23112 20460
rect 23063 20420 23112 20448
rect 23063 20417 23075 20420
rect 23017 20411 23075 20417
rect 23106 20408 23112 20420
rect 23164 20408 23170 20460
rect 23290 20457 23296 20460
rect 23284 20411 23296 20457
rect 23348 20448 23354 20460
rect 23348 20420 23384 20448
rect 23290 20408 23296 20411
rect 23348 20408 23354 20420
rect 18966 20380 18972 20392
rect 18748 20352 18828 20380
rect 18927 20352 18972 20380
rect 18748 20340 18754 20352
rect 18966 20340 18972 20352
rect 19024 20340 19030 20392
rect 19061 20383 19119 20389
rect 19061 20349 19073 20383
rect 19107 20349 19119 20383
rect 19061 20343 19119 20349
rect 18598 20272 18604 20324
rect 18656 20312 18662 20324
rect 19076 20312 19104 20343
rect 24412 20321 24440 20488
rect 25130 20476 25136 20528
rect 25188 20516 25194 20528
rect 25225 20519 25283 20525
rect 25225 20516 25237 20519
rect 25188 20488 25237 20516
rect 25188 20476 25194 20488
rect 25225 20485 25237 20488
rect 25271 20485 25283 20519
rect 25225 20479 25283 20485
rect 25409 20519 25467 20525
rect 25409 20485 25421 20519
rect 25455 20516 25467 20519
rect 26050 20516 26056 20528
rect 25455 20488 26056 20516
rect 25455 20485 25467 20488
rect 25409 20479 25467 20485
rect 26050 20476 26056 20488
rect 26108 20476 26114 20528
rect 28442 20476 28448 20528
rect 28500 20516 28506 20528
rect 28721 20519 28779 20525
rect 28721 20516 28733 20519
rect 28500 20488 28733 20516
rect 28500 20476 28506 20488
rect 28721 20485 28733 20488
rect 28767 20485 28779 20519
rect 28721 20479 28779 20485
rect 28902 20476 28908 20528
rect 28960 20525 28966 20528
rect 28960 20519 28979 20525
rect 28967 20485 28979 20519
rect 28960 20479 28979 20485
rect 28960 20476 28966 20479
rect 32674 20476 32680 20528
rect 32732 20516 32738 20528
rect 33505 20519 33563 20525
rect 32732 20488 32777 20516
rect 32732 20476 32738 20488
rect 33505 20485 33517 20519
rect 33551 20516 33563 20519
rect 33594 20516 33600 20528
rect 33551 20488 33600 20516
rect 33551 20485 33563 20488
rect 33505 20479 33563 20485
rect 33594 20476 33600 20488
rect 33652 20476 33658 20528
rect 37366 20476 37372 20528
rect 37424 20516 37430 20528
rect 37614 20519 37672 20525
rect 37614 20516 37626 20519
rect 37424 20488 37626 20516
rect 37424 20476 37430 20488
rect 37614 20485 37626 20488
rect 37660 20485 37672 20519
rect 37614 20479 37672 20485
rect 37734 20476 37740 20528
rect 37792 20476 37798 20528
rect 25682 20448 25688 20460
rect 25595 20420 25688 20448
rect 25682 20408 25688 20420
rect 25740 20448 25746 20460
rect 31662 20448 31668 20460
rect 25740 20420 31668 20448
rect 25740 20408 25746 20420
rect 31662 20408 31668 20420
rect 31720 20408 31726 20460
rect 31754 20408 31760 20460
rect 31812 20448 31818 20460
rect 32950 20457 32956 20460
rect 32408 20451 32466 20457
rect 32408 20448 32420 20451
rect 31812 20420 32420 20448
rect 31812 20408 31818 20420
rect 32408 20417 32420 20420
rect 32454 20417 32466 20451
rect 32408 20411 32466 20417
rect 32494 20451 32552 20457
rect 32494 20417 32506 20451
rect 32540 20417 32552 20451
rect 32494 20411 32552 20417
rect 32769 20451 32827 20457
rect 32769 20417 32781 20451
rect 32815 20417 32827 20451
rect 32769 20411 32827 20417
rect 32907 20451 32956 20457
rect 32907 20417 32919 20451
rect 32953 20417 32956 20451
rect 32907 20411 32956 20417
rect 18656 20284 19104 20312
rect 24397 20315 24455 20321
rect 18656 20272 18662 20284
rect 24397 20281 24409 20315
rect 24443 20281 24455 20315
rect 24397 20275 24455 20281
rect 24486 20272 24492 20324
rect 24544 20312 24550 20324
rect 28810 20312 28816 20324
rect 24544 20284 28816 20312
rect 24544 20272 24550 20284
rect 28810 20272 28816 20284
rect 28868 20272 28874 20324
rect 29086 20312 29092 20324
rect 29047 20284 29092 20312
rect 29086 20272 29092 20284
rect 29144 20272 29150 20324
rect 32509 20312 32537 20411
rect 32784 20380 32812 20411
rect 32950 20408 32956 20411
rect 33008 20408 33014 20460
rect 33042 20408 33048 20460
rect 33100 20448 33106 20460
rect 33781 20451 33839 20457
rect 33781 20448 33793 20451
rect 33100 20420 33793 20448
rect 33100 20408 33106 20420
rect 33781 20417 33793 20420
rect 33827 20417 33839 20451
rect 34514 20448 34520 20460
rect 34475 20420 34520 20448
rect 33781 20411 33839 20417
rect 34514 20408 34520 20420
rect 34572 20408 34578 20460
rect 34698 20448 34704 20460
rect 34659 20420 34704 20448
rect 34698 20408 34704 20420
rect 34756 20408 34762 20460
rect 37752 20448 37780 20476
rect 37384 20420 37780 20448
rect 33226 20380 33232 20392
rect 32784 20352 33232 20380
rect 33226 20340 33232 20352
rect 33284 20340 33290 20392
rect 37384 20389 37412 20420
rect 37369 20383 37427 20389
rect 37369 20349 37381 20383
rect 37415 20349 37427 20383
rect 37369 20343 37427 20349
rect 33594 20312 33600 20324
rect 32509 20284 33600 20312
rect 33594 20272 33600 20284
rect 33652 20272 33658 20324
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 2501 20247 2559 20253
rect 2501 20213 2513 20247
rect 2547 20244 2559 20247
rect 2774 20244 2780 20256
rect 2547 20216 2780 20244
rect 2547 20213 2559 20216
rect 2501 20207 2559 20213
rect 2774 20204 2780 20216
rect 2832 20204 2838 20256
rect 18966 20204 18972 20256
rect 19024 20244 19030 20256
rect 21082 20244 21088 20256
rect 19024 20216 21088 20244
rect 19024 20204 19030 20216
rect 21082 20204 21088 20216
rect 21140 20244 21146 20256
rect 21269 20247 21327 20253
rect 21269 20244 21281 20247
rect 21140 20216 21281 20244
rect 21140 20204 21146 20216
rect 21269 20213 21281 20216
rect 21315 20213 21327 20247
rect 21269 20207 21327 20213
rect 21910 20204 21916 20256
rect 21968 20244 21974 20256
rect 24857 20247 24915 20253
rect 24857 20244 24869 20247
rect 21968 20216 24869 20244
rect 21968 20204 21974 20216
rect 24857 20213 24869 20216
rect 24903 20244 24915 20247
rect 25409 20247 25467 20253
rect 25409 20244 25421 20247
rect 24903 20216 25421 20244
rect 24903 20213 24915 20216
rect 24857 20207 24915 20213
rect 25409 20213 25421 20216
rect 25455 20244 25467 20247
rect 28626 20244 28632 20256
rect 25455 20216 28632 20244
rect 25455 20213 25467 20216
rect 25409 20207 25467 20213
rect 28626 20204 28632 20216
rect 28684 20204 28690 20256
rect 28902 20244 28908 20256
rect 28863 20216 28908 20244
rect 28902 20204 28908 20216
rect 28960 20204 28966 20256
rect 28994 20204 29000 20256
rect 29052 20244 29058 20256
rect 33410 20244 33416 20256
rect 29052 20216 33416 20244
rect 29052 20204 29058 20216
rect 33410 20204 33416 20216
rect 33468 20204 33474 20256
rect 34054 20244 34060 20256
rect 34015 20216 34060 20244
rect 34054 20204 34060 20216
rect 34112 20204 34118 20256
rect 38010 20204 38016 20256
rect 38068 20244 38074 20256
rect 38749 20247 38807 20253
rect 38749 20244 38761 20247
rect 38068 20216 38761 20244
rect 38068 20204 38074 20216
rect 38749 20213 38761 20216
rect 38795 20213 38807 20247
rect 38749 20207 38807 20213
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 7834 20040 7840 20052
rect 7795 20012 7840 20040
rect 7834 20000 7840 20012
rect 7892 20000 7898 20052
rect 7944 20012 17448 20040
rect 2590 19932 2596 19984
rect 2648 19972 2654 19984
rect 7944 19972 7972 20012
rect 16666 19972 16672 19984
rect 2648 19944 7972 19972
rect 8036 19944 16672 19972
rect 2648 19932 2654 19944
rect 1394 19836 1400 19848
rect 1355 19808 1400 19836
rect 1394 19796 1400 19808
rect 1452 19796 1458 19848
rect 2774 19796 2780 19848
rect 2832 19836 2838 19848
rect 5074 19836 5080 19848
rect 2832 19808 2877 19836
rect 5035 19808 5080 19836
rect 2832 19796 2838 19808
rect 5074 19796 5080 19808
rect 5132 19796 5138 19848
rect 8036 19845 8064 19944
rect 16666 19932 16672 19944
rect 16724 19932 16730 19984
rect 8110 19864 8116 19916
rect 8168 19904 8174 19916
rect 10229 19907 10287 19913
rect 10229 19904 10241 19907
rect 8168 19876 10241 19904
rect 8168 19864 8174 19876
rect 10229 19873 10241 19876
rect 10275 19904 10287 19907
rect 11422 19904 11428 19916
rect 10275 19876 11428 19904
rect 10275 19873 10287 19876
rect 10229 19867 10287 19873
rect 11422 19864 11428 19876
rect 11480 19864 11486 19916
rect 11514 19864 11520 19916
rect 11572 19904 11578 19916
rect 11977 19907 12035 19913
rect 11977 19904 11989 19907
rect 11572 19876 11989 19904
rect 11572 19864 11578 19876
rect 11977 19873 11989 19876
rect 12023 19873 12035 19907
rect 11977 19867 12035 19873
rect 8021 19839 8079 19845
rect 8021 19805 8033 19839
rect 8067 19805 8079 19839
rect 8294 19836 8300 19848
rect 8255 19808 8300 19836
rect 8021 19799 8079 19805
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 11238 19836 11244 19848
rect 8404 19808 11244 19836
rect 2038 19728 2044 19780
rect 2096 19768 2102 19780
rect 8404 19768 8432 19808
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 11701 19839 11759 19845
rect 11701 19805 11713 19839
rect 11747 19805 11759 19839
rect 11992 19836 12020 19867
rect 13538 19864 13544 19916
rect 13596 19904 13602 19916
rect 15286 19904 15292 19916
rect 13596 19876 15148 19904
rect 15247 19876 15292 19904
rect 13596 19864 13602 19876
rect 14458 19836 14464 19848
rect 11992 19808 14464 19836
rect 11701 19799 11759 19805
rect 2096 19740 8432 19768
rect 10045 19771 10103 19777
rect 2096 19728 2102 19740
rect 10045 19737 10057 19771
rect 10091 19768 10103 19771
rect 11606 19768 11612 19780
rect 10091 19740 11612 19768
rect 10091 19737 10103 19740
rect 10045 19731 10103 19737
rect 11606 19728 11612 19740
rect 11664 19728 11670 19780
rect 11716 19768 11744 19799
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 14826 19796 14832 19848
rect 14884 19836 14890 19848
rect 15013 19839 15071 19845
rect 15013 19836 15025 19839
rect 14884 19808 15025 19836
rect 14884 19796 14890 19808
rect 15013 19805 15025 19808
rect 15059 19805 15071 19839
rect 15120 19836 15148 19876
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 16574 19904 16580 19916
rect 15764 19876 16436 19904
rect 16535 19876 16580 19904
rect 15764 19836 15792 19876
rect 16298 19836 16304 19848
rect 15120 19808 15792 19836
rect 16259 19808 16304 19836
rect 15013 19799 15071 19805
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 16408 19836 16436 19876
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 16408 19808 17080 19836
rect 16942 19768 16948 19780
rect 11716 19740 16948 19768
rect 16942 19728 16948 19740
rect 17000 19728 17006 19780
rect 1581 19703 1639 19709
rect 1581 19669 1593 19703
rect 1627 19700 1639 19703
rect 1762 19700 1768 19712
rect 1627 19672 1768 19700
rect 1627 19669 1639 19672
rect 1581 19663 1639 19669
rect 1762 19660 1768 19672
rect 1820 19660 1826 19712
rect 2590 19700 2596 19712
rect 2551 19672 2596 19700
rect 2590 19660 2596 19672
rect 2648 19660 2654 19712
rect 4890 19700 4896 19712
rect 4851 19672 4896 19700
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 8202 19700 8208 19712
rect 8163 19672 8208 19700
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 9674 19700 9680 19712
rect 9635 19672 9680 19700
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 9766 19660 9772 19712
rect 9824 19700 9830 19712
rect 10137 19703 10195 19709
rect 10137 19700 10149 19703
rect 9824 19672 10149 19700
rect 9824 19660 9830 19672
rect 10137 19669 10149 19672
rect 10183 19669 10195 19703
rect 10137 19663 10195 19669
rect 11238 19660 11244 19712
rect 11296 19700 11302 19712
rect 15746 19700 15752 19712
rect 11296 19672 15752 19700
rect 11296 19660 11302 19672
rect 15746 19660 15752 19672
rect 15804 19660 15810 19712
rect 17052 19700 17080 19808
rect 17420 19768 17448 20012
rect 18322 20000 18328 20052
rect 18380 20040 18386 20052
rect 18690 20040 18696 20052
rect 18380 20012 18696 20040
rect 18380 20000 18386 20012
rect 18690 20000 18696 20012
rect 18748 20040 18754 20052
rect 18874 20040 18880 20052
rect 18748 20012 18880 20040
rect 18748 20000 18754 20012
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 20714 20040 20720 20052
rect 20675 20012 20720 20040
rect 20714 20000 20720 20012
rect 20772 20000 20778 20052
rect 21450 20000 21456 20052
rect 21508 20040 21514 20052
rect 22002 20040 22008 20052
rect 21508 20012 22008 20040
rect 21508 20000 21514 20012
rect 22002 20000 22008 20012
rect 22060 20000 22066 20052
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 22189 20043 22247 20049
rect 22189 20040 22201 20043
rect 22152 20012 22201 20040
rect 22152 20000 22158 20012
rect 22189 20009 22201 20012
rect 22235 20009 22247 20043
rect 22189 20003 22247 20009
rect 23290 20000 23296 20052
rect 23348 20040 23354 20052
rect 23385 20043 23443 20049
rect 23385 20040 23397 20043
rect 23348 20012 23397 20040
rect 23348 20000 23354 20012
rect 23385 20009 23397 20012
rect 23431 20009 23443 20043
rect 23385 20003 23443 20009
rect 24670 20000 24676 20052
rect 24728 20040 24734 20052
rect 24949 20043 25007 20049
rect 24949 20040 24961 20043
rect 24728 20012 24961 20040
rect 24728 20000 24734 20012
rect 24949 20009 24961 20012
rect 24995 20009 25007 20043
rect 24949 20003 25007 20009
rect 26528 20012 27476 20040
rect 17678 19932 17684 19984
rect 17736 19972 17742 19984
rect 26528 19972 26556 20012
rect 17736 19944 26556 19972
rect 27448 19972 27476 20012
rect 28534 20000 28540 20052
rect 28592 20040 28598 20052
rect 28629 20043 28687 20049
rect 28629 20040 28641 20043
rect 28592 20012 28641 20040
rect 28592 20000 28598 20012
rect 28629 20009 28641 20012
rect 28675 20009 28687 20043
rect 28629 20003 28687 20009
rect 28810 20000 28816 20052
rect 28868 20040 28874 20052
rect 30098 20040 30104 20052
rect 28868 20012 29132 20040
rect 30059 20012 30104 20040
rect 28868 20000 28874 20012
rect 28994 19972 29000 19984
rect 27448 19944 29000 19972
rect 17736 19932 17742 19944
rect 28994 19932 29000 19944
rect 29052 19932 29058 19984
rect 29104 19972 29132 20012
rect 30098 20000 30104 20012
rect 30156 20000 30162 20052
rect 30190 20000 30196 20052
rect 30248 20040 30254 20052
rect 32401 20043 32459 20049
rect 32401 20040 32413 20043
rect 30248 20012 32413 20040
rect 30248 20000 30254 20012
rect 32401 20009 32413 20012
rect 32447 20009 32459 20043
rect 32401 20003 32459 20009
rect 33410 20000 33416 20052
rect 33468 20040 33474 20052
rect 33505 20043 33563 20049
rect 33505 20040 33517 20043
rect 33468 20012 33517 20040
rect 33468 20000 33474 20012
rect 33505 20009 33517 20012
rect 33551 20009 33563 20043
rect 33505 20003 33563 20009
rect 37001 20043 37059 20049
rect 37001 20009 37013 20043
rect 37047 20040 37059 20043
rect 37458 20040 37464 20052
rect 37047 20012 37464 20040
rect 37047 20009 37059 20012
rect 37001 20003 37059 20009
rect 37458 20000 37464 20012
rect 37516 20000 37522 20052
rect 37553 20043 37611 20049
rect 37553 20009 37565 20043
rect 37599 20040 37611 20043
rect 37642 20040 37648 20052
rect 37599 20012 37648 20040
rect 37599 20009 37611 20012
rect 37553 20003 37611 20009
rect 37642 20000 37648 20012
rect 37700 20000 37706 20052
rect 34698 19972 34704 19984
rect 29104 19944 34704 19972
rect 34698 19932 34704 19944
rect 34756 19932 34762 19984
rect 18046 19864 18052 19916
rect 18104 19904 18110 19916
rect 20714 19904 20720 19916
rect 18104 19876 20720 19904
rect 18104 19864 18110 19876
rect 20714 19864 20720 19876
rect 20772 19864 20778 19916
rect 22186 19904 22192 19916
rect 20916 19876 22192 19904
rect 17494 19796 17500 19848
rect 17552 19836 17558 19848
rect 17589 19839 17647 19845
rect 17589 19836 17601 19839
rect 17552 19808 17601 19836
rect 17552 19796 17558 19808
rect 17589 19805 17601 19808
rect 17635 19805 17647 19839
rect 17589 19799 17647 19805
rect 17865 19839 17923 19845
rect 17865 19805 17877 19839
rect 17911 19836 17923 19839
rect 18598 19836 18604 19848
rect 17911 19808 18604 19836
rect 17911 19805 17923 19808
rect 17865 19799 17923 19805
rect 18598 19796 18604 19808
rect 18656 19796 18662 19848
rect 20916 19845 20944 19876
rect 22186 19864 22192 19876
rect 22244 19864 22250 19916
rect 23658 19904 23664 19916
rect 23571 19876 23664 19904
rect 20901 19839 20959 19845
rect 20901 19805 20913 19839
rect 20947 19805 20959 19839
rect 21082 19836 21088 19848
rect 21043 19808 21088 19836
rect 20901 19799 20959 19805
rect 21082 19796 21088 19808
rect 21140 19796 21146 19848
rect 21174 19796 21180 19848
rect 21232 19836 21238 19848
rect 23584 19845 23612 19876
rect 23658 19864 23664 19876
rect 23716 19904 23722 19916
rect 24486 19904 24492 19916
rect 23716 19876 24492 19904
rect 23716 19864 23722 19876
rect 24486 19864 24492 19876
rect 24544 19864 24550 19916
rect 28442 19864 28448 19916
rect 28500 19904 28506 19916
rect 29178 19904 29184 19916
rect 28500 19876 29184 19904
rect 28500 19864 28506 19876
rect 23569 19839 23627 19845
rect 21232 19808 21277 19836
rect 21232 19796 21238 19808
rect 23569 19805 23581 19839
rect 23615 19805 23627 19839
rect 23750 19836 23756 19848
rect 23711 19808 23756 19836
rect 23569 19799 23627 19805
rect 23750 19796 23756 19808
rect 23808 19796 23814 19848
rect 23842 19796 23848 19848
rect 23900 19836 23906 19848
rect 26513 19839 26571 19845
rect 23900 19808 23945 19836
rect 23900 19796 23906 19808
rect 26513 19805 26525 19839
rect 26559 19836 26571 19839
rect 27614 19836 27620 19848
rect 26559 19808 27620 19836
rect 26559 19805 26571 19808
rect 26513 19799 26571 19805
rect 27614 19796 27620 19808
rect 27672 19796 27678 19848
rect 28644 19845 28672 19876
rect 29178 19864 29184 19876
rect 29236 19904 29242 19916
rect 29730 19904 29736 19916
rect 29236 19876 29736 19904
rect 29236 19864 29242 19876
rect 29730 19864 29736 19876
rect 29788 19864 29794 19916
rect 32674 19904 32680 19916
rect 32048 19876 32680 19904
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19805 28687 19839
rect 28629 19799 28687 19805
rect 28810 19796 28816 19848
rect 28868 19836 28874 19848
rect 28905 19839 28963 19845
rect 28905 19836 28917 19839
rect 28868 19808 28917 19836
rect 28868 19796 28874 19808
rect 28905 19805 28917 19808
rect 28951 19805 28963 19839
rect 29825 19839 29883 19845
rect 29825 19836 29837 19839
rect 28905 19799 28963 19805
rect 29012 19808 29837 19836
rect 21450 19768 21456 19780
rect 17420 19740 21456 19768
rect 21450 19728 21456 19740
rect 21508 19728 21514 19780
rect 21818 19768 21824 19780
rect 21779 19740 21824 19768
rect 21818 19728 21824 19740
rect 21876 19728 21882 19780
rect 22094 19777 22100 19780
rect 22037 19771 22100 19777
rect 22037 19737 22049 19771
rect 22083 19737 22100 19771
rect 22037 19731 22100 19737
rect 22094 19728 22100 19731
rect 22152 19728 22158 19780
rect 24857 19771 24915 19777
rect 24857 19737 24869 19771
rect 24903 19737 24915 19771
rect 24857 19731 24915 19737
rect 26780 19771 26838 19777
rect 26780 19737 26792 19771
rect 26826 19768 26838 19771
rect 26970 19768 26976 19780
rect 26826 19740 26976 19768
rect 26826 19737 26838 19740
rect 26780 19731 26838 19737
rect 21726 19700 21732 19712
rect 17052 19672 21732 19700
rect 21726 19660 21732 19672
rect 21784 19660 21790 19712
rect 24210 19660 24216 19712
rect 24268 19700 24274 19712
rect 24872 19700 24900 19731
rect 26970 19728 26976 19740
rect 27028 19728 27034 19780
rect 29012 19768 29040 19808
rect 29825 19805 29837 19808
rect 29871 19805 29883 19839
rect 31754 19836 31760 19848
rect 31715 19808 31760 19836
rect 29825 19799 29883 19805
rect 31754 19796 31760 19808
rect 31812 19796 31818 19848
rect 31938 19845 31944 19848
rect 31905 19839 31944 19845
rect 31905 19805 31917 19839
rect 31905 19799 31944 19805
rect 31938 19796 31944 19799
rect 31996 19796 32002 19848
rect 32048 19845 32076 19876
rect 32033 19839 32091 19845
rect 32033 19805 32045 19839
rect 32079 19805 32091 19839
rect 32033 19799 32091 19805
rect 32263 19839 32321 19845
rect 32263 19805 32275 19839
rect 32309 19836 32321 19839
rect 32309 19808 32537 19836
rect 32309 19805 32321 19808
rect 32263 19799 32321 19805
rect 29546 19768 29552 19780
rect 28736 19740 29040 19768
rect 29507 19740 29552 19768
rect 27062 19700 27068 19712
rect 24268 19672 27068 19700
rect 24268 19660 24274 19672
rect 27062 19660 27068 19672
rect 27120 19660 27126 19712
rect 27893 19703 27951 19709
rect 27893 19669 27905 19703
rect 27939 19700 27951 19703
rect 28534 19700 28540 19712
rect 27939 19672 28540 19700
rect 27939 19669 27951 19672
rect 27893 19663 27951 19669
rect 28534 19660 28540 19672
rect 28592 19700 28598 19712
rect 28736 19700 28764 19740
rect 29546 19728 29552 19740
rect 29604 19728 29610 19780
rect 29638 19728 29644 19780
rect 29696 19768 29702 19780
rect 29917 19771 29975 19777
rect 29917 19768 29929 19771
rect 29696 19740 29929 19768
rect 29696 19728 29702 19740
rect 29917 19737 29929 19740
rect 29963 19737 29975 19771
rect 29917 19731 29975 19737
rect 32125 19771 32183 19777
rect 32125 19737 32137 19771
rect 32171 19768 32183 19771
rect 32171 19740 32260 19768
rect 32171 19737 32183 19740
rect 32125 19731 32183 19737
rect 32232 19712 32260 19740
rect 28592 19672 28764 19700
rect 28813 19703 28871 19709
rect 28592 19660 28598 19672
rect 28813 19669 28825 19703
rect 28859 19700 28871 19703
rect 28902 19700 28908 19712
rect 28859 19672 28908 19700
rect 28859 19669 28871 19672
rect 28813 19663 28871 19669
rect 28902 19660 28908 19672
rect 28960 19660 28966 19712
rect 29730 19700 29736 19712
rect 29691 19672 29736 19700
rect 29730 19660 29736 19672
rect 29788 19660 29794 19712
rect 32214 19660 32220 19712
rect 32272 19660 32278 19712
rect 32509 19700 32537 19808
rect 32600 19768 32628 19876
rect 32674 19864 32680 19876
rect 32732 19864 32738 19916
rect 33686 19904 33692 19916
rect 33244 19876 33692 19904
rect 32858 19836 32864 19848
rect 32819 19808 32864 19836
rect 32858 19796 32864 19808
rect 32916 19796 32922 19848
rect 33009 19839 33067 19845
rect 33009 19805 33021 19839
rect 33055 19836 33067 19839
rect 33244 19836 33272 19876
rect 33686 19864 33692 19876
rect 33744 19864 33750 19916
rect 37921 19907 37979 19913
rect 37921 19904 37933 19907
rect 36924 19876 37933 19904
rect 36924 19848 36952 19876
rect 37921 19873 37933 19876
rect 37967 19873 37979 19907
rect 37921 19867 37979 19873
rect 33055 19808 33272 19836
rect 33326 19839 33384 19845
rect 33055 19805 33067 19808
rect 33009 19799 33067 19805
rect 33326 19805 33338 19839
rect 33372 19836 33384 19839
rect 36906 19836 36912 19848
rect 33372 19808 33456 19836
rect 36867 19808 36912 19836
rect 33372 19805 33384 19808
rect 33326 19799 33384 19805
rect 33137 19771 33195 19777
rect 33137 19768 33149 19771
rect 32600 19740 33149 19768
rect 32876 19712 32904 19740
rect 33137 19737 33149 19740
rect 33183 19737 33195 19771
rect 33137 19731 33195 19737
rect 33226 19728 33232 19780
rect 33284 19768 33290 19780
rect 33284 19740 33329 19768
rect 33284 19728 33290 19740
rect 32674 19700 32680 19712
rect 32509 19672 32680 19700
rect 32674 19660 32680 19672
rect 32732 19660 32738 19712
rect 32858 19660 32864 19712
rect 32916 19660 32922 19712
rect 33042 19660 33048 19712
rect 33100 19700 33106 19712
rect 33428 19700 33456 19808
rect 36906 19796 36912 19808
rect 36964 19796 36970 19848
rect 37093 19839 37151 19845
rect 37093 19805 37105 19839
rect 37139 19805 37151 19839
rect 37734 19836 37740 19848
rect 37695 19808 37740 19836
rect 37093 19799 37151 19805
rect 37108 19768 37136 19799
rect 37734 19796 37740 19808
rect 37792 19796 37798 19848
rect 38013 19839 38071 19845
rect 38013 19805 38025 19839
rect 38059 19836 38071 19839
rect 38286 19836 38292 19848
rect 38059 19808 38292 19836
rect 38059 19805 38071 19808
rect 38013 19799 38071 19805
rect 38028 19768 38056 19799
rect 38286 19796 38292 19808
rect 38344 19796 38350 19848
rect 37108 19740 38056 19768
rect 33100 19672 33456 19700
rect 33100 19660 33106 19672
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 3694 19456 3700 19508
rect 3752 19496 3758 19508
rect 3973 19499 4031 19505
rect 3973 19496 3985 19499
rect 3752 19468 3985 19496
rect 3752 19456 3758 19468
rect 3973 19465 3985 19468
rect 4019 19496 4031 19499
rect 7190 19496 7196 19508
rect 4019 19468 7196 19496
rect 4019 19465 4031 19468
rect 3973 19459 4031 19465
rect 7190 19456 7196 19468
rect 7248 19456 7254 19508
rect 10965 19499 11023 19505
rect 10965 19465 10977 19499
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 2590 19388 2596 19440
rect 2648 19428 2654 19440
rect 2838 19431 2896 19437
rect 2838 19428 2850 19431
rect 2648 19400 2850 19428
rect 2648 19388 2654 19400
rect 2838 19397 2850 19400
rect 2884 19397 2896 19431
rect 2838 19391 2896 19397
rect 4700 19431 4758 19437
rect 4700 19397 4712 19431
rect 4746 19428 4758 19431
rect 4890 19428 4896 19440
rect 4746 19400 4896 19428
rect 4746 19397 4758 19400
rect 4700 19391 4758 19397
rect 4890 19388 4896 19400
rect 4948 19388 4954 19440
rect 1394 19360 1400 19372
rect 1355 19332 1400 19360
rect 1394 19320 1400 19332
rect 1452 19320 1458 19372
rect 2682 19360 2688 19372
rect 2608 19332 2688 19360
rect 1486 19252 1492 19304
rect 1544 19292 1550 19304
rect 2498 19292 2504 19304
rect 1544 19264 2504 19292
rect 1544 19252 1550 19264
rect 2498 19252 2504 19264
rect 2556 19292 2562 19304
rect 2608 19301 2636 19332
rect 2682 19320 2688 19332
rect 2740 19360 2746 19372
rect 4433 19363 4491 19369
rect 4433 19360 4445 19363
rect 2740 19332 4445 19360
rect 2740 19320 2746 19332
rect 4433 19329 4445 19332
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 7098 19320 7104 19372
rect 7156 19360 7162 19372
rect 8202 19360 8208 19372
rect 7156 19332 8208 19360
rect 7156 19320 7162 19332
rect 8202 19320 8208 19332
rect 8260 19360 8266 19372
rect 9490 19360 9496 19372
rect 8260 19332 9496 19360
rect 8260 19320 8266 19332
rect 9490 19320 9496 19332
rect 9548 19360 9554 19372
rect 9858 19369 9864 19372
rect 9585 19363 9643 19369
rect 9585 19360 9597 19363
rect 9548 19332 9597 19360
rect 9548 19320 9554 19332
rect 9585 19329 9597 19332
rect 9631 19329 9643 19363
rect 9585 19323 9643 19329
rect 9852 19323 9864 19369
rect 9916 19360 9922 19372
rect 10980 19360 11008 19459
rect 11422 19456 11428 19508
rect 11480 19496 11486 19508
rect 12066 19496 12072 19508
rect 11480 19468 12072 19496
rect 11480 19456 11486 19468
rect 12066 19456 12072 19468
rect 12124 19456 12130 19508
rect 13906 19456 13912 19508
rect 13964 19496 13970 19508
rect 14001 19499 14059 19505
rect 14001 19496 14013 19499
rect 13964 19468 14013 19496
rect 13964 19456 13970 19468
rect 14001 19465 14013 19468
rect 14047 19465 14059 19499
rect 14001 19459 14059 19465
rect 14458 19456 14464 19508
rect 14516 19496 14522 19508
rect 15562 19496 15568 19508
rect 14516 19468 15568 19496
rect 14516 19456 14522 19468
rect 12802 19360 12808 19372
rect 9916 19332 9952 19360
rect 10980 19332 12808 19360
rect 9858 19320 9864 19323
rect 9916 19320 9922 19332
rect 12802 19320 12808 19332
rect 12860 19360 12866 19372
rect 13357 19363 13415 19369
rect 13357 19360 13369 19363
rect 12860 19332 13369 19360
rect 12860 19320 12866 19332
rect 13357 19329 13369 19332
rect 13403 19329 13415 19363
rect 13357 19323 13415 19329
rect 13722 19320 13728 19372
rect 13780 19360 13786 19372
rect 15194 19360 15200 19372
rect 13780 19332 15056 19360
rect 15155 19332 15200 19360
rect 13780 19320 13786 19332
rect 2593 19295 2651 19301
rect 2593 19292 2605 19295
rect 2556 19264 2605 19292
rect 2556 19252 2562 19264
rect 2593 19261 2605 19264
rect 2639 19261 2651 19295
rect 2593 19255 2651 19261
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19292 13599 19295
rect 13814 19292 13820 19304
rect 13587 19264 13820 19292
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 13814 19252 13820 19264
rect 13872 19252 13878 19304
rect 14182 19292 14188 19304
rect 14144 19264 14188 19292
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14278 19295 14336 19301
rect 14278 19261 14290 19295
rect 14324 19261 14336 19295
rect 14278 19255 14336 19261
rect 14369 19295 14427 19301
rect 14369 19261 14381 19295
rect 14415 19261 14427 19295
rect 14369 19255 14427 19261
rect 14292 19168 14320 19255
rect 14384 19224 14412 19255
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 15028 19301 15056 19332
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 15488 19369 15516 19468
rect 15562 19456 15568 19468
rect 15620 19456 15626 19508
rect 17402 19456 17408 19508
rect 17460 19496 17466 19508
rect 18325 19499 18383 19505
rect 18325 19496 18337 19499
rect 17460 19468 18337 19496
rect 17460 19456 17466 19468
rect 18325 19465 18337 19468
rect 18371 19465 18383 19499
rect 22026 19499 22084 19505
rect 18325 19459 18383 19465
rect 18525 19468 20760 19496
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 15746 19320 15752 19372
rect 15804 19360 15810 19372
rect 18525 19360 18553 19468
rect 20622 19428 20628 19440
rect 18616 19400 20628 19428
rect 18616 19369 18644 19400
rect 20622 19388 20628 19400
rect 20680 19388 20686 19440
rect 15804 19332 18553 19360
rect 18601 19363 18659 19369
rect 15804 19320 15810 19332
rect 18601 19329 18613 19363
rect 18647 19329 18659 19363
rect 20732 19360 20760 19468
rect 22026 19465 22038 19499
rect 22072 19496 22084 19499
rect 22072 19468 22140 19496
rect 22072 19465 22084 19468
rect 22026 19459 22084 19465
rect 20806 19388 20812 19440
rect 20864 19428 20870 19440
rect 21818 19428 21824 19440
rect 20864 19400 21824 19428
rect 20864 19388 20870 19400
rect 21818 19388 21824 19400
rect 21876 19388 21882 19440
rect 22112 19372 22140 19468
rect 22186 19456 22192 19508
rect 22244 19496 22250 19508
rect 22244 19468 22337 19496
rect 22244 19456 22250 19468
rect 23842 19456 23848 19508
rect 23900 19496 23906 19508
rect 24397 19499 24455 19505
rect 24397 19496 24409 19499
rect 23900 19468 24409 19496
rect 23900 19456 23906 19468
rect 24397 19465 24409 19468
rect 24443 19465 24455 19499
rect 26970 19496 26976 19508
rect 26931 19468 26976 19496
rect 24397 19459 24455 19465
rect 26970 19456 26976 19468
rect 27028 19456 27034 19508
rect 27062 19456 27068 19508
rect 27120 19496 27126 19508
rect 27120 19468 33088 19496
rect 27120 19456 27126 19468
rect 22204 19428 22232 19456
rect 28810 19428 28816 19440
rect 22204 19400 27476 19428
rect 21910 19360 21916 19372
rect 20732 19332 21916 19360
rect 18601 19323 18659 19329
rect 21910 19320 21916 19332
rect 21968 19320 21974 19372
rect 22094 19320 22100 19372
rect 22152 19320 22158 19372
rect 24210 19360 24216 19372
rect 24171 19332 24216 19360
rect 24210 19320 24216 19332
rect 24268 19320 24274 19372
rect 27448 19369 27476 19400
rect 28000 19400 28816 19428
rect 28000 19372 28028 19400
rect 28810 19388 28816 19400
rect 28868 19388 28874 19440
rect 29546 19388 29552 19440
rect 29604 19428 29610 19440
rect 32401 19431 32459 19437
rect 29604 19400 32261 19428
rect 29604 19388 29610 19400
rect 27433 19363 27491 19369
rect 27433 19329 27445 19363
rect 27479 19329 27491 19363
rect 27982 19360 27988 19372
rect 27943 19332 27988 19360
rect 27433 19323 27491 19329
rect 27982 19320 27988 19332
rect 28040 19320 28046 19372
rect 28169 19363 28227 19369
rect 28169 19329 28181 19363
rect 28215 19360 28227 19363
rect 28215 19332 28488 19360
rect 28215 19329 28227 19332
rect 28169 19323 28227 19329
rect 15013 19295 15071 19301
rect 14516 19264 14561 19292
rect 14516 19252 14522 19264
rect 15013 19261 15025 19295
rect 15059 19261 15071 19295
rect 15286 19292 15292 19304
rect 15247 19264 15292 19292
rect 15013 19255 15071 19261
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15378 19252 15384 19304
rect 15436 19292 15442 19304
rect 15436 19264 15481 19292
rect 15436 19252 15442 19264
rect 16298 19252 16304 19304
rect 16356 19292 16362 19304
rect 17037 19295 17095 19301
rect 17037 19292 17049 19295
rect 16356 19264 17049 19292
rect 16356 19252 16362 19264
rect 17037 19261 17049 19264
rect 17083 19261 17095 19295
rect 17037 19255 17095 19261
rect 17313 19295 17371 19301
rect 17313 19261 17325 19295
rect 17359 19292 17371 19295
rect 17586 19292 17592 19304
rect 17359 19264 17592 19292
rect 17359 19261 17371 19264
rect 17313 19255 17371 19261
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 18506 19292 18512 19304
rect 18468 19264 18512 19292
rect 18506 19252 18512 19264
rect 18564 19252 18570 19304
rect 18690 19292 18696 19304
rect 18651 19264 18696 19292
rect 18690 19252 18696 19264
rect 18748 19252 18754 19304
rect 18785 19295 18843 19301
rect 18785 19261 18797 19295
rect 18831 19292 18843 19295
rect 18966 19292 18972 19304
rect 18831 19264 18972 19292
rect 18831 19261 18843 19264
rect 18785 19255 18843 19261
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 27154 19292 27160 19304
rect 27115 19264 27160 19292
rect 27154 19252 27160 19264
rect 27212 19252 27218 19304
rect 27249 19295 27307 19301
rect 27249 19261 27261 19295
rect 27295 19261 27307 19295
rect 27249 19255 27307 19261
rect 27341 19295 27399 19301
rect 27341 19261 27353 19295
rect 27387 19292 27399 19295
rect 28460 19292 28488 19332
rect 28534 19320 28540 19372
rect 28592 19360 28598 19372
rect 28629 19363 28687 19369
rect 28629 19360 28641 19363
rect 28592 19332 28641 19360
rect 28592 19320 28598 19332
rect 28629 19329 28641 19332
rect 28675 19329 28687 19363
rect 28902 19360 28908 19372
rect 28863 19332 28908 19360
rect 28629 19323 28687 19329
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 32233 19369 32261 19400
rect 32401 19397 32413 19431
rect 32447 19428 32459 19431
rect 32858 19428 32864 19440
rect 32447 19400 32864 19428
rect 32447 19397 32459 19400
rect 32401 19391 32459 19397
rect 32858 19388 32864 19400
rect 32916 19388 32922 19440
rect 33060 19428 33088 19468
rect 33134 19456 33140 19508
rect 33192 19496 33198 19508
rect 33689 19499 33747 19505
rect 33689 19496 33701 19499
rect 33192 19468 33701 19496
rect 33192 19456 33198 19468
rect 33689 19465 33701 19468
rect 33735 19465 33747 19499
rect 33689 19459 33747 19465
rect 33873 19499 33931 19505
rect 33873 19465 33885 19499
rect 33919 19496 33931 19499
rect 34514 19496 34520 19508
rect 33919 19468 34520 19496
rect 33919 19465 33931 19468
rect 33873 19459 33931 19465
rect 34514 19456 34520 19468
rect 34572 19456 34578 19508
rect 37734 19428 37740 19440
rect 33060 19400 37740 19428
rect 37734 19388 37740 19400
rect 37792 19388 37798 19440
rect 32114 19363 32172 19369
rect 32114 19329 32126 19363
rect 32160 19329 32172 19363
rect 32114 19323 32172 19329
rect 32218 19363 32276 19369
rect 32218 19329 32230 19363
rect 32264 19329 32276 19363
rect 32218 19323 32276 19329
rect 28920 19292 28948 19320
rect 27387 19264 28212 19292
rect 28460 19264 28948 19292
rect 27387 19261 27399 19264
rect 27341 19255 27399 19261
rect 15396 19224 15424 19252
rect 14384 19196 15424 19224
rect 20622 19184 20628 19236
rect 20680 19224 20686 19236
rect 24210 19224 24216 19236
rect 20680 19196 24216 19224
rect 20680 19184 20686 19196
rect 24210 19184 24216 19196
rect 24268 19184 24274 19236
rect 27264 19224 27292 19255
rect 28077 19227 28135 19233
rect 28077 19224 28089 19227
rect 27264 19196 28089 19224
rect 28077 19193 28089 19196
rect 28123 19193 28135 19227
rect 28184 19224 28212 19264
rect 31846 19252 31852 19304
rect 31904 19292 31910 19304
rect 32140 19292 32168 19323
rect 32490 19320 32496 19372
rect 32548 19360 32554 19372
rect 32674 19369 32680 19372
rect 32631 19363 32680 19369
rect 32548 19332 32593 19360
rect 32548 19320 32554 19332
rect 32631 19329 32643 19363
rect 32677 19329 32680 19363
rect 32631 19323 32680 19329
rect 32674 19320 32680 19323
rect 32732 19360 32738 19372
rect 33042 19360 33048 19372
rect 32732 19332 33048 19360
rect 32732 19320 32738 19332
rect 33042 19320 33048 19332
rect 33100 19320 33106 19372
rect 33321 19363 33379 19369
rect 33321 19329 33333 19363
rect 33367 19360 33379 19363
rect 34054 19360 34060 19372
rect 33367 19332 34060 19360
rect 33367 19329 33379 19332
rect 33321 19323 33379 19329
rect 34054 19320 34060 19332
rect 34112 19360 34118 19372
rect 34422 19360 34428 19372
rect 34112 19332 34428 19360
rect 34112 19320 34118 19332
rect 34422 19320 34428 19332
rect 34480 19320 34486 19372
rect 44082 19360 44088 19372
rect 44043 19332 44088 19360
rect 44082 19320 44088 19332
rect 44140 19320 44146 19372
rect 32950 19292 32956 19304
rect 31904 19264 32956 19292
rect 31904 19252 31910 19264
rect 32600 19236 32628 19264
rect 32950 19252 32956 19264
rect 33008 19252 33014 19304
rect 35434 19252 35440 19304
rect 35492 19292 35498 19304
rect 37829 19295 37887 19301
rect 37829 19292 37841 19295
rect 35492 19264 37841 19292
rect 35492 19252 35498 19264
rect 37829 19261 37841 19264
rect 37875 19292 37887 19295
rect 38010 19292 38016 19304
rect 37875 19264 38016 19292
rect 37875 19261 37887 19264
rect 37829 19255 37887 19261
rect 38010 19252 38016 19264
rect 38068 19252 38074 19304
rect 38105 19295 38163 19301
rect 38105 19261 38117 19295
rect 38151 19292 38163 19295
rect 38286 19292 38292 19304
rect 38151 19264 38292 19292
rect 38151 19261 38163 19264
rect 38105 19255 38163 19261
rect 38286 19252 38292 19264
rect 38344 19252 38350 19304
rect 30374 19224 30380 19236
rect 28184 19196 30380 19224
rect 28077 19187 28135 19193
rect 30374 19184 30380 19196
rect 30432 19184 30438 19236
rect 32582 19184 32588 19236
rect 32640 19184 32646 19236
rect 32766 19224 32772 19236
rect 32727 19196 32772 19224
rect 32766 19184 32772 19196
rect 32824 19184 32830 19236
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 5813 19159 5871 19165
rect 5813 19125 5825 19159
rect 5859 19156 5871 19159
rect 5994 19156 6000 19168
rect 5859 19128 6000 19156
rect 5859 19125 5871 19128
rect 5813 19119 5871 19125
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 14274 19116 14280 19168
rect 14332 19116 14338 19168
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 19058 19156 19064 19168
rect 16448 19128 19064 19156
rect 16448 19116 16454 19128
rect 19058 19116 19064 19128
rect 19116 19116 19122 19168
rect 21634 19116 21640 19168
rect 21692 19156 21698 19168
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 21692 19128 22017 19156
rect 21692 19116 21698 19128
rect 22005 19125 22017 19128
rect 22051 19125 22063 19159
rect 22005 19119 22063 19125
rect 26878 19116 26884 19168
rect 26936 19156 26942 19168
rect 32674 19156 32680 19168
rect 26936 19128 32680 19156
rect 26936 19116 26942 19128
rect 32674 19116 32680 19128
rect 32732 19116 32738 19168
rect 33686 19156 33692 19168
rect 33647 19128 33692 19156
rect 33686 19116 33692 19128
rect 33744 19116 33750 19168
rect 43898 19156 43904 19168
rect 43859 19128 43904 19156
rect 43898 19116 43904 19128
rect 43956 19116 43962 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 1394 18912 1400 18964
rect 1452 18952 1458 18964
rect 2682 18952 2688 18964
rect 1452 18924 2688 18952
rect 1452 18912 1458 18924
rect 2682 18912 2688 18924
rect 2740 18952 2746 18964
rect 2961 18955 3019 18961
rect 2961 18952 2973 18955
rect 2740 18924 2973 18952
rect 2740 18912 2746 18924
rect 2961 18921 2973 18924
rect 3007 18921 3019 18955
rect 2961 18915 3019 18921
rect 4893 18955 4951 18961
rect 4893 18921 4905 18955
rect 4939 18952 4951 18955
rect 5074 18952 5080 18964
rect 4939 18924 5080 18952
rect 4939 18921 4951 18924
rect 4893 18915 4951 18921
rect 5074 18912 5080 18924
rect 5132 18912 5138 18964
rect 13078 18952 13084 18964
rect 7576 18924 13084 18952
rect 7576 18884 7604 18924
rect 13078 18912 13084 18924
rect 13136 18912 13142 18964
rect 13170 18912 13176 18964
rect 13228 18952 13234 18964
rect 15470 18952 15476 18964
rect 13228 18924 15476 18952
rect 13228 18912 13234 18924
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 15654 18952 15660 18964
rect 15615 18924 15660 18952
rect 15654 18912 15660 18924
rect 15712 18952 15718 18964
rect 15930 18952 15936 18964
rect 15712 18924 15936 18952
rect 15712 18912 15718 18924
rect 15930 18912 15936 18924
rect 15988 18912 15994 18964
rect 16114 18912 16120 18964
rect 16172 18952 16178 18964
rect 20990 18952 20996 18964
rect 16172 18924 20996 18952
rect 16172 18912 16178 18924
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 27154 18912 27160 18964
rect 27212 18952 27218 18964
rect 27525 18955 27583 18961
rect 27525 18952 27537 18955
rect 27212 18924 27537 18952
rect 27212 18912 27218 18924
rect 27525 18921 27537 18924
rect 27571 18921 27583 18955
rect 27525 18915 27583 18921
rect 32674 18912 32680 18964
rect 32732 18952 32738 18964
rect 33229 18955 33287 18961
rect 33229 18952 33241 18955
rect 32732 18924 33241 18952
rect 32732 18912 32738 18924
rect 33229 18921 33241 18924
rect 33275 18921 33287 18955
rect 33229 18915 33287 18921
rect 37274 18912 37280 18964
rect 37332 18952 37338 18964
rect 41233 18955 41291 18961
rect 41233 18952 41245 18955
rect 37332 18924 41245 18952
rect 37332 18912 37338 18924
rect 41233 18921 41245 18924
rect 41279 18921 41291 18955
rect 41233 18915 41291 18921
rect 9858 18884 9864 18896
rect 2608 18856 7604 18884
rect 9819 18856 9864 18884
rect 1486 18776 1492 18828
rect 1544 18816 1550 18828
rect 1581 18819 1639 18825
rect 1581 18816 1593 18819
rect 1544 18788 1593 18816
rect 1544 18776 1550 18788
rect 1581 18785 1593 18788
rect 1627 18785 1639 18819
rect 1581 18779 1639 18785
rect 1670 18708 1676 18760
rect 1728 18748 1734 18760
rect 2608 18748 2636 18856
rect 9858 18844 9864 18856
rect 9916 18844 9922 18896
rect 15838 18844 15844 18896
rect 15896 18884 15902 18896
rect 27706 18884 27712 18896
rect 15896 18856 15941 18884
rect 17926 18856 27712 18884
rect 15896 18844 15902 18856
rect 5537 18819 5595 18825
rect 5537 18785 5549 18819
rect 5583 18816 5595 18819
rect 6730 18816 6736 18828
rect 5583 18788 6736 18816
rect 5583 18785 5595 18788
rect 5537 18779 5595 18785
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 14277 18819 14335 18825
rect 14277 18785 14289 18819
rect 14323 18816 14335 18819
rect 14918 18816 14924 18828
rect 14323 18788 14924 18816
rect 14323 18785 14335 18788
rect 14277 18779 14335 18785
rect 14918 18776 14924 18788
rect 14976 18776 14982 18828
rect 15286 18776 15292 18828
rect 15344 18816 15350 18828
rect 17926 18816 17954 18856
rect 27706 18844 27712 18856
rect 27764 18844 27770 18896
rect 27798 18844 27804 18896
rect 27856 18884 27862 18896
rect 33686 18884 33692 18896
rect 27856 18856 33692 18884
rect 27856 18844 27862 18856
rect 33686 18844 33692 18856
rect 33744 18844 33750 18896
rect 37826 18844 37832 18896
rect 37884 18884 37890 18896
rect 38562 18884 38568 18896
rect 37884 18856 38568 18884
rect 37884 18844 37890 18856
rect 38562 18844 38568 18856
rect 38620 18884 38626 18896
rect 38620 18856 39896 18884
rect 38620 18844 38626 18856
rect 15344 18788 17954 18816
rect 18417 18819 18475 18825
rect 15344 18776 15350 18788
rect 18417 18785 18429 18819
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 3970 18748 3976 18760
rect 1728 18720 2636 18748
rect 3931 18720 3976 18748
rect 1728 18708 1734 18720
rect 3970 18708 3976 18720
rect 4028 18708 4034 18760
rect 7098 18748 7104 18760
rect 7059 18720 7104 18748
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 10045 18751 10103 18757
rect 10045 18748 10057 18751
rect 9732 18720 10057 18748
rect 9732 18708 9738 18720
rect 10045 18717 10057 18720
rect 10091 18717 10103 18751
rect 11422 18748 11428 18760
rect 11383 18720 11428 18748
rect 10045 18711 10103 18717
rect 11422 18708 11428 18720
rect 11480 18748 11486 18760
rect 12158 18748 12164 18760
rect 11480 18720 12164 18748
rect 11480 18708 11486 18720
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18748 14611 18751
rect 16114 18748 16120 18760
rect 14599 18720 16120 18748
rect 14599 18717 14611 18720
rect 14553 18711 14611 18717
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 16850 18708 16856 18760
rect 16908 18748 16914 18760
rect 17129 18751 17187 18757
rect 16908 18720 16953 18748
rect 16908 18708 16914 18720
rect 17129 18717 17141 18751
rect 17175 18748 17187 18751
rect 18138 18748 18144 18760
rect 17175 18720 18144 18748
rect 17175 18717 17187 18720
rect 17129 18711 17187 18717
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 18322 18748 18328 18760
rect 18283 18720 18328 18748
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 1848 18683 1906 18689
rect 1848 18649 1860 18683
rect 1894 18680 1906 18683
rect 2314 18680 2320 18692
rect 1894 18652 2320 18680
rect 1894 18649 1906 18652
rect 1848 18643 1906 18649
rect 2314 18640 2320 18652
rect 2372 18640 2378 18692
rect 5353 18683 5411 18689
rect 5353 18680 5365 18683
rect 3804 18652 5365 18680
rect 3804 18621 3832 18652
rect 5353 18649 5365 18652
rect 5399 18649 5411 18683
rect 5353 18643 5411 18649
rect 11692 18683 11750 18689
rect 11692 18649 11704 18683
rect 11738 18680 11750 18683
rect 12618 18680 12624 18692
rect 11738 18652 12624 18680
rect 11738 18649 11750 18652
rect 11692 18643 11750 18649
rect 12618 18640 12624 18652
rect 12676 18640 12682 18692
rect 14461 18683 14519 18689
rect 14461 18680 14473 18683
rect 12728 18652 14473 18680
rect 3789 18615 3847 18621
rect 3789 18581 3801 18615
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 5261 18615 5319 18621
rect 5261 18581 5273 18615
rect 5307 18612 5319 18615
rect 5994 18612 6000 18624
rect 5307 18584 6000 18612
rect 5307 18581 5319 18584
rect 5261 18575 5319 18581
rect 5994 18572 6000 18584
rect 6052 18572 6058 18624
rect 6914 18612 6920 18624
rect 6875 18584 6920 18612
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7558 18572 7564 18624
rect 7616 18612 7622 18624
rect 12728 18612 12756 18652
rect 14461 18649 14473 18652
rect 14507 18649 14519 18683
rect 15010 18680 15016 18692
rect 14971 18652 15016 18680
rect 14461 18643 14519 18649
rect 15010 18640 15016 18652
rect 15068 18640 15074 18692
rect 15286 18640 15292 18692
rect 15344 18680 15350 18692
rect 15473 18683 15531 18689
rect 15473 18680 15485 18683
rect 15344 18652 15485 18680
rect 15344 18640 15350 18652
rect 15473 18649 15485 18652
rect 15519 18649 15531 18683
rect 15838 18680 15844 18692
rect 15473 18643 15531 18649
rect 15580 18652 15844 18680
rect 7616 18584 12756 18612
rect 12805 18615 12863 18621
rect 7616 18572 7622 18584
rect 12805 18581 12817 18615
rect 12851 18612 12863 18615
rect 12986 18612 12992 18624
rect 12851 18584 12992 18612
rect 12851 18581 12863 18584
rect 12805 18575 12863 18581
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 15580 18612 15608 18652
rect 15838 18640 15844 18652
rect 15896 18640 15902 18692
rect 16298 18680 16304 18692
rect 15948 18652 16304 18680
rect 13320 18584 15608 18612
rect 15683 18615 15741 18621
rect 13320 18572 13326 18584
rect 15683 18581 15695 18615
rect 15729 18612 15741 18615
rect 15948 18612 15976 18652
rect 16298 18640 16304 18652
rect 16356 18640 16362 18692
rect 16390 18640 16396 18692
rect 16448 18680 16454 18692
rect 17494 18680 17500 18692
rect 16448 18652 17500 18680
rect 16448 18640 16454 18652
rect 17494 18640 17500 18652
rect 17552 18640 17558 18692
rect 15729 18584 15976 18612
rect 15729 18581 15741 18584
rect 15683 18575 15741 18581
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 18141 18615 18199 18621
rect 18141 18612 18153 18615
rect 16080 18584 18153 18612
rect 16080 18572 16086 18584
rect 18141 18581 18153 18584
rect 18187 18581 18199 18615
rect 18432 18612 18460 18779
rect 18506 18776 18512 18828
rect 18564 18816 18570 18828
rect 18564 18788 18609 18816
rect 18564 18776 18570 18788
rect 18966 18776 18972 18828
rect 19024 18776 19030 18828
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 26878 18816 26884 18828
rect 19116 18788 26884 18816
rect 19116 18776 19122 18788
rect 26878 18776 26884 18788
rect 26936 18776 26942 18828
rect 28810 18776 28816 18828
rect 28868 18816 28874 18828
rect 29825 18819 29883 18825
rect 29825 18816 29837 18819
rect 28868 18788 29837 18816
rect 28868 18776 28874 18788
rect 29825 18785 29837 18788
rect 29871 18785 29883 18819
rect 35434 18816 35440 18828
rect 29825 18779 29883 18785
rect 32968 18788 35440 18816
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18748 18659 18751
rect 18984 18748 19012 18776
rect 18647 18720 19012 18748
rect 18647 18717 18659 18720
rect 18601 18711 18659 18717
rect 18506 18640 18512 18692
rect 18564 18680 18570 18692
rect 18616 18680 18644 18711
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 27246 18748 27252 18760
rect 20036 18720 27252 18748
rect 20036 18708 20042 18720
rect 27246 18708 27252 18720
rect 27304 18708 27310 18760
rect 27341 18751 27399 18757
rect 27341 18717 27353 18751
rect 27387 18748 27399 18751
rect 28902 18748 28908 18760
rect 27387 18720 28908 18748
rect 27387 18717 27399 18720
rect 27341 18711 27399 18717
rect 28902 18708 28908 18720
rect 28960 18708 28966 18760
rect 28994 18708 29000 18760
rect 29052 18748 29058 18760
rect 29549 18751 29607 18757
rect 29549 18748 29561 18751
rect 29052 18720 29561 18748
rect 29052 18708 29058 18720
rect 29549 18717 29561 18720
rect 29595 18748 29607 18751
rect 29638 18748 29644 18760
rect 29595 18720 29644 18748
rect 29595 18717 29607 18720
rect 29549 18711 29607 18717
rect 29638 18708 29644 18720
rect 29696 18708 29702 18760
rect 32582 18748 32588 18760
rect 32543 18720 32588 18748
rect 32582 18708 32588 18720
rect 32640 18708 32646 18760
rect 32733 18751 32791 18757
rect 32733 18717 32745 18751
rect 32779 18748 32791 18751
rect 32968 18748 32996 18788
rect 35434 18776 35440 18788
rect 35492 18776 35498 18828
rect 39868 18825 39896 18856
rect 39853 18819 39911 18825
rect 38120 18788 39160 18816
rect 32779 18720 32996 18748
rect 32779 18717 32791 18720
rect 32733 18711 32791 18717
rect 33042 18708 33048 18760
rect 33100 18757 33106 18760
rect 33100 18748 33108 18757
rect 36630 18748 36636 18760
rect 33100 18720 33145 18748
rect 36591 18720 36636 18748
rect 33100 18711 33108 18720
rect 33100 18708 33106 18711
rect 36630 18708 36636 18720
rect 36688 18708 36694 18760
rect 36906 18748 36912 18760
rect 36867 18720 36912 18748
rect 36906 18708 36912 18720
rect 36964 18708 36970 18760
rect 37182 18708 37188 18760
rect 37240 18748 37246 18760
rect 38120 18757 38148 18788
rect 39132 18757 39160 18788
rect 39853 18785 39865 18819
rect 39899 18785 39911 18819
rect 39853 18779 39911 18785
rect 38105 18751 38163 18757
rect 38105 18748 38117 18751
rect 37240 18720 38117 18748
rect 37240 18708 37246 18720
rect 38105 18717 38117 18720
rect 38151 18717 38163 18751
rect 38105 18711 38163 18717
rect 38381 18751 38439 18757
rect 38381 18717 38393 18751
rect 38427 18748 38439 18751
rect 38841 18751 38899 18757
rect 38841 18748 38853 18751
rect 38427 18720 38853 18748
rect 38427 18717 38439 18720
rect 38381 18711 38439 18717
rect 38841 18717 38853 18720
rect 38887 18717 38899 18751
rect 38841 18711 38899 18717
rect 39117 18751 39175 18757
rect 39117 18717 39129 18751
rect 39163 18717 39175 18751
rect 43070 18748 43076 18760
rect 43031 18720 43076 18748
rect 39117 18711 39175 18717
rect 18564 18652 18644 18680
rect 18564 18640 18570 18652
rect 18966 18640 18972 18692
rect 19024 18680 19030 18692
rect 23658 18680 23664 18692
rect 19024 18652 23664 18680
rect 19024 18640 19030 18652
rect 23658 18640 23664 18652
rect 23716 18640 23722 18692
rect 27154 18680 27160 18692
rect 27115 18652 27160 18680
rect 27154 18640 27160 18652
rect 27212 18680 27218 18692
rect 27982 18680 27988 18692
rect 27212 18652 27988 18680
rect 27212 18640 27218 18652
rect 27982 18640 27988 18652
rect 28040 18640 28046 18692
rect 32858 18680 32864 18692
rect 32819 18652 32864 18680
rect 32858 18640 32864 18652
rect 32916 18640 32922 18692
rect 32953 18683 33011 18689
rect 32953 18649 32965 18683
rect 32999 18680 33011 18683
rect 36924 18680 36952 18708
rect 38396 18680 38424 18711
rect 43070 18708 43076 18720
rect 43128 18708 43134 18760
rect 43340 18751 43398 18757
rect 43340 18717 43352 18751
rect 43386 18748 43398 18751
rect 43898 18748 43904 18760
rect 43386 18720 43904 18748
rect 43386 18717 43398 18720
rect 43340 18711 43398 18717
rect 43898 18708 43904 18720
rect 43956 18708 43962 18760
rect 47486 18748 47492 18760
rect 47447 18720 47492 18748
rect 47486 18708 47492 18720
rect 47544 18708 47550 18760
rect 39025 18683 39083 18689
rect 39025 18680 39037 18683
rect 32999 18652 33088 18680
rect 36924 18652 38424 18680
rect 38488 18652 39037 18680
rect 32999 18649 33011 18652
rect 32953 18643 33011 18649
rect 33060 18624 33088 18652
rect 30190 18612 30196 18624
rect 18432 18584 30196 18612
rect 18141 18575 18199 18581
rect 30190 18572 30196 18584
rect 30248 18572 30254 18624
rect 33042 18572 33048 18624
rect 33100 18572 33106 18624
rect 37826 18572 37832 18624
rect 37884 18612 37890 18624
rect 37921 18615 37979 18621
rect 37921 18612 37933 18615
rect 37884 18584 37933 18612
rect 37884 18572 37890 18584
rect 37921 18581 37933 18584
rect 37967 18581 37979 18615
rect 38286 18612 38292 18624
rect 38247 18584 38292 18612
rect 37921 18575 37979 18581
rect 38286 18572 38292 18584
rect 38344 18612 38350 18624
rect 38488 18612 38516 18652
rect 39025 18649 39037 18652
rect 39071 18649 39083 18683
rect 39025 18643 39083 18649
rect 39206 18640 39212 18692
rect 39264 18680 39270 18692
rect 40098 18683 40156 18689
rect 40098 18680 40110 18683
rect 39264 18652 40110 18680
rect 39264 18640 39270 18652
rect 40098 18649 40110 18652
rect 40144 18649 40156 18683
rect 40098 18643 40156 18649
rect 38930 18612 38936 18624
rect 38344 18584 38516 18612
rect 38891 18584 38936 18612
rect 38344 18572 38350 18584
rect 38930 18572 38936 18584
rect 38988 18572 38994 18624
rect 44358 18572 44364 18624
rect 44416 18612 44422 18624
rect 44453 18615 44511 18621
rect 44453 18612 44465 18615
rect 44416 18584 44465 18612
rect 44416 18572 44422 18584
rect 44453 18581 44465 18584
rect 44499 18581 44511 18615
rect 47302 18612 47308 18624
rect 47263 18584 47308 18612
rect 44453 18575 44511 18581
rect 47302 18572 47308 18584
rect 47360 18572 47366 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 1670 18408 1676 18420
rect 1627 18380 1676 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 1670 18368 1676 18380
rect 1728 18368 1734 18420
rect 2314 18408 2320 18420
rect 2275 18380 2320 18408
rect 2314 18368 2320 18380
rect 2372 18368 2378 18420
rect 2682 18408 2688 18420
rect 2643 18380 2688 18408
rect 2682 18368 2688 18380
rect 2740 18368 2746 18420
rect 7558 18408 7564 18420
rect 6840 18380 7564 18408
rect 1946 18300 1952 18352
rect 2004 18340 2010 18352
rect 6840 18340 6868 18380
rect 7558 18368 7564 18380
rect 7616 18368 7622 18420
rect 12618 18408 12624 18420
rect 12579 18380 12624 18408
rect 12618 18368 12624 18380
rect 12676 18368 12682 18420
rect 14185 18411 14243 18417
rect 14185 18377 14197 18411
rect 14231 18408 14243 18411
rect 15194 18408 15200 18420
rect 14231 18380 15200 18408
rect 14231 18377 14243 18380
rect 14185 18371 14243 18377
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 15286 18368 15292 18420
rect 15344 18368 15350 18420
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 17221 18411 17279 18417
rect 17221 18408 17233 18411
rect 15528 18380 17233 18408
rect 15528 18368 15534 18380
rect 17221 18377 17233 18380
rect 17267 18377 17279 18411
rect 18230 18408 18236 18420
rect 17221 18371 17279 18377
rect 17328 18380 18236 18408
rect 2004 18312 6868 18340
rect 2004 18300 2010 18312
rect 6914 18300 6920 18352
rect 6972 18340 6978 18352
rect 7438 18343 7496 18349
rect 7438 18340 7450 18343
rect 6972 18312 7450 18340
rect 6972 18300 6978 18312
rect 7438 18309 7450 18312
rect 7484 18309 7496 18343
rect 12986 18340 12992 18352
rect 12899 18312 12992 18340
rect 7438 18303 7496 18309
rect 12986 18300 12992 18312
rect 13044 18340 13050 18352
rect 15304 18340 15332 18368
rect 17328 18340 17356 18380
rect 18230 18368 18236 18380
rect 18288 18368 18294 18420
rect 18414 18368 18420 18420
rect 18472 18408 18478 18420
rect 19245 18411 19303 18417
rect 19245 18408 19257 18411
rect 18472 18380 19257 18408
rect 18472 18368 18478 18380
rect 19245 18377 19257 18380
rect 19291 18377 19303 18411
rect 19245 18371 19303 18377
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 20990 18408 20996 18420
rect 19392 18380 20484 18408
rect 20951 18380 20996 18408
rect 19392 18368 19398 18380
rect 19978 18340 19984 18352
rect 13044 18312 14596 18340
rect 15304 18312 17356 18340
rect 17512 18312 19984 18340
rect 13044 18300 13050 18312
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 2590 18272 2596 18284
rect 2547 18244 2596 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 2590 18232 2596 18244
rect 2648 18232 2654 18284
rect 2774 18232 2780 18284
rect 2832 18272 2838 18284
rect 3418 18272 3424 18284
rect 2832 18244 2877 18272
rect 3379 18244 3424 18272
rect 2832 18232 2838 18244
rect 3418 18232 3424 18244
rect 3476 18232 3482 18284
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 6549 18275 6607 18281
rect 6549 18272 6561 18275
rect 6512 18244 6561 18272
rect 6512 18232 6518 18244
rect 6549 18241 6561 18244
rect 6595 18241 6607 18275
rect 8202 18272 8208 18284
rect 6549 18235 6607 18241
rect 7208 18244 8208 18272
rect 6914 18164 6920 18216
rect 6972 18204 6978 18216
rect 7208 18213 7236 18244
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 12805 18275 12863 18281
rect 12805 18241 12817 18275
rect 12851 18272 12863 18275
rect 12851 18244 13032 18272
rect 12851 18241 12863 18244
rect 12805 18235 12863 18241
rect 7193 18207 7251 18213
rect 7193 18204 7205 18207
rect 6972 18176 7205 18204
rect 6972 18164 6978 18176
rect 7193 18173 7205 18176
rect 7239 18173 7251 18207
rect 7193 18167 7251 18173
rect 6730 18136 6736 18148
rect 6691 18108 6736 18136
rect 6730 18096 6736 18108
rect 6788 18096 6794 18148
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18068 3295 18071
rect 6546 18068 6552 18080
rect 3283 18040 6552 18068
rect 3283 18037 3295 18040
rect 3237 18031 3295 18037
rect 6546 18028 6552 18040
rect 6604 18028 6610 18080
rect 6822 18028 6828 18080
rect 6880 18068 6886 18080
rect 8573 18071 8631 18077
rect 8573 18068 8585 18071
rect 6880 18040 8585 18068
rect 6880 18028 6886 18040
rect 8573 18037 8585 18040
rect 8619 18037 8631 18071
rect 13004 18068 13032 18244
rect 13078 18232 13084 18284
rect 13136 18272 13142 18284
rect 13538 18272 13544 18284
rect 13136 18244 13544 18272
rect 13136 18232 13142 18244
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14568 18281 14596 18312
rect 14461 18275 14519 18281
rect 14461 18272 14473 18275
rect 13872 18244 14473 18272
rect 13872 18232 13878 18244
rect 14461 18241 14473 18244
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 14553 18275 14611 18281
rect 14553 18241 14565 18275
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 14826 18232 14832 18284
rect 14884 18272 14890 18284
rect 15289 18275 15347 18281
rect 15289 18272 15301 18275
rect 14884 18244 15301 18272
rect 14884 18232 14890 18244
rect 15289 18241 15301 18244
rect 15335 18272 15347 18275
rect 16850 18272 16856 18284
rect 15335 18244 16856 18272
rect 15335 18241 15347 18244
rect 15289 18235 15347 18241
rect 16850 18232 16856 18244
rect 16908 18232 16914 18284
rect 17512 18281 17540 18312
rect 19978 18300 19984 18312
rect 20036 18300 20042 18352
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 18196 18244 18429 18272
rect 18196 18232 18202 18244
rect 18417 18241 18429 18244
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 18607 18272 18736 18278
rect 19334 18272 19340 18284
rect 18607 18250 19340 18272
rect 14369 18207 14427 18213
rect 14369 18173 14381 18207
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 14645 18207 14703 18213
rect 14645 18173 14657 18207
rect 14691 18204 14703 18207
rect 15654 18204 15660 18216
rect 14691 18176 15660 18204
rect 14691 18173 14703 18176
rect 14645 18167 14703 18173
rect 14384 18136 14412 18167
rect 15654 18164 15660 18176
rect 15712 18204 15718 18216
rect 16022 18204 16028 18216
rect 15712 18176 16028 18204
rect 15712 18164 15718 18176
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 17405 18207 17463 18213
rect 17405 18173 17417 18207
rect 17451 18173 17463 18207
rect 17586 18204 17592 18216
rect 17547 18176 17592 18204
rect 17405 18167 17463 18173
rect 15473 18139 15531 18145
rect 15473 18136 15485 18139
rect 14384 18108 15485 18136
rect 15473 18105 15485 18108
rect 15519 18136 15531 18139
rect 16574 18136 16580 18148
rect 15519 18108 16580 18136
rect 15519 18105 15531 18108
rect 15473 18099 15531 18105
rect 16574 18096 16580 18108
rect 16632 18096 16638 18148
rect 17420 18136 17448 18167
rect 17586 18164 17592 18176
rect 17644 18164 17650 18216
rect 17678 18164 17684 18216
rect 17736 18204 17742 18216
rect 18506 18204 18512 18216
rect 17736 18176 18368 18204
rect 18467 18176 18512 18204
rect 17736 18164 17742 18176
rect 18233 18139 18291 18145
rect 18233 18136 18245 18139
rect 17420 18108 18245 18136
rect 18233 18105 18245 18108
rect 18279 18105 18291 18139
rect 18340 18136 18368 18176
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 18607 18213 18635 18250
rect 18708 18244 19340 18250
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18241 19579 18275
rect 20456 18272 20484 18380
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 33870 18408 33876 18420
rect 21928 18380 33876 18408
rect 20806 18340 20812 18352
rect 20767 18312 20812 18340
rect 20806 18300 20812 18312
rect 20864 18300 20870 18352
rect 21928 18340 21956 18380
rect 33870 18368 33876 18380
rect 33928 18368 33934 18420
rect 34790 18408 34796 18420
rect 33980 18380 34796 18408
rect 20916 18312 21956 18340
rect 20916 18272 20944 18312
rect 22186 18300 22192 18352
rect 22244 18340 22250 18352
rect 27433 18343 27491 18349
rect 27433 18340 27445 18343
rect 22244 18312 22289 18340
rect 26988 18312 27445 18340
rect 22244 18300 22250 18312
rect 20456 18244 20944 18272
rect 21269 18275 21327 18281
rect 19521 18235 19579 18241
rect 21269 18241 21281 18275
rect 21315 18272 21327 18275
rect 21910 18272 21916 18284
rect 21315 18244 21916 18272
rect 21315 18241 21327 18244
rect 21269 18235 21327 18241
rect 18601 18207 18659 18213
rect 18601 18173 18613 18207
rect 18647 18173 18659 18207
rect 18601 18167 18659 18173
rect 18693 18207 18751 18213
rect 18693 18173 18705 18207
rect 18739 18173 18751 18207
rect 18693 18167 18751 18173
rect 18414 18136 18420 18148
rect 18340 18108 18420 18136
rect 18233 18099 18291 18105
rect 18414 18096 18420 18108
rect 18472 18096 18478 18148
rect 18708 18136 18736 18167
rect 18874 18164 18880 18216
rect 18932 18204 18938 18216
rect 19429 18207 19487 18213
rect 19429 18204 19441 18207
rect 18932 18176 19441 18204
rect 18932 18164 18938 18176
rect 19429 18173 19441 18176
rect 19475 18173 19487 18207
rect 19429 18167 19487 18173
rect 18616 18108 18736 18136
rect 18616 18080 18644 18108
rect 19058 18096 19064 18148
rect 19116 18136 19122 18148
rect 19536 18136 19564 18235
rect 21910 18232 21916 18244
rect 21968 18272 21974 18284
rect 22024 18278 22082 18281
rect 22020 18275 22082 18278
rect 22020 18272 22036 18275
rect 21968 18244 22036 18272
rect 21968 18232 21974 18244
rect 22024 18241 22036 18244
rect 22070 18241 22082 18275
rect 22024 18235 22082 18241
rect 22278 18275 22336 18281
rect 22278 18241 22290 18275
rect 22324 18272 22336 18275
rect 22370 18272 22376 18284
rect 22324 18244 22376 18272
rect 22324 18241 22336 18244
rect 22278 18235 22336 18241
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 23468 18275 23526 18281
rect 23468 18241 23480 18275
rect 23514 18272 23526 18275
rect 24394 18272 24400 18284
rect 23514 18244 24400 18272
rect 23514 18241 23526 18244
rect 23468 18235 23526 18241
rect 24394 18232 24400 18244
rect 24452 18232 24458 18284
rect 25314 18232 25320 18284
rect 25372 18272 25378 18284
rect 26988 18272 27016 18312
rect 27433 18309 27445 18312
rect 27479 18340 27491 18343
rect 27798 18340 27804 18352
rect 27479 18312 27804 18340
rect 27479 18309 27491 18312
rect 27433 18303 27491 18309
rect 27798 18300 27804 18312
rect 27856 18300 27862 18352
rect 29178 18300 29184 18352
rect 29236 18340 29242 18352
rect 29825 18343 29883 18349
rect 29825 18340 29837 18343
rect 29236 18312 29837 18340
rect 29236 18300 29242 18312
rect 29825 18309 29837 18312
rect 29871 18309 29883 18343
rect 32950 18340 32956 18352
rect 29825 18303 29883 18309
rect 31726 18312 32956 18340
rect 25372 18244 27016 18272
rect 27065 18275 27123 18281
rect 25372 18232 25378 18244
rect 27065 18241 27077 18275
rect 27111 18272 27123 18275
rect 27154 18272 27160 18284
rect 27111 18244 27160 18272
rect 27111 18241 27123 18244
rect 27065 18235 27123 18241
rect 27154 18232 27160 18244
rect 27212 18232 27218 18284
rect 29454 18272 29460 18284
rect 29415 18244 29460 18272
rect 29454 18232 29460 18244
rect 29512 18232 29518 18284
rect 29638 18281 29644 18284
rect 29605 18275 29644 18281
rect 29605 18241 29617 18275
rect 29605 18235 29644 18241
rect 29638 18232 29644 18235
rect 29696 18232 29702 18284
rect 29730 18232 29736 18284
rect 29788 18272 29794 18284
rect 30006 18281 30012 18284
rect 29963 18275 30012 18281
rect 29788 18244 29833 18272
rect 29788 18232 29794 18244
rect 29963 18241 29975 18275
rect 30009 18241 30012 18275
rect 29963 18235 30012 18241
rect 30006 18232 30012 18235
rect 30064 18232 30070 18284
rect 31021 18275 31079 18281
rect 31021 18241 31033 18275
rect 31067 18272 31079 18275
rect 31726 18272 31754 18312
rect 32950 18300 32956 18312
rect 33008 18300 33014 18352
rect 33980 18340 34008 18380
rect 34790 18368 34796 18380
rect 34848 18368 34854 18420
rect 35434 18408 35440 18420
rect 35395 18380 35440 18408
rect 35434 18368 35440 18380
rect 35492 18368 35498 18420
rect 35529 18411 35587 18417
rect 35529 18377 35541 18411
rect 35575 18408 35587 18411
rect 35575 18380 36768 18408
rect 35575 18377 35587 18380
rect 35529 18371 35587 18377
rect 33888 18312 34008 18340
rect 31067 18244 31754 18272
rect 32677 18275 32735 18281
rect 31067 18241 31079 18244
rect 31021 18235 31079 18241
rect 32677 18241 32689 18275
rect 32723 18272 32735 18275
rect 32858 18272 32864 18284
rect 32723 18244 32864 18272
rect 32723 18241 32735 18244
rect 32677 18235 32735 18241
rect 32858 18232 32864 18244
rect 32916 18232 32922 18284
rect 33134 18232 33140 18284
rect 33192 18272 33198 18284
rect 33888 18281 33916 18312
rect 34054 18300 34060 18352
rect 34112 18340 34118 18352
rect 36630 18340 36636 18352
rect 34112 18312 34157 18340
rect 35360 18312 36636 18340
rect 34112 18300 34118 18312
rect 33689 18275 33747 18281
rect 33689 18272 33701 18275
rect 33192 18244 33701 18272
rect 33192 18232 33198 18244
rect 33689 18241 33701 18244
rect 33735 18241 33747 18275
rect 33689 18235 33747 18241
rect 33837 18275 33916 18281
rect 33837 18241 33849 18275
rect 33883 18244 33916 18275
rect 33965 18275 34023 18281
rect 33883 18241 33895 18244
rect 33837 18235 33895 18241
rect 33965 18241 33977 18275
rect 34011 18241 34023 18275
rect 33965 18235 34023 18241
rect 19614 18207 19672 18213
rect 19614 18173 19626 18207
rect 19660 18173 19672 18207
rect 19614 18167 19672 18173
rect 19116 18108 19564 18136
rect 19628 18136 19656 18167
rect 19702 18164 19708 18216
rect 19760 18204 19766 18216
rect 23198 18204 23204 18216
rect 19760 18176 19805 18204
rect 23159 18176 23204 18204
rect 19760 18164 19766 18176
rect 23198 18164 23204 18176
rect 23256 18164 23262 18216
rect 24210 18164 24216 18216
rect 24268 18204 24274 18216
rect 24268 18176 30144 18204
rect 24268 18164 24274 18176
rect 28166 18136 28172 18148
rect 19628 18108 23060 18136
rect 19116 18096 19122 18108
rect 15010 18068 15016 18080
rect 13004 18040 15016 18068
rect 8573 18031 8631 18037
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 15102 18028 15108 18080
rect 15160 18068 15166 18080
rect 18138 18068 18144 18080
rect 15160 18040 18144 18068
rect 15160 18028 15166 18040
rect 18138 18028 18144 18040
rect 18196 18028 18202 18080
rect 18598 18068 18604 18080
rect 18511 18040 18604 18068
rect 18598 18028 18604 18040
rect 18656 18068 18662 18080
rect 19150 18068 19156 18080
rect 18656 18040 19156 18068
rect 18656 18028 18662 18040
rect 19150 18028 19156 18040
rect 19208 18068 19214 18080
rect 19702 18068 19708 18080
rect 19208 18040 19708 18068
rect 19208 18028 19214 18040
rect 19702 18028 19708 18040
rect 19760 18028 19766 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20993 18071 21051 18077
rect 20993 18068 21005 18071
rect 20772 18040 21005 18068
rect 20772 18028 20778 18040
rect 20993 18037 21005 18040
rect 21039 18037 21051 18071
rect 21818 18068 21824 18080
rect 21779 18040 21824 18068
rect 20993 18031 21051 18037
rect 21818 18028 21824 18040
rect 21876 18028 21882 18080
rect 23032 18068 23060 18108
rect 27448 18108 28172 18136
rect 24578 18068 24584 18080
rect 23032 18040 24584 18068
rect 24578 18028 24584 18040
rect 24636 18028 24642 18080
rect 27448 18077 27476 18108
rect 28166 18096 28172 18108
rect 28224 18096 28230 18148
rect 30116 18145 30144 18176
rect 30374 18164 30380 18216
rect 30432 18204 30438 18216
rect 30745 18207 30803 18213
rect 30745 18204 30757 18207
rect 30432 18176 30757 18204
rect 30432 18164 30438 18176
rect 30745 18173 30757 18176
rect 30791 18173 30803 18207
rect 32398 18204 32404 18216
rect 32359 18176 32404 18204
rect 30745 18167 30803 18173
rect 32398 18164 32404 18176
rect 32456 18164 32462 18216
rect 30101 18139 30159 18145
rect 30101 18105 30113 18139
rect 30147 18105 30159 18139
rect 30101 18099 30159 18105
rect 33594 18096 33600 18148
rect 33652 18136 33658 18148
rect 33980 18136 34008 18235
rect 34146 18232 34152 18284
rect 34204 18281 34210 18284
rect 34204 18272 34212 18281
rect 34204 18244 34249 18272
rect 34204 18235 34212 18244
rect 34204 18232 34210 18235
rect 34422 18232 34428 18284
rect 34480 18272 34486 18284
rect 35360 18281 35388 18312
rect 35345 18275 35403 18281
rect 35345 18272 35357 18275
rect 34480 18244 35357 18272
rect 34480 18232 34486 18244
rect 35345 18241 35357 18244
rect 35391 18241 35403 18275
rect 35345 18235 35403 18241
rect 35434 18232 35440 18284
rect 35492 18272 35498 18284
rect 36372 18281 36400 18312
rect 36630 18300 36636 18312
rect 36688 18300 36694 18352
rect 36357 18275 36415 18281
rect 35492 18244 36308 18272
rect 35492 18232 35498 18244
rect 35713 18207 35771 18213
rect 35713 18173 35725 18207
rect 35759 18173 35771 18207
rect 36280 18204 36308 18244
rect 36357 18241 36369 18275
rect 36403 18241 36415 18275
rect 36357 18235 36415 18241
rect 36541 18275 36599 18281
rect 36541 18241 36553 18275
rect 36587 18272 36599 18275
rect 36740 18272 36768 18380
rect 43162 18368 43168 18420
rect 43220 18408 43226 18420
rect 43917 18411 43975 18417
rect 43917 18408 43929 18411
rect 43220 18380 43929 18408
rect 43220 18368 43226 18380
rect 43917 18377 43929 18380
rect 43963 18377 43975 18411
rect 44082 18408 44088 18420
rect 44043 18380 44088 18408
rect 43917 18371 43975 18377
rect 44082 18368 44088 18380
rect 44140 18368 44146 18420
rect 53377 18411 53435 18417
rect 53377 18377 53389 18411
rect 53423 18377 53435 18411
rect 55398 18408 55404 18420
rect 55359 18380 55404 18408
rect 53377 18371 53435 18377
rect 42610 18300 42616 18352
rect 42668 18340 42674 18352
rect 43717 18343 43775 18349
rect 43717 18340 43729 18343
rect 42668 18312 43729 18340
rect 42668 18300 42674 18312
rect 43717 18309 43729 18312
rect 43763 18309 43775 18343
rect 43717 18303 43775 18309
rect 46492 18312 47256 18340
rect 37182 18272 37188 18284
rect 36587 18244 37188 18272
rect 36587 18241 36599 18244
rect 36541 18235 36599 18241
rect 37182 18232 37188 18244
rect 37240 18272 37246 18284
rect 37553 18275 37611 18281
rect 37553 18272 37565 18275
rect 37240 18244 37565 18272
rect 37240 18232 37246 18244
rect 37553 18241 37565 18244
rect 37599 18241 37611 18275
rect 37553 18235 37611 18241
rect 43070 18232 43076 18284
rect 43128 18272 43134 18284
rect 46492 18272 46520 18312
rect 46658 18272 46664 18284
rect 43128 18244 46520 18272
rect 46619 18244 46664 18272
rect 43128 18232 43134 18244
rect 46658 18232 46664 18244
rect 46716 18232 46722 18284
rect 46845 18275 46903 18281
rect 46845 18241 46857 18275
rect 46891 18272 46903 18275
rect 47228 18272 47256 18312
rect 47302 18300 47308 18352
rect 47360 18340 47366 18352
rect 47826 18343 47884 18349
rect 47826 18340 47838 18343
rect 47360 18312 47838 18340
rect 47360 18300 47366 18312
rect 47826 18309 47838 18312
rect 47872 18309 47884 18343
rect 53392 18340 53420 18371
rect 55398 18368 55404 18380
rect 55456 18368 55462 18420
rect 54266 18343 54324 18349
rect 54266 18340 54278 18343
rect 53392 18312 54278 18340
rect 47826 18303 47884 18309
rect 54266 18309 54278 18312
rect 54312 18309 54324 18343
rect 54266 18303 54324 18309
rect 47578 18272 47584 18284
rect 46891 18244 47164 18272
rect 47228 18244 47584 18272
rect 46891 18241 46903 18244
rect 46845 18235 46903 18241
rect 36449 18207 36507 18213
rect 36449 18204 36461 18207
rect 36280 18176 36461 18204
rect 35713 18167 35771 18173
rect 36449 18173 36461 18176
rect 36495 18173 36507 18207
rect 36449 18167 36507 18173
rect 36633 18207 36691 18213
rect 36633 18173 36645 18207
rect 36679 18204 36691 18207
rect 36998 18204 37004 18216
rect 36679 18176 37004 18204
rect 36679 18173 36691 18176
rect 36633 18167 36691 18173
rect 33652 18108 34008 18136
rect 35728 18136 35756 18167
rect 35894 18136 35900 18148
rect 35728 18108 35900 18136
rect 33652 18096 33658 18108
rect 35894 18096 35900 18108
rect 35952 18136 35958 18148
rect 36648 18136 36676 18167
rect 36998 18164 37004 18176
rect 37056 18164 37062 18216
rect 37274 18204 37280 18216
rect 37235 18176 37280 18204
rect 37274 18164 37280 18176
rect 37332 18164 37338 18216
rect 35952 18108 36676 18136
rect 35952 18096 35958 18108
rect 27433 18071 27491 18077
rect 27433 18037 27445 18071
rect 27479 18037 27491 18071
rect 27433 18031 27491 18037
rect 27522 18028 27528 18080
rect 27580 18068 27586 18080
rect 27617 18071 27675 18077
rect 27617 18068 27629 18071
rect 27580 18040 27629 18068
rect 27580 18028 27586 18040
rect 27617 18037 27629 18040
rect 27663 18037 27675 18071
rect 27617 18031 27675 18037
rect 27706 18028 27712 18080
rect 27764 18068 27770 18080
rect 34333 18071 34391 18077
rect 34333 18068 34345 18071
rect 27764 18040 34345 18068
rect 27764 18028 27770 18040
rect 34333 18037 34345 18040
rect 34379 18037 34391 18071
rect 34333 18031 34391 18037
rect 35621 18071 35679 18077
rect 35621 18037 35633 18071
rect 35667 18068 35679 18071
rect 36078 18068 36084 18080
rect 35667 18040 36084 18068
rect 35667 18037 35679 18040
rect 35621 18031 35679 18037
rect 36078 18028 36084 18040
rect 36136 18028 36142 18080
rect 36173 18071 36231 18077
rect 36173 18037 36185 18071
rect 36219 18068 36231 18071
rect 36538 18068 36544 18080
rect 36219 18040 36544 18068
rect 36219 18037 36231 18040
rect 36173 18031 36231 18037
rect 36538 18028 36544 18040
rect 36596 18028 36602 18080
rect 43898 18068 43904 18080
rect 43859 18040 43904 18068
rect 43898 18028 43904 18040
rect 43956 18028 43962 18080
rect 47026 18068 47032 18080
rect 46987 18040 47032 18068
rect 47026 18028 47032 18040
rect 47084 18028 47090 18080
rect 47136 18068 47164 18244
rect 47578 18232 47584 18244
rect 47636 18232 47642 18284
rect 53558 18272 53564 18284
rect 53519 18244 53564 18272
rect 53558 18232 53564 18244
rect 53616 18232 53622 18284
rect 53374 18164 53380 18216
rect 53432 18204 53438 18216
rect 54021 18207 54079 18213
rect 54021 18204 54033 18207
rect 53432 18176 54033 18204
rect 53432 18164 53438 18176
rect 54021 18173 54033 18176
rect 54067 18173 54079 18207
rect 54021 18167 54079 18173
rect 47854 18068 47860 18080
rect 47136 18040 47860 18068
rect 47854 18028 47860 18040
rect 47912 18068 47918 18080
rect 48961 18071 49019 18077
rect 48961 18068 48973 18071
rect 47912 18040 48973 18068
rect 47912 18028 47918 18040
rect 48961 18037 48973 18040
rect 49007 18037 49019 18071
rect 48961 18031 49019 18037
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 6365 17867 6423 17873
rect 6365 17833 6377 17867
rect 6411 17864 6423 17867
rect 7098 17864 7104 17876
rect 6411 17836 7104 17864
rect 6411 17833 6423 17836
rect 6365 17827 6423 17833
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 8938 17824 8944 17876
rect 8996 17864 9002 17876
rect 16666 17864 16672 17876
rect 8996 17836 16672 17864
rect 8996 17824 9002 17836
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 16850 17824 16856 17876
rect 16908 17864 16914 17876
rect 18874 17864 18880 17876
rect 16908 17836 18880 17864
rect 16908 17824 16914 17836
rect 18874 17824 18880 17836
rect 18932 17824 18938 17876
rect 18966 17824 18972 17876
rect 19024 17864 19030 17876
rect 33873 17867 33931 17873
rect 33873 17864 33885 17867
rect 19024 17836 33885 17864
rect 19024 17824 19030 17836
rect 33873 17833 33885 17836
rect 33919 17833 33931 17867
rect 33873 17827 33931 17833
rect 37645 17867 37703 17873
rect 37645 17833 37657 17867
rect 37691 17864 37703 17867
rect 39206 17864 39212 17876
rect 37691 17836 39212 17864
rect 37691 17833 37703 17836
rect 37645 17827 37703 17833
rect 39206 17824 39212 17836
rect 39264 17824 39270 17876
rect 43070 17864 43076 17876
rect 41800 17836 43076 17864
rect 14274 17756 14280 17808
rect 14332 17796 14338 17808
rect 19978 17796 19984 17808
rect 14332 17768 19984 17796
rect 14332 17756 14338 17768
rect 19978 17756 19984 17768
rect 20036 17756 20042 17808
rect 22097 17799 22155 17805
rect 22097 17765 22109 17799
rect 22143 17796 22155 17799
rect 22186 17796 22192 17808
rect 22143 17768 22192 17796
rect 22143 17765 22155 17768
rect 22097 17759 22155 17765
rect 22186 17756 22192 17768
rect 22244 17756 22250 17808
rect 24394 17796 24400 17808
rect 24355 17768 24400 17796
rect 24394 17756 24400 17768
rect 24452 17756 24458 17808
rect 27154 17756 27160 17808
rect 27212 17796 27218 17808
rect 32398 17796 32404 17808
rect 27212 17768 32404 17796
rect 27212 17756 27218 17768
rect 32398 17756 32404 17768
rect 32456 17756 32462 17808
rect 37274 17796 37280 17808
rect 33612 17768 37280 17796
rect 2498 17688 2504 17740
rect 2556 17728 2562 17740
rect 2556 17700 3832 17728
rect 2556 17688 2562 17700
rect 3804 17672 3832 17700
rect 6546 17688 6552 17740
rect 6604 17728 6610 17740
rect 6825 17731 6883 17737
rect 6825 17728 6837 17731
rect 6604 17700 6837 17728
rect 6604 17688 6610 17700
rect 6825 17697 6837 17700
rect 6871 17697 6883 17731
rect 6825 17691 6883 17697
rect 6917 17731 6975 17737
rect 6917 17697 6929 17731
rect 6963 17697 6975 17731
rect 6917 17691 6975 17697
rect 1394 17660 1400 17672
rect 1355 17632 1400 17660
rect 1394 17620 1400 17632
rect 1452 17620 1458 17672
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17660 2191 17663
rect 3786 17660 3792 17672
rect 2179 17632 2774 17660
rect 3747 17632 3792 17660
rect 2179 17629 2191 17632
rect 2133 17623 2191 17629
rect 1578 17524 1584 17536
rect 1539 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 2314 17524 2320 17536
rect 2275 17496 2320 17524
rect 2314 17484 2320 17496
rect 2372 17484 2378 17536
rect 2746 17524 2774 17632
rect 3786 17620 3792 17632
rect 3844 17620 3850 17672
rect 6730 17620 6736 17672
rect 6788 17660 6794 17672
rect 6932 17660 6960 17691
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 8938 17728 8944 17740
rect 8352 17700 8944 17728
rect 8352 17688 8358 17700
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 16301 17731 16359 17737
rect 14568 17700 16160 17728
rect 6788 17632 6960 17660
rect 8956 17660 8984 17688
rect 11422 17660 11428 17672
rect 8956 17632 11428 17660
rect 6788 17620 6794 17632
rect 11422 17620 11428 17632
rect 11480 17620 11486 17672
rect 12526 17620 12532 17672
rect 12584 17660 12590 17672
rect 12986 17660 12992 17672
rect 12584 17632 12992 17660
rect 12584 17620 12590 17632
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 13446 17620 13452 17672
rect 13504 17660 13510 17672
rect 14568 17669 14596 17700
rect 14553 17663 14611 17669
rect 14553 17660 14565 17663
rect 13504 17632 14565 17660
rect 13504 17620 13510 17632
rect 14553 17629 14565 17632
rect 14599 17629 14611 17663
rect 15930 17660 15936 17672
rect 14553 17623 14611 17629
rect 14936 17632 15936 17660
rect 3878 17552 3884 17604
rect 3936 17592 3942 17604
rect 4034 17595 4092 17601
rect 4034 17592 4046 17595
rect 3936 17564 4046 17592
rect 3936 17552 3942 17564
rect 4034 17561 4046 17564
rect 4080 17561 4092 17595
rect 4034 17555 4092 17561
rect 5626 17552 5632 17604
rect 5684 17592 5690 17604
rect 5721 17595 5779 17601
rect 5721 17592 5733 17595
rect 5684 17564 5733 17592
rect 5684 17552 5690 17564
rect 5721 17561 5733 17564
rect 5767 17561 5779 17595
rect 5721 17555 5779 17561
rect 7834 17552 7840 17604
rect 7892 17592 7898 17604
rect 9186 17595 9244 17601
rect 9186 17592 9198 17595
rect 7892 17564 9198 17592
rect 7892 17552 7898 17564
rect 9186 17561 9198 17564
rect 9232 17561 9244 17595
rect 9186 17555 9244 17561
rect 13354 17552 13360 17604
rect 13412 17592 13418 17604
rect 14936 17592 14964 17632
rect 15930 17620 15936 17632
rect 15988 17660 15994 17672
rect 16025 17663 16083 17669
rect 16025 17660 16037 17663
rect 15988 17632 16037 17660
rect 15988 17620 15994 17632
rect 16025 17629 16037 17632
rect 16071 17629 16083 17663
rect 16132 17660 16160 17700
rect 16301 17697 16313 17731
rect 16347 17728 16359 17731
rect 16390 17728 16396 17740
rect 16347 17700 16396 17728
rect 16347 17697 16359 17700
rect 16301 17691 16359 17697
rect 16390 17688 16396 17700
rect 16448 17688 16454 17740
rect 16482 17688 16488 17740
rect 16540 17728 16546 17740
rect 17497 17731 17555 17737
rect 16540 17700 17448 17728
rect 16540 17688 16546 17700
rect 16850 17660 16856 17672
rect 16132 17632 16856 17660
rect 16025 17623 16083 17629
rect 16850 17620 16856 17632
rect 16908 17620 16914 17672
rect 16942 17620 16948 17672
rect 17000 17660 17006 17672
rect 17221 17663 17279 17669
rect 17221 17660 17233 17663
rect 17000 17632 17233 17660
rect 17000 17620 17006 17632
rect 17221 17629 17233 17632
rect 17267 17629 17279 17663
rect 17420 17660 17448 17700
rect 17497 17697 17509 17731
rect 17543 17728 17555 17731
rect 17678 17728 17684 17740
rect 17543 17700 17684 17728
rect 17543 17697 17555 17700
rect 17497 17691 17555 17697
rect 17678 17688 17684 17700
rect 17736 17688 17742 17740
rect 17770 17688 17776 17740
rect 17828 17728 17834 17740
rect 20530 17728 20536 17740
rect 17828 17700 20536 17728
rect 17828 17688 17834 17700
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 25516 17700 26280 17728
rect 18966 17660 18972 17672
rect 17420 17632 18972 17660
rect 17221 17623 17279 17629
rect 18966 17620 18972 17632
rect 19024 17620 19030 17672
rect 20162 17620 20168 17672
rect 20220 17660 20226 17672
rect 20717 17663 20775 17669
rect 20717 17660 20729 17663
rect 20220 17632 20729 17660
rect 20220 17620 20226 17632
rect 20717 17629 20729 17632
rect 20763 17629 20775 17663
rect 20717 17623 20775 17629
rect 20984 17663 21042 17669
rect 20984 17629 20996 17663
rect 21030 17660 21042 17663
rect 21818 17660 21824 17672
rect 21030 17632 21824 17660
rect 21030 17629 21042 17632
rect 20984 17623 21042 17629
rect 21818 17620 21824 17632
rect 21876 17620 21882 17672
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 24762 17660 24768 17672
rect 24627 17632 24768 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 24857 17663 24915 17669
rect 24857 17629 24869 17663
rect 24903 17660 24915 17663
rect 24946 17660 24952 17672
rect 24903 17632 24952 17660
rect 24903 17629 24915 17632
rect 24857 17623 24915 17629
rect 24946 17620 24952 17632
rect 25004 17620 25010 17672
rect 25516 17669 25544 17700
rect 25501 17663 25559 17669
rect 25501 17629 25513 17663
rect 25547 17629 25559 17663
rect 26145 17663 26203 17669
rect 26145 17660 26157 17663
rect 25501 17623 25559 17629
rect 25608 17632 26157 17660
rect 13412 17564 14964 17592
rect 13412 17552 13418 17564
rect 15010 17552 15016 17604
rect 15068 17592 15074 17604
rect 18782 17592 18788 17604
rect 15068 17564 18788 17592
rect 15068 17552 15074 17564
rect 18782 17552 18788 17564
rect 18840 17552 18846 17604
rect 18874 17552 18880 17604
rect 18932 17592 18938 17604
rect 20898 17592 20904 17604
rect 18932 17564 20904 17592
rect 18932 17552 18938 17564
rect 20898 17552 20904 17564
rect 20956 17552 20962 17604
rect 24780 17592 24808 17620
rect 25317 17595 25375 17601
rect 25317 17592 25329 17595
rect 24780 17564 25329 17592
rect 25317 17561 25329 17564
rect 25363 17561 25375 17595
rect 25317 17555 25375 17561
rect 25406 17552 25412 17604
rect 25464 17592 25470 17604
rect 25608 17592 25636 17632
rect 26145 17629 26157 17632
rect 26191 17629 26203 17663
rect 26252 17660 26280 17700
rect 28902 17688 28908 17740
rect 28960 17728 28966 17740
rect 28960 17700 29684 17728
rect 28960 17688 28966 17700
rect 27522 17660 27528 17672
rect 26252 17632 27528 17660
rect 26145 17623 26203 17629
rect 27522 17620 27528 17632
rect 27580 17620 27586 17672
rect 29086 17620 29092 17672
rect 29144 17660 29150 17672
rect 29454 17660 29460 17672
rect 29144 17632 29460 17660
rect 29144 17620 29150 17632
rect 29454 17620 29460 17632
rect 29512 17660 29518 17672
rect 29656 17669 29684 17700
rect 29730 17688 29736 17740
rect 29788 17728 29794 17740
rect 31113 17731 31171 17737
rect 31113 17728 31125 17731
rect 29788 17700 31125 17728
rect 29788 17688 29794 17700
rect 31113 17697 31125 17700
rect 31159 17697 31171 17731
rect 31113 17691 31171 17697
rect 31389 17731 31447 17737
rect 31389 17697 31401 17731
rect 31435 17728 31447 17731
rect 32582 17728 32588 17740
rect 31435 17700 32588 17728
rect 31435 17697 31447 17700
rect 31389 17691 31447 17697
rect 29549 17663 29607 17669
rect 29549 17660 29561 17663
rect 29512 17632 29561 17660
rect 29512 17620 29518 17632
rect 29549 17629 29561 17632
rect 29595 17629 29607 17663
rect 29549 17623 29607 17629
rect 29642 17663 29700 17669
rect 29642 17629 29654 17663
rect 29688 17629 29700 17663
rect 29642 17623 29700 17629
rect 30006 17620 30012 17672
rect 30064 17669 30070 17672
rect 30064 17660 30072 17669
rect 30064 17632 30109 17660
rect 30064 17623 30072 17632
rect 30064 17620 30070 17623
rect 25464 17564 25636 17592
rect 25464 17552 25470 17564
rect 25958 17552 25964 17604
rect 26016 17592 26022 17604
rect 26390 17595 26448 17601
rect 26390 17592 26402 17595
rect 26016 17564 26402 17592
rect 26016 17552 26022 17564
rect 26390 17561 26402 17564
rect 26436 17561 26448 17595
rect 26390 17555 26448 17561
rect 26510 17552 26516 17604
rect 26568 17592 26574 17604
rect 29822 17592 29828 17604
rect 26568 17564 29684 17592
rect 29783 17564 29828 17592
rect 26568 17552 26574 17564
rect 4154 17524 4160 17536
rect 2746 17496 4160 17524
rect 4154 17484 4160 17496
rect 4212 17524 4218 17536
rect 5169 17527 5227 17533
rect 5169 17524 5181 17527
rect 4212 17496 5181 17524
rect 4212 17484 4218 17496
rect 5169 17493 5181 17496
rect 5215 17493 5227 17527
rect 5810 17524 5816 17536
rect 5771 17496 5816 17524
rect 5169 17487 5227 17493
rect 5810 17484 5816 17496
rect 5868 17484 5874 17536
rect 6362 17484 6368 17536
rect 6420 17524 6426 17536
rect 6733 17527 6791 17533
rect 6733 17524 6745 17527
rect 6420 17496 6745 17524
rect 6420 17484 6426 17496
rect 6733 17493 6745 17496
rect 6779 17524 6791 17527
rect 6822 17524 6828 17536
rect 6779 17496 6828 17524
rect 6779 17493 6791 17496
rect 6733 17487 6791 17493
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 10318 17524 10324 17536
rect 10279 17496 10324 17524
rect 10318 17484 10324 17496
rect 10376 17484 10382 17536
rect 14829 17527 14887 17533
rect 14829 17493 14841 17527
rect 14875 17524 14887 17527
rect 15286 17524 15292 17536
rect 14875 17496 15292 17524
rect 14875 17493 14887 17496
rect 14829 17487 14887 17493
rect 15286 17484 15292 17496
rect 15344 17524 15350 17536
rect 15838 17524 15844 17536
rect 15344 17496 15844 17524
rect 15344 17484 15350 17496
rect 15838 17484 15844 17496
rect 15896 17484 15902 17536
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 20806 17524 20812 17536
rect 16540 17496 20812 17524
rect 16540 17484 16546 17496
rect 20806 17484 20812 17496
rect 20864 17484 20870 17536
rect 24578 17484 24584 17536
rect 24636 17524 24642 17536
rect 24765 17527 24823 17533
rect 24765 17524 24777 17527
rect 24636 17496 24777 17524
rect 24636 17484 24642 17496
rect 24765 17493 24777 17496
rect 24811 17493 24823 17527
rect 24765 17487 24823 17493
rect 25685 17527 25743 17533
rect 25685 17493 25697 17527
rect 25731 17524 25743 17527
rect 26142 17524 26148 17536
rect 25731 17496 26148 17524
rect 25731 17493 25743 17496
rect 25685 17487 25743 17493
rect 26142 17484 26148 17496
rect 26200 17484 26206 17536
rect 27525 17527 27583 17533
rect 27525 17493 27537 17527
rect 27571 17524 27583 17527
rect 28442 17524 28448 17536
rect 27571 17496 28448 17524
rect 27571 17493 27583 17496
rect 27525 17487 27583 17493
rect 28442 17484 28448 17496
rect 28500 17484 28506 17536
rect 29656 17524 29684 17564
rect 29822 17552 29828 17564
rect 29880 17552 29886 17604
rect 29914 17552 29920 17604
rect 29972 17592 29978 17604
rect 30374 17592 30380 17604
rect 29972 17564 30017 17592
rect 30116 17564 30380 17592
rect 29972 17552 29978 17564
rect 30116 17524 30144 17564
rect 30374 17552 30380 17564
rect 30432 17552 30438 17604
rect 29656 17496 30144 17524
rect 30190 17484 30196 17536
rect 30248 17524 30254 17536
rect 31128 17524 31156 17691
rect 32582 17688 32588 17700
rect 32640 17688 32646 17740
rect 33134 17620 33140 17672
rect 33192 17660 33198 17672
rect 33229 17663 33287 17669
rect 33229 17660 33241 17663
rect 33192 17632 33241 17660
rect 33192 17620 33198 17632
rect 33229 17629 33241 17632
rect 33275 17629 33287 17663
rect 33229 17623 33287 17629
rect 33377 17663 33435 17669
rect 33377 17629 33389 17663
rect 33423 17660 33435 17663
rect 33612 17660 33640 17768
rect 37274 17756 37280 17768
rect 37332 17756 37338 17808
rect 36906 17688 36912 17740
rect 36964 17728 36970 17740
rect 37185 17731 37243 17737
rect 37185 17728 37197 17731
rect 36964 17700 37197 17728
rect 36964 17688 36970 17700
rect 37185 17697 37197 17700
rect 37231 17697 37243 17731
rect 37826 17728 37832 17740
rect 37787 17700 37832 17728
rect 37185 17691 37243 17697
rect 37826 17688 37832 17700
rect 37884 17688 37890 17740
rect 37921 17731 37979 17737
rect 37921 17697 37933 17731
rect 37967 17728 37979 17731
rect 38930 17728 38936 17740
rect 37967 17700 38936 17728
rect 37967 17697 37979 17700
rect 37921 17691 37979 17697
rect 38930 17688 38936 17700
rect 38988 17688 38994 17740
rect 33423 17632 33640 17660
rect 33735 17663 33793 17669
rect 33423 17629 33435 17632
rect 33377 17623 33435 17629
rect 33735 17629 33747 17663
rect 33781 17660 33793 17663
rect 33870 17660 33876 17672
rect 33781 17632 33876 17660
rect 33781 17629 33793 17632
rect 33735 17623 33793 17629
rect 33870 17620 33876 17632
rect 33928 17620 33934 17672
rect 34790 17620 34796 17672
rect 34848 17660 34854 17672
rect 36722 17660 36728 17672
rect 34848 17632 36728 17660
rect 34848 17620 34854 17632
rect 36722 17620 36728 17632
rect 36780 17620 36786 17672
rect 36817 17663 36875 17669
rect 36817 17629 36829 17663
rect 36863 17660 36875 17663
rect 36998 17660 37004 17672
rect 36863 17632 37004 17660
rect 36863 17629 36875 17632
rect 36817 17623 36875 17629
rect 36998 17620 37004 17632
rect 37056 17620 37062 17672
rect 38010 17660 38016 17672
rect 37971 17632 38016 17660
rect 38010 17620 38016 17632
rect 38068 17620 38074 17672
rect 38105 17663 38163 17669
rect 38105 17629 38117 17663
rect 38151 17660 38163 17663
rect 38194 17660 38200 17672
rect 38151 17632 38200 17660
rect 38151 17629 38163 17632
rect 38105 17623 38163 17629
rect 38194 17620 38200 17632
rect 38252 17620 38258 17672
rect 38562 17620 38568 17672
rect 38620 17660 38626 17672
rect 40773 17663 40831 17669
rect 40773 17660 40785 17663
rect 38620 17632 40785 17660
rect 38620 17620 38626 17632
rect 40773 17629 40785 17632
rect 40819 17660 40831 17663
rect 41800 17660 41828 17836
rect 43070 17824 43076 17836
rect 43128 17824 43134 17876
rect 43898 17864 43904 17876
rect 43859 17836 43904 17864
rect 43898 17824 43904 17836
rect 43956 17824 43962 17876
rect 47026 17864 47032 17876
rect 46987 17836 47032 17864
rect 47026 17824 47032 17836
rect 47084 17824 47090 17876
rect 47213 17867 47271 17873
rect 47213 17833 47225 17867
rect 47259 17864 47271 17867
rect 47486 17864 47492 17876
rect 47259 17836 47492 17864
rect 47259 17833 47271 17836
rect 47213 17827 47271 17833
rect 47486 17824 47492 17836
rect 47544 17824 47550 17876
rect 42794 17756 42800 17808
rect 42852 17796 42858 17808
rect 42852 17768 43116 17796
rect 42852 17756 42858 17768
rect 43088 17728 43116 17768
rect 44177 17731 44235 17737
rect 44177 17728 44189 17731
rect 42628 17700 43024 17728
rect 43088 17700 44189 17728
rect 42628 17672 42656 17700
rect 42610 17660 42616 17672
rect 40819 17632 41828 17660
rect 42571 17632 42616 17660
rect 40819 17629 40831 17632
rect 40773 17623 40831 17629
rect 42610 17620 42616 17632
rect 42668 17620 42674 17672
rect 42797 17663 42855 17669
rect 42797 17629 42809 17663
rect 42843 17629 42855 17663
rect 42797 17623 42855 17629
rect 32398 17552 32404 17604
rect 32456 17592 32462 17604
rect 33502 17592 33508 17604
rect 32456 17564 33508 17592
rect 32456 17552 32462 17564
rect 33502 17552 33508 17564
rect 33560 17552 33566 17604
rect 33597 17595 33655 17601
rect 33597 17561 33609 17595
rect 33643 17592 33655 17595
rect 34330 17592 34336 17604
rect 33643 17564 34336 17592
rect 33643 17561 33655 17564
rect 33597 17555 33655 17561
rect 34330 17552 34336 17564
rect 34388 17552 34394 17604
rect 37093 17595 37151 17601
rect 37093 17561 37105 17595
rect 37139 17592 37151 17595
rect 38286 17592 38292 17604
rect 37139 17564 38292 17592
rect 37139 17561 37151 17564
rect 37093 17555 37151 17561
rect 38286 17552 38292 17564
rect 38344 17552 38350 17604
rect 32122 17524 32128 17536
rect 30248 17496 30293 17524
rect 31128 17496 32128 17524
rect 30248 17484 30254 17496
rect 32122 17484 32128 17496
rect 32180 17484 32186 17536
rect 36262 17484 36268 17536
rect 36320 17524 36326 17536
rect 36541 17527 36599 17533
rect 36541 17524 36553 17527
rect 36320 17496 36553 17524
rect 36320 17484 36326 17496
rect 36541 17493 36553 17496
rect 36587 17493 36599 17527
rect 36541 17487 36599 17493
rect 37001 17527 37059 17533
rect 37001 17493 37013 17527
rect 37047 17524 37059 17527
rect 37182 17524 37188 17536
rect 37047 17496 37188 17524
rect 37047 17493 37059 17496
rect 37001 17487 37059 17493
rect 37182 17484 37188 17496
rect 37240 17484 37246 17536
rect 37550 17484 37556 17536
rect 37608 17524 37614 17536
rect 38580 17524 38608 17620
rect 41040 17595 41098 17601
rect 41040 17561 41052 17595
rect 41086 17592 41098 17595
rect 42812 17592 42840 17623
rect 41086 17564 42840 17592
rect 42996 17592 43024 17700
rect 44177 17697 44189 17700
rect 44223 17697 44235 17731
rect 44177 17691 44235 17697
rect 44269 17731 44327 17737
rect 44269 17697 44281 17731
rect 44315 17728 44327 17731
rect 44450 17728 44456 17740
rect 44315 17700 44456 17728
rect 44315 17697 44327 17700
rect 44269 17691 44327 17697
rect 44450 17688 44456 17700
rect 44508 17688 44514 17740
rect 43073 17663 43131 17669
rect 43073 17629 43085 17663
rect 43119 17660 43131 17663
rect 43162 17660 43168 17672
rect 43119 17632 43168 17660
rect 43119 17629 43131 17632
rect 43073 17623 43131 17629
rect 43162 17620 43168 17632
rect 43220 17620 43226 17672
rect 44082 17620 44088 17672
rect 44140 17660 44146 17672
rect 44358 17660 44364 17672
rect 44140 17632 44185 17660
rect 44319 17632 44364 17660
rect 44140 17620 44146 17632
rect 44358 17620 44364 17632
rect 44416 17620 44422 17672
rect 46658 17620 46664 17672
rect 46716 17660 46722 17672
rect 47673 17663 47731 17669
rect 47673 17660 47685 17663
rect 46716 17632 47685 17660
rect 46716 17620 46722 17632
rect 47673 17629 47685 17632
rect 47719 17629 47731 17663
rect 47854 17660 47860 17672
rect 47815 17632 47860 17660
rect 47673 17623 47731 17629
rect 47854 17620 47860 17632
rect 47912 17620 47918 17672
rect 46845 17595 46903 17601
rect 46845 17592 46857 17595
rect 42996 17564 46857 17592
rect 41086 17561 41098 17564
rect 41040 17555 41098 17561
rect 46845 17561 46857 17564
rect 46891 17592 46903 17595
rect 46934 17592 46940 17604
rect 46891 17564 46940 17592
rect 46891 17561 46903 17564
rect 46845 17555 46903 17561
rect 46934 17552 46940 17564
rect 46992 17552 46998 17604
rect 47061 17595 47119 17601
rect 47061 17561 47073 17595
rect 47107 17592 47119 17595
rect 47765 17595 47823 17601
rect 47765 17592 47777 17595
rect 47107 17564 47777 17592
rect 47107 17561 47119 17564
rect 47061 17555 47119 17561
rect 47765 17561 47777 17564
rect 47811 17561 47823 17595
rect 47765 17555 47823 17561
rect 42150 17524 42156 17536
rect 37608 17496 38608 17524
rect 42111 17496 42156 17524
rect 37608 17484 37614 17496
rect 42150 17484 42156 17496
rect 42208 17484 42214 17536
rect 42518 17484 42524 17536
rect 42576 17524 42582 17536
rect 42981 17527 43039 17533
rect 42981 17524 42993 17527
rect 42576 17496 42993 17524
rect 42576 17484 42582 17496
rect 42981 17493 42993 17496
rect 43027 17493 43039 17527
rect 42981 17487 43039 17493
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 3789 17323 3847 17329
rect 3789 17289 3801 17323
rect 3835 17320 3847 17323
rect 3878 17320 3884 17332
rect 3835 17292 3884 17320
rect 3835 17289 3847 17292
rect 3789 17283 3847 17289
rect 3878 17280 3884 17292
rect 3936 17280 3942 17332
rect 4154 17320 4160 17332
rect 4115 17292 4160 17320
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 7009 17323 7067 17329
rect 7009 17289 7021 17323
rect 7055 17289 7067 17323
rect 7834 17320 7840 17332
rect 7795 17292 7840 17320
rect 7009 17283 7067 17289
rect 2774 17212 2780 17264
rect 2832 17252 2838 17264
rect 7024 17252 7052 17283
rect 7834 17280 7840 17292
rect 7892 17280 7898 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17320 13231 17323
rect 16482 17320 16488 17332
rect 13219 17292 16488 17320
rect 13219 17289 13231 17292
rect 13173 17283 13231 17289
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 16666 17320 16672 17332
rect 16627 17292 16672 17320
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 16776 17292 18000 17320
rect 7650 17252 7656 17264
rect 2832 17224 4292 17252
rect 7024 17224 7656 17252
rect 2832 17212 2838 17224
rect 1854 17184 1860 17196
rect 1815 17156 1860 17184
rect 1854 17144 1860 17156
rect 1912 17144 1918 17196
rect 2866 17184 2872 17196
rect 2827 17156 2872 17184
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 3970 17184 3976 17196
rect 3931 17156 3976 17184
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 4264 17193 4292 17224
rect 7650 17212 7656 17224
rect 7708 17252 7714 17264
rect 10318 17252 10324 17264
rect 7708 17224 10324 17252
rect 7708 17212 7714 17224
rect 10318 17212 10324 17224
rect 10376 17212 10382 17264
rect 12802 17252 12808 17264
rect 12763 17224 12808 17252
rect 12802 17212 12808 17224
rect 12860 17212 12866 17264
rect 12989 17255 13047 17261
rect 12989 17221 13001 17255
rect 13035 17252 13047 17255
rect 14366 17252 14372 17264
rect 13035 17224 14372 17252
rect 13035 17221 13047 17224
rect 12989 17215 13047 17221
rect 14366 17212 14372 17224
rect 14424 17212 14430 17264
rect 16114 17212 16120 17264
rect 16172 17252 16178 17264
rect 16776 17252 16804 17292
rect 17862 17252 17868 17264
rect 16172 17224 16804 17252
rect 16868 17224 17868 17252
rect 16172 17212 16178 17224
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17184 4307 17187
rect 5810 17184 5816 17196
rect 4295 17156 5816 17184
rect 4295 17153 4307 17156
rect 4249 17147 4307 17153
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 16868 17193 16896 17224
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 8021 17187 8079 17193
rect 6788 17156 7236 17184
rect 6788 17144 6794 17156
rect 7208 17125 7236 17156
rect 8021 17153 8033 17187
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17153 16911 17187
rect 17126 17184 17132 17196
rect 17039 17156 17132 17184
rect 16853 17147 16911 17153
rect 7101 17119 7159 17125
rect 7101 17116 7113 17119
rect 4908 17088 7113 17116
rect 2685 17051 2743 17057
rect 2685 17017 2697 17051
rect 2731 17048 2743 17051
rect 4908 17048 4936 17088
rect 7101 17085 7113 17088
rect 7147 17085 7159 17119
rect 7101 17079 7159 17085
rect 7193 17119 7251 17125
rect 7193 17085 7205 17119
rect 7239 17085 7251 17119
rect 7193 17079 7251 17085
rect 2731 17020 4936 17048
rect 6641 17051 6699 17057
rect 2731 17017 2743 17020
rect 2685 17011 2743 17017
rect 6641 17017 6653 17051
rect 6687 17048 6699 17051
rect 8036 17048 8064 17147
rect 17126 17144 17132 17156
rect 17184 17184 17190 17196
rect 17678 17184 17684 17196
rect 17184 17156 17684 17184
rect 17184 17144 17190 17156
rect 17678 17144 17684 17156
rect 17736 17144 17742 17196
rect 13725 17119 13783 17125
rect 13725 17085 13737 17119
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17116 14059 17119
rect 14274 17116 14280 17128
rect 14047 17088 14280 17116
rect 14047 17085 14059 17088
rect 14001 17079 14059 17085
rect 13740 17048 13768 17079
rect 14274 17076 14280 17088
rect 14332 17116 14338 17128
rect 14826 17116 14832 17128
rect 14332 17088 14832 17116
rect 14332 17076 14338 17088
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 15010 17116 15016 17128
rect 14971 17088 15016 17116
rect 15010 17076 15016 17088
rect 15068 17076 15074 17128
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17116 15347 17119
rect 15930 17116 15936 17128
rect 15335 17088 15936 17116
rect 15335 17085 15347 17088
rect 15289 17079 15347 17085
rect 15930 17076 15936 17088
rect 15988 17076 15994 17128
rect 16945 17119 17003 17125
rect 16945 17085 16957 17119
rect 16991 17085 17003 17119
rect 16945 17079 17003 17085
rect 17037 17119 17095 17125
rect 17037 17085 17049 17119
rect 17083 17116 17095 17119
rect 17586 17116 17592 17128
rect 17083 17088 17592 17116
rect 17083 17085 17095 17088
rect 17037 17079 17095 17085
rect 6687 17020 8064 17048
rect 13004 17020 13768 17048
rect 16960 17048 16988 17079
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 17862 17116 17868 17128
rect 17823 17088 17868 17116
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 17972 17125 18000 17292
rect 18322 17280 18328 17332
rect 18380 17320 18386 17332
rect 18693 17323 18751 17329
rect 18693 17320 18705 17323
rect 18380 17292 18705 17320
rect 18380 17280 18386 17292
rect 18693 17289 18705 17292
rect 18739 17289 18751 17323
rect 18693 17283 18751 17289
rect 18782 17280 18788 17332
rect 18840 17320 18846 17332
rect 31938 17320 31944 17332
rect 18840 17292 31944 17320
rect 18840 17280 18846 17292
rect 31938 17280 31944 17292
rect 31996 17280 32002 17332
rect 35894 17320 35900 17332
rect 33336 17292 35900 17320
rect 20622 17252 20628 17264
rect 18064 17224 20628 17252
rect 18064 17193 18092 17224
rect 20622 17212 20628 17224
rect 20680 17212 20686 17264
rect 23198 17212 23204 17264
rect 23256 17252 23262 17264
rect 25406 17252 25412 17264
rect 23256 17224 25412 17252
rect 23256 17212 23262 17224
rect 25406 17212 25412 17224
rect 25464 17212 25470 17264
rect 25516 17224 33088 17252
rect 18049 17187 18107 17193
rect 18049 17153 18061 17187
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 18230 17144 18236 17196
rect 18288 17184 18294 17196
rect 18966 17184 18972 17196
rect 18288 17156 18972 17184
rect 18288 17144 18294 17156
rect 18966 17144 18972 17156
rect 19024 17144 19030 17196
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17184 19119 17187
rect 19107 17156 19334 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 17957 17119 18015 17125
rect 17957 17085 17969 17119
rect 18003 17085 18015 17119
rect 17957 17079 18015 17085
rect 18138 17076 18144 17128
rect 18196 17116 18202 17128
rect 18598 17116 18604 17128
rect 18196 17088 18604 17116
rect 18196 17076 18202 17088
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 18690 17076 18696 17128
rect 18748 17116 18754 17128
rect 18877 17119 18935 17125
rect 18877 17116 18889 17119
rect 18748 17088 18889 17116
rect 18748 17076 18754 17088
rect 18877 17085 18889 17088
rect 18923 17085 18935 17119
rect 19150 17116 19156 17128
rect 19111 17088 19156 17116
rect 18877 17079 18935 17085
rect 19150 17076 19156 17088
rect 19208 17076 19214 17128
rect 19306 17116 19334 17156
rect 20530 17144 20536 17196
rect 20588 17184 20594 17196
rect 23014 17184 23020 17196
rect 20588 17156 23020 17184
rect 20588 17144 20594 17156
rect 23014 17144 23020 17156
rect 23072 17144 23078 17196
rect 25516 17116 25544 17224
rect 26142 17184 26148 17196
rect 26103 17156 26148 17184
rect 26142 17144 26148 17156
rect 26200 17144 26206 17196
rect 29086 17144 29092 17196
rect 29144 17184 29150 17196
rect 29181 17187 29239 17193
rect 29181 17184 29193 17187
rect 29144 17156 29193 17184
rect 29144 17144 29150 17156
rect 29181 17153 29193 17156
rect 29227 17153 29239 17187
rect 29181 17147 29239 17153
rect 29274 17187 29332 17193
rect 29274 17153 29286 17187
rect 29320 17153 29332 17187
rect 29454 17184 29460 17196
rect 29415 17156 29460 17184
rect 29274 17147 29332 17153
rect 19306 17088 25544 17116
rect 28442 17076 28448 17128
rect 28500 17116 28506 17128
rect 29288 17116 29316 17147
rect 29454 17144 29460 17156
rect 29512 17144 29518 17196
rect 29546 17144 29552 17196
rect 29604 17184 29610 17196
rect 29687 17187 29745 17193
rect 29604 17156 29649 17184
rect 29604 17144 29610 17156
rect 29687 17153 29699 17187
rect 29733 17184 29745 17187
rect 30006 17184 30012 17196
rect 29733 17156 30012 17184
rect 29733 17153 29745 17156
rect 29687 17147 29745 17153
rect 30006 17144 30012 17156
rect 30064 17184 30070 17196
rect 32122 17184 32128 17196
rect 30064 17156 30604 17184
rect 32083 17156 32128 17184
rect 30064 17144 30070 17156
rect 28500 17088 29316 17116
rect 29472 17116 29500 17144
rect 29822 17116 29828 17128
rect 29472 17088 29828 17116
rect 28500 17076 28506 17088
rect 29822 17076 29828 17088
rect 29880 17076 29886 17128
rect 30285 17119 30343 17125
rect 30285 17085 30297 17119
rect 30331 17116 30343 17119
rect 30374 17116 30380 17128
rect 30331 17088 30380 17116
rect 30331 17085 30343 17088
rect 30285 17079 30343 17085
rect 30374 17076 30380 17088
rect 30432 17076 30438 17128
rect 30576 17125 30604 17156
rect 32122 17144 32128 17156
rect 32180 17144 32186 17196
rect 30561 17119 30619 17125
rect 30561 17085 30573 17119
rect 30607 17116 30619 17119
rect 31478 17116 31484 17128
rect 30607 17088 31484 17116
rect 30607 17085 30619 17088
rect 30561 17079 30619 17085
rect 31478 17076 31484 17088
rect 31536 17076 31542 17128
rect 33060 17116 33088 17224
rect 33134 17144 33140 17196
rect 33192 17184 33198 17196
rect 33336 17193 33364 17292
rect 35894 17280 35900 17292
rect 35952 17280 35958 17332
rect 36078 17280 36084 17332
rect 36136 17320 36142 17332
rect 36557 17323 36615 17329
rect 36557 17320 36569 17323
rect 36136 17292 36569 17320
rect 36136 17280 36142 17292
rect 36557 17289 36569 17292
rect 36603 17289 36615 17323
rect 42518 17320 42524 17332
rect 42479 17292 42524 17320
rect 36557 17283 36615 17289
rect 42518 17280 42524 17292
rect 42576 17280 42582 17332
rect 43162 17280 43168 17332
rect 43220 17320 43226 17332
rect 44177 17323 44235 17329
rect 44177 17320 44189 17323
rect 43220 17292 44189 17320
rect 43220 17280 43226 17292
rect 44177 17289 44189 17292
rect 44223 17289 44235 17323
rect 44177 17283 44235 17289
rect 33502 17252 33508 17264
rect 33463 17224 33508 17252
rect 33502 17212 33508 17224
rect 33560 17212 33566 17264
rect 33597 17255 33655 17261
rect 33597 17221 33609 17255
rect 33643 17252 33655 17255
rect 34422 17252 34428 17264
rect 33643 17224 34428 17252
rect 33643 17221 33655 17224
rect 33597 17215 33655 17221
rect 34422 17212 34428 17224
rect 34480 17212 34486 17264
rect 36357 17255 36415 17261
rect 36357 17221 36369 17255
rect 36403 17221 36415 17255
rect 36357 17215 36415 17221
rect 33229 17187 33287 17193
rect 33229 17184 33241 17187
rect 33192 17156 33241 17184
rect 33192 17144 33198 17156
rect 33229 17153 33241 17156
rect 33275 17153 33287 17187
rect 33229 17147 33287 17153
rect 33322 17187 33380 17193
rect 33322 17153 33334 17187
rect 33368 17153 33380 17187
rect 33322 17147 33380 17153
rect 33735 17187 33793 17193
rect 33735 17153 33747 17187
rect 33781 17184 33793 17187
rect 33870 17184 33876 17196
rect 33781 17156 33876 17184
rect 33781 17153 33793 17156
rect 33735 17147 33793 17153
rect 33870 17144 33876 17156
rect 33928 17144 33934 17196
rect 36372 17184 36400 17215
rect 36446 17212 36452 17264
rect 36504 17252 36510 17264
rect 42978 17252 42984 17264
rect 36504 17224 42984 17252
rect 36504 17212 36510 17224
rect 42978 17212 42984 17224
rect 43036 17212 43042 17264
rect 44082 17252 44088 17264
rect 44043 17224 44088 17252
rect 44082 17212 44088 17224
rect 44140 17212 44146 17264
rect 44269 17255 44327 17261
rect 44269 17221 44281 17255
rect 44315 17252 44327 17255
rect 44450 17252 44456 17264
rect 44315 17224 44456 17252
rect 44315 17221 44327 17224
rect 44269 17215 44327 17221
rect 44450 17212 44456 17224
rect 44508 17252 44514 17264
rect 45278 17252 45284 17264
rect 44508 17224 45284 17252
rect 44508 17212 44514 17224
rect 45278 17212 45284 17224
rect 45336 17252 45342 17264
rect 47854 17252 47860 17264
rect 45336 17224 47860 17252
rect 45336 17212 45342 17224
rect 47854 17212 47860 17224
rect 47912 17212 47918 17264
rect 36630 17184 36636 17196
rect 36372 17156 36636 17184
rect 36630 17144 36636 17156
rect 36688 17144 36694 17196
rect 41690 17144 41696 17196
rect 41748 17184 41754 17196
rect 42150 17184 42156 17196
rect 41748 17156 42156 17184
rect 41748 17144 41754 17156
rect 42150 17144 42156 17156
rect 42208 17184 42214 17196
rect 42429 17187 42487 17193
rect 42429 17184 42441 17187
rect 42208 17156 42441 17184
rect 42208 17144 42214 17156
rect 42429 17153 42441 17156
rect 42475 17153 42487 17187
rect 44358 17184 44364 17196
rect 44319 17156 44364 17184
rect 42429 17147 42487 17153
rect 44358 17144 44364 17156
rect 44416 17144 44422 17196
rect 51442 17184 51448 17196
rect 51403 17156 51448 17184
rect 51442 17144 51448 17156
rect 51500 17144 51506 17196
rect 34606 17116 34612 17128
rect 33060 17088 34612 17116
rect 34606 17076 34612 17088
rect 34664 17076 34670 17128
rect 16960 17020 19564 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 2133 16983 2191 16989
rect 2133 16949 2145 16983
rect 2179 16980 2191 16983
rect 7558 16980 7564 16992
rect 2179 16952 7564 16980
rect 2179 16949 2191 16952
rect 2133 16943 2191 16949
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 13004 16989 13032 17020
rect 12989 16983 13047 16989
rect 12989 16980 13001 16983
rect 10744 16952 13001 16980
rect 10744 16940 10750 16952
rect 12989 16949 13001 16952
rect 13035 16949 13047 16983
rect 12989 16943 13047 16949
rect 16850 16940 16856 16992
rect 16908 16980 16914 16992
rect 17681 16983 17739 16989
rect 17681 16980 17693 16983
rect 16908 16952 17693 16980
rect 16908 16940 16914 16952
rect 17681 16949 17693 16952
rect 17727 16949 17739 16983
rect 19536 16980 19564 17020
rect 19978 17008 19984 17060
rect 20036 17048 20042 17060
rect 33873 17051 33931 17057
rect 33873 17048 33885 17051
rect 20036 17020 33885 17048
rect 20036 17008 20042 17020
rect 33873 17017 33885 17020
rect 33919 17017 33931 17051
rect 33873 17011 33931 17017
rect 25774 16980 25780 16992
rect 19536 16952 25780 16980
rect 17681 16943 17739 16949
rect 25774 16940 25780 16952
rect 25832 16940 25838 16992
rect 25958 16980 25964 16992
rect 25919 16952 25964 16980
rect 25958 16940 25964 16952
rect 26016 16940 26022 16992
rect 27246 16940 27252 16992
rect 27304 16980 27310 16992
rect 29825 16983 29883 16989
rect 29825 16980 29837 16983
rect 27304 16952 29837 16980
rect 27304 16940 27310 16952
rect 29825 16949 29837 16952
rect 29871 16949 29883 16983
rect 32306 16980 32312 16992
rect 32267 16952 32312 16980
rect 29825 16943 29883 16949
rect 32306 16940 32312 16952
rect 32364 16980 32370 16992
rect 33134 16980 33140 16992
rect 32364 16952 33140 16980
rect 32364 16940 32370 16952
rect 33134 16940 33140 16952
rect 33192 16940 33198 16992
rect 36538 16980 36544 16992
rect 36499 16952 36544 16980
rect 36538 16940 36544 16952
rect 36596 16940 36602 16992
rect 36725 16983 36783 16989
rect 36725 16949 36737 16983
rect 36771 16980 36783 16983
rect 37090 16980 37096 16992
rect 36771 16952 37096 16980
rect 36771 16949 36783 16952
rect 36725 16943 36783 16949
rect 37090 16940 37096 16952
rect 37148 16940 37154 16992
rect 51074 16940 51080 16992
rect 51132 16980 51138 16992
rect 51261 16983 51319 16989
rect 51261 16980 51273 16983
rect 51132 16952 51273 16980
rect 51132 16940 51138 16952
rect 51261 16949 51273 16952
rect 51307 16949 51319 16983
rect 51261 16943 51319 16949
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 7558 16736 7564 16788
rect 7616 16776 7622 16788
rect 7616 16748 14228 16776
rect 7616 16736 7622 16748
rect 3970 16668 3976 16720
rect 4028 16708 4034 16720
rect 9950 16708 9956 16720
rect 4028 16680 9956 16708
rect 4028 16668 4034 16680
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 14200 16708 14228 16748
rect 14274 16736 14280 16788
rect 14332 16776 14338 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 14332 16748 14381 16776
rect 14332 16736 14338 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 16666 16776 16672 16788
rect 14369 16739 14427 16745
rect 14476 16748 16672 16776
rect 14476 16708 14504 16748
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 16960 16748 22094 16776
rect 14200 16680 14504 16708
rect 1486 16600 1492 16652
rect 1544 16640 1550 16652
rect 1581 16643 1639 16649
rect 1581 16640 1593 16643
rect 1544 16612 1593 16640
rect 1544 16600 1550 16612
rect 1581 16609 1593 16612
rect 1627 16609 1639 16643
rect 1581 16603 1639 16609
rect 11422 16600 11428 16652
rect 11480 16640 11486 16652
rect 12158 16640 12164 16652
rect 11480 16612 12164 16640
rect 11480 16600 11486 16612
rect 12158 16600 12164 16612
rect 12216 16600 12222 16652
rect 16114 16640 16120 16652
rect 16075 16612 16120 16640
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 16850 16640 16856 16652
rect 16811 16612 16856 16640
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 16960 16649 16988 16748
rect 22066 16708 22094 16748
rect 22738 16736 22744 16788
rect 22796 16776 22802 16788
rect 24394 16776 24400 16788
rect 22796 16748 24400 16776
rect 22796 16736 22802 16748
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 24486 16736 24492 16788
rect 24544 16776 24550 16788
rect 24581 16779 24639 16785
rect 24581 16776 24593 16779
rect 24544 16748 24593 16776
rect 24544 16736 24550 16748
rect 24581 16745 24593 16748
rect 24627 16776 24639 16779
rect 25133 16779 25191 16785
rect 25133 16776 25145 16779
rect 24627 16748 25145 16776
rect 24627 16745 24639 16748
rect 24581 16739 24639 16745
rect 25133 16745 25145 16748
rect 25179 16776 25191 16779
rect 25682 16776 25688 16788
rect 25179 16748 25688 16776
rect 25179 16745 25191 16748
rect 25133 16739 25191 16745
rect 25682 16736 25688 16748
rect 25740 16736 25746 16788
rect 25774 16736 25780 16788
rect 25832 16776 25838 16788
rect 28994 16776 29000 16788
rect 25832 16748 28580 16776
rect 28955 16748 29000 16776
rect 25832 16736 25838 16748
rect 27522 16708 27528 16720
rect 22066 16680 27528 16708
rect 27522 16668 27528 16680
rect 27580 16668 27586 16720
rect 28442 16708 28448 16720
rect 28403 16680 28448 16708
rect 28442 16668 28448 16680
rect 28500 16668 28506 16720
rect 28552 16708 28580 16748
rect 28994 16736 29000 16748
rect 29052 16736 29058 16788
rect 31665 16779 31723 16785
rect 31665 16776 31677 16779
rect 29104 16748 31677 16776
rect 29104 16708 29132 16748
rect 31665 16745 31677 16748
rect 31711 16745 31723 16779
rect 31665 16739 31723 16745
rect 31938 16736 31944 16788
rect 31996 16776 32002 16788
rect 37366 16776 37372 16788
rect 31996 16748 37372 16776
rect 31996 16736 32002 16748
rect 37366 16736 37372 16748
rect 37424 16776 37430 16788
rect 38194 16776 38200 16788
rect 37424 16748 38200 16776
rect 37424 16736 37430 16748
rect 38194 16736 38200 16748
rect 38252 16736 38258 16788
rect 44082 16736 44088 16788
rect 44140 16776 44146 16788
rect 46109 16779 46167 16785
rect 46109 16776 46121 16779
rect 44140 16748 46121 16776
rect 44140 16736 44146 16748
rect 46109 16745 46121 16748
rect 46155 16776 46167 16779
rect 46658 16776 46664 16788
rect 46155 16748 46664 16776
rect 46155 16745 46167 16748
rect 46109 16739 46167 16745
rect 28552 16680 29132 16708
rect 29270 16668 29276 16720
rect 29328 16708 29334 16720
rect 36446 16708 36452 16720
rect 29328 16680 36452 16708
rect 29328 16668 29334 16680
rect 36446 16668 36452 16680
rect 36504 16668 36510 16720
rect 40681 16711 40739 16717
rect 40681 16677 40693 16711
rect 40727 16708 40739 16711
rect 40727 16680 41276 16708
rect 40727 16677 40739 16680
rect 40681 16671 40739 16677
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16609 17003 16643
rect 17126 16640 17132 16652
rect 17087 16612 17132 16640
rect 16945 16603 17003 16609
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 17494 16600 17500 16652
rect 17552 16640 17558 16652
rect 17681 16643 17739 16649
rect 17681 16640 17693 16643
rect 17552 16612 17693 16640
rect 17552 16600 17558 16612
rect 17681 16609 17693 16612
rect 17727 16609 17739 16643
rect 17681 16603 17739 16609
rect 17957 16643 18015 16649
rect 17957 16609 17969 16643
rect 18003 16640 18015 16643
rect 18138 16640 18144 16652
rect 18003 16612 18144 16640
rect 18003 16609 18015 16612
rect 17957 16603 18015 16609
rect 18138 16600 18144 16612
rect 18196 16640 18202 16652
rect 18414 16640 18420 16652
rect 18196 16612 18420 16640
rect 18196 16600 18202 16612
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 20162 16600 20168 16652
rect 20220 16640 20226 16652
rect 20257 16643 20315 16649
rect 20257 16640 20269 16643
rect 20220 16612 20269 16640
rect 20220 16600 20226 16612
rect 20257 16609 20269 16612
rect 20303 16609 20315 16643
rect 20257 16603 20315 16609
rect 23014 16600 23020 16652
rect 23072 16640 23078 16652
rect 23072 16612 29132 16640
rect 23072 16600 23078 16612
rect 6546 16532 6552 16584
rect 6604 16572 6610 16584
rect 6917 16575 6975 16581
rect 6917 16572 6929 16575
rect 6604 16544 6929 16572
rect 6604 16532 6610 16544
rect 6917 16541 6929 16544
rect 6963 16541 6975 16575
rect 10962 16572 10968 16584
rect 10923 16544 10968 16572
rect 6917 16535 6975 16541
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 17034 16572 17040 16584
rect 12268 16544 16896 16572
rect 16995 16544 17040 16572
rect 1848 16507 1906 16513
rect 1848 16473 1860 16507
rect 1894 16504 1906 16507
rect 2314 16504 2320 16516
rect 1894 16476 2320 16504
rect 1894 16473 1906 16476
rect 1848 16467 1906 16473
rect 2314 16464 2320 16476
rect 2372 16464 2378 16516
rect 2406 16464 2412 16516
rect 2464 16504 2470 16516
rect 12268 16504 12296 16544
rect 12434 16513 12440 16516
rect 2464 16476 12296 16504
rect 2464 16464 2470 16476
rect 12428 16467 12440 16513
rect 12492 16504 12498 16516
rect 14185 16507 14243 16513
rect 14185 16504 14197 16507
rect 12492 16476 12528 16504
rect 13556 16476 14197 16504
rect 12434 16464 12440 16467
rect 12492 16464 12498 16476
rect 1394 16396 1400 16448
rect 1452 16436 1458 16448
rect 2682 16436 2688 16448
rect 1452 16408 2688 16436
rect 1452 16396 1458 16408
rect 2682 16396 2688 16408
rect 2740 16436 2746 16448
rect 2961 16439 3019 16445
rect 2961 16436 2973 16439
rect 2740 16408 2973 16436
rect 2740 16396 2746 16408
rect 2961 16405 2973 16408
rect 3007 16405 3019 16439
rect 2961 16399 3019 16405
rect 6733 16439 6791 16445
rect 6733 16405 6745 16439
rect 6779 16436 6791 16439
rect 6822 16436 6828 16448
rect 6779 16408 6828 16436
rect 6779 16405 6791 16408
rect 6733 16399 6791 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 13556 16445 13584 16476
rect 14185 16473 14197 16476
rect 14231 16504 14243 16507
rect 15010 16504 15016 16516
rect 14231 16476 15016 16504
rect 14231 16473 14243 16476
rect 14185 16467 14243 16473
rect 15010 16464 15016 16476
rect 15068 16464 15074 16516
rect 15194 16504 15200 16516
rect 15155 16476 15200 16504
rect 15194 16464 15200 16476
rect 15252 16464 15258 16516
rect 15378 16464 15384 16516
rect 15436 16504 15442 16516
rect 15746 16504 15752 16516
rect 15436 16476 15752 16504
rect 15436 16464 15442 16476
rect 15746 16464 15752 16476
rect 15804 16464 15810 16516
rect 15930 16464 15936 16516
rect 15988 16504 15994 16516
rect 16868 16504 16896 16544
rect 17034 16532 17040 16544
rect 17092 16532 17098 16584
rect 23106 16572 23112 16584
rect 17144 16544 23112 16572
rect 17144 16504 17172 16544
rect 23106 16532 23112 16544
rect 23164 16532 23170 16584
rect 24627 16541 24685 16547
rect 15988 16476 16804 16504
rect 16868 16476 17172 16504
rect 20524 16507 20582 16513
rect 15988 16464 15994 16476
rect 11057 16439 11115 16445
rect 11057 16436 11069 16439
rect 10928 16408 11069 16436
rect 10928 16396 10934 16408
rect 11057 16405 11069 16408
rect 11103 16405 11115 16439
rect 11057 16399 11115 16405
rect 13541 16439 13599 16445
rect 13541 16405 13553 16439
rect 13587 16405 13599 16439
rect 14366 16436 14372 16448
rect 14327 16408 14372 16436
rect 13541 16399 13599 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 14550 16436 14556 16448
rect 14511 16408 14556 16436
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 15212 16436 15240 16464
rect 16298 16436 16304 16448
rect 15212 16408 16304 16436
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16666 16436 16672 16448
rect 16627 16408 16672 16436
rect 16666 16396 16672 16408
rect 16724 16396 16730 16448
rect 16776 16436 16804 16476
rect 20524 16473 20536 16507
rect 20570 16504 20582 16507
rect 21818 16504 21824 16516
rect 20570 16476 21824 16504
rect 20570 16473 20582 16476
rect 20524 16467 20582 16473
rect 21818 16464 21824 16476
rect 21876 16464 21882 16516
rect 23474 16464 23480 16516
rect 23532 16504 23538 16516
rect 24397 16507 24455 16513
rect 24397 16504 24409 16507
rect 23532 16476 24409 16504
rect 23532 16464 23538 16476
rect 24397 16473 24409 16476
rect 24443 16473 24455 16507
rect 24627 16507 24639 16541
rect 24673 16538 24685 16541
rect 24673 16516 24716 16538
rect 24762 16532 24768 16584
rect 24820 16532 24826 16584
rect 28074 16532 28080 16584
rect 28132 16572 28138 16584
rect 28721 16575 28779 16581
rect 28721 16572 28733 16575
rect 28132 16544 28733 16572
rect 28132 16532 28138 16544
rect 28721 16541 28733 16544
rect 28767 16541 28779 16575
rect 28721 16535 28779 16541
rect 28813 16575 28871 16581
rect 28813 16541 28825 16575
rect 28859 16572 28871 16575
rect 28994 16572 29000 16584
rect 28859 16544 29000 16572
rect 28859 16541 28871 16544
rect 28813 16535 28871 16541
rect 28994 16532 29000 16544
rect 29052 16532 29058 16584
rect 29104 16572 29132 16612
rect 29638 16600 29644 16652
rect 29696 16640 29702 16652
rect 29696 16612 30052 16640
rect 29696 16600 29702 16612
rect 29730 16572 29736 16584
rect 29104 16544 29736 16572
rect 29730 16532 29736 16544
rect 29788 16532 29794 16584
rect 30024 16581 30052 16612
rect 35526 16600 35532 16652
rect 35584 16640 35590 16652
rect 37550 16640 37556 16652
rect 35584 16612 36492 16640
rect 37511 16612 37556 16640
rect 35584 16600 35590 16612
rect 30009 16575 30067 16581
rect 30009 16541 30021 16575
rect 30055 16572 30067 16575
rect 31021 16575 31079 16581
rect 31021 16572 31033 16575
rect 30055 16544 31033 16572
rect 30055 16541 30067 16544
rect 30009 16535 30067 16541
rect 31021 16541 31033 16544
rect 31067 16541 31079 16575
rect 31021 16535 31079 16541
rect 31169 16575 31227 16581
rect 31169 16541 31181 16575
rect 31215 16572 31227 16575
rect 31215 16541 31248 16572
rect 31169 16535 31248 16541
rect 24673 16507 24676 16516
rect 24627 16501 24676 16507
rect 24397 16467 24455 16473
rect 24670 16464 24676 16501
rect 24728 16464 24734 16516
rect 18230 16436 18236 16448
rect 16776 16408 18236 16436
rect 18230 16396 18236 16408
rect 18288 16396 18294 16448
rect 20622 16396 20628 16448
rect 20680 16436 20686 16448
rect 21637 16439 21695 16445
rect 21637 16436 21649 16439
rect 20680 16408 21649 16436
rect 20680 16396 20686 16408
rect 21637 16405 21649 16408
rect 21683 16436 21695 16439
rect 22186 16436 22192 16448
rect 21683 16408 22192 16436
rect 21683 16405 21695 16408
rect 21637 16399 21695 16405
rect 22186 16396 22192 16408
rect 22244 16396 22250 16448
rect 24780 16445 24808 16532
rect 25682 16504 25688 16516
rect 25643 16476 25688 16504
rect 25682 16464 25688 16476
rect 25740 16504 25746 16516
rect 25740 16476 28488 16504
rect 25740 16464 25746 16476
rect 24765 16439 24823 16445
rect 24765 16405 24777 16439
rect 24811 16405 24823 16439
rect 25774 16436 25780 16448
rect 25735 16408 25780 16436
rect 24765 16399 24823 16405
rect 25774 16396 25780 16408
rect 25832 16396 25838 16448
rect 28460 16436 28488 16476
rect 28534 16464 28540 16516
rect 28592 16504 28598 16516
rect 28629 16507 28687 16513
rect 28629 16504 28641 16507
rect 28592 16476 28641 16504
rect 28592 16464 28598 16476
rect 28629 16473 28641 16476
rect 28675 16504 28687 16507
rect 31220 16504 31248 16535
rect 31294 16532 31300 16584
rect 31352 16572 31358 16584
rect 31478 16572 31484 16584
rect 31536 16581 31542 16584
rect 31352 16544 31397 16572
rect 31444 16544 31484 16572
rect 31352 16532 31358 16544
rect 31478 16532 31484 16544
rect 31536 16535 31544 16581
rect 31536 16532 31542 16535
rect 34790 16532 34796 16584
rect 34848 16572 34854 16584
rect 35161 16575 35219 16581
rect 35161 16572 35173 16575
rect 34848 16544 35173 16572
rect 34848 16532 34854 16544
rect 35161 16541 35173 16544
rect 35207 16541 35219 16575
rect 35161 16535 35219 16541
rect 35253 16575 35311 16581
rect 35253 16541 35265 16575
rect 35299 16572 35311 16575
rect 36035 16575 36093 16581
rect 36035 16572 36047 16575
rect 35299 16544 36047 16572
rect 35299 16541 35311 16544
rect 35253 16535 35311 16541
rect 36035 16541 36047 16544
rect 36081 16541 36093 16575
rect 36167 16572 36173 16584
rect 36128 16544 36173 16572
rect 36035 16535 36093 16541
rect 36167 16532 36173 16544
rect 36225 16532 36231 16584
rect 36262 16532 36268 16584
rect 36320 16569 36326 16584
rect 36464 16581 36492 16612
rect 37550 16600 37556 16612
rect 37608 16600 37614 16652
rect 40788 16612 41000 16640
rect 36449 16575 36507 16581
rect 36320 16541 36362 16569
rect 36449 16541 36461 16575
rect 36495 16541 36507 16575
rect 37090 16572 37096 16584
rect 37051 16544 37096 16572
rect 36320 16532 36326 16541
rect 36449 16535 36507 16541
rect 37090 16532 37096 16544
rect 37148 16532 37154 16584
rect 38746 16532 38752 16584
rect 38804 16572 38810 16584
rect 40788 16572 40816 16612
rect 38804 16544 40816 16572
rect 40865 16575 40923 16581
rect 38804 16532 38810 16544
rect 40865 16541 40877 16575
rect 40911 16541 40923 16575
rect 40972 16572 41000 16612
rect 41141 16575 41199 16581
rect 41141 16572 41153 16575
rect 40972 16544 41153 16572
rect 40865 16535 40923 16541
rect 41141 16541 41153 16544
rect 41187 16541 41199 16575
rect 41141 16535 41199 16541
rect 31386 16504 31392 16516
rect 28675 16476 31248 16504
rect 31347 16476 31392 16504
rect 28675 16473 28687 16476
rect 28629 16467 28687 16473
rect 29454 16436 29460 16448
rect 28460 16408 29460 16436
rect 29454 16396 29460 16408
rect 29512 16396 29518 16448
rect 31220 16436 31248 16476
rect 31386 16464 31392 16476
rect 31444 16464 31450 16516
rect 37798 16507 37856 16513
rect 37798 16504 37810 16507
rect 36924 16476 37810 16504
rect 32766 16436 32772 16448
rect 31220 16408 32772 16436
rect 32766 16396 32772 16408
rect 32824 16396 32830 16448
rect 35802 16436 35808 16448
rect 35763 16408 35808 16436
rect 35802 16396 35808 16408
rect 35860 16396 35866 16448
rect 36924 16445 36952 16476
rect 37798 16473 37810 16476
rect 37844 16473 37856 16507
rect 37798 16467 37856 16473
rect 36909 16439 36967 16445
rect 36909 16405 36921 16439
rect 36955 16405 36967 16439
rect 36909 16399 36967 16405
rect 36998 16396 37004 16448
rect 37056 16436 37062 16448
rect 38933 16439 38991 16445
rect 38933 16436 38945 16439
rect 37056 16408 38945 16436
rect 37056 16396 37062 16408
rect 38933 16405 38945 16408
rect 38979 16405 38991 16439
rect 40880 16436 40908 16535
rect 41248 16504 41276 16680
rect 42886 16668 42892 16720
rect 42944 16708 42950 16720
rect 46584 16717 46612 16748
rect 46658 16736 46664 16748
rect 46716 16736 46722 16788
rect 46934 16776 46940 16788
rect 46895 16748 46940 16776
rect 46934 16736 46940 16748
rect 46992 16736 46998 16788
rect 53374 16776 53380 16788
rect 47872 16748 53380 16776
rect 45097 16711 45155 16717
rect 45097 16708 45109 16711
rect 42944 16680 45109 16708
rect 42944 16668 42950 16680
rect 45097 16677 45109 16680
rect 45143 16677 45155 16711
rect 45097 16671 45155 16677
rect 46569 16711 46627 16717
rect 46569 16677 46581 16711
rect 46615 16677 46627 16711
rect 46569 16671 46627 16677
rect 42518 16640 42524 16652
rect 41892 16612 42380 16640
rect 42479 16612 42524 16640
rect 41325 16575 41383 16581
rect 41325 16541 41337 16575
rect 41371 16572 41383 16575
rect 41690 16572 41696 16584
rect 41371 16544 41696 16572
rect 41371 16541 41383 16544
rect 41325 16535 41383 16541
rect 41690 16532 41696 16544
rect 41748 16532 41754 16584
rect 41785 16575 41843 16581
rect 41785 16541 41797 16575
rect 41831 16541 41843 16575
rect 41785 16535 41843 16541
rect 41800 16504 41828 16535
rect 41248 16476 41828 16504
rect 41892 16436 41920 16612
rect 41969 16575 42027 16581
rect 41969 16541 41981 16575
rect 42015 16541 42027 16575
rect 42242 16572 42248 16584
rect 42203 16544 42248 16572
rect 41969 16535 42027 16541
rect 41984 16504 42012 16535
rect 42242 16532 42248 16544
rect 42300 16532 42306 16584
rect 42352 16572 42380 16612
rect 42518 16600 42524 16612
rect 42576 16600 42582 16652
rect 47578 16600 47584 16652
rect 47636 16640 47642 16652
rect 47872 16649 47900 16748
rect 50816 16652 50844 16748
rect 53374 16736 53380 16748
rect 53432 16736 53438 16788
rect 47857 16643 47915 16649
rect 47857 16640 47869 16643
rect 47636 16612 47869 16640
rect 47636 16600 47642 16612
rect 47857 16609 47869 16612
rect 47903 16609 47915 16643
rect 50798 16640 50804 16652
rect 50711 16612 50804 16640
rect 47857 16603 47915 16609
rect 50798 16600 50804 16612
rect 50856 16600 50862 16652
rect 53392 16649 53420 16736
rect 53377 16643 53435 16649
rect 53377 16609 53389 16643
rect 53423 16609 53435 16643
rect 53377 16603 53435 16609
rect 42613 16575 42671 16581
rect 42613 16572 42625 16575
rect 42352 16544 42625 16572
rect 42613 16541 42625 16544
rect 42659 16572 42671 16575
rect 44358 16572 44364 16584
rect 42659 16544 44364 16572
rect 42659 16541 42671 16544
rect 42613 16535 42671 16541
rect 44358 16532 44364 16544
rect 44416 16532 44422 16584
rect 45278 16572 45284 16584
rect 45239 16544 45284 16572
rect 45278 16532 45284 16544
rect 45336 16532 45342 16584
rect 45830 16572 45836 16584
rect 45791 16544 45836 16572
rect 45830 16532 45836 16544
rect 45888 16532 45894 16584
rect 45922 16532 45928 16584
rect 45980 16572 45986 16584
rect 51074 16581 51080 16584
rect 45980 16544 46025 16572
rect 45980 16532 45986 16544
rect 51068 16535 51080 16581
rect 51132 16572 51138 16584
rect 51132 16544 51168 16572
rect 51074 16532 51080 16535
rect 51132 16532 51138 16544
rect 42886 16504 42892 16516
rect 41984 16476 42892 16504
rect 42886 16464 42892 16476
rect 42944 16464 42950 16516
rect 45002 16504 45008 16516
rect 44963 16476 45008 16504
rect 45002 16464 45008 16476
rect 45060 16464 45066 16516
rect 45189 16507 45247 16513
rect 45189 16473 45201 16507
rect 45235 16504 45247 16507
rect 45848 16504 45876 16532
rect 45235 16476 45876 16504
rect 45235 16473 45247 16476
rect 45189 16467 45247 16473
rect 47670 16464 47676 16516
rect 47728 16504 47734 16516
rect 48102 16507 48160 16513
rect 48102 16504 48114 16507
rect 47728 16476 48114 16504
rect 47728 16464 47734 16476
rect 48102 16473 48114 16476
rect 48148 16473 48160 16507
rect 48102 16467 48160 16473
rect 53190 16464 53196 16516
rect 53248 16504 53254 16516
rect 53622 16507 53680 16513
rect 53622 16504 53634 16507
rect 53248 16476 53634 16504
rect 53248 16464 53254 16476
rect 53622 16473 53634 16476
rect 53668 16473 53680 16507
rect 53622 16467 53680 16473
rect 40880 16408 41920 16436
rect 38933 16399 38991 16405
rect 42518 16396 42524 16448
rect 42576 16436 42582 16448
rect 42797 16439 42855 16445
rect 42797 16436 42809 16439
rect 42576 16408 42809 16436
rect 42576 16396 42582 16408
rect 42797 16405 42809 16408
rect 42843 16405 42855 16439
rect 42797 16399 42855 16405
rect 46750 16396 46756 16448
rect 46808 16436 46814 16448
rect 46937 16439 46995 16445
rect 46937 16436 46949 16439
rect 46808 16408 46949 16436
rect 46808 16396 46814 16408
rect 46937 16405 46949 16408
rect 46983 16405 46995 16439
rect 46937 16399 46995 16405
rect 47121 16439 47179 16445
rect 47121 16405 47133 16439
rect 47167 16436 47179 16439
rect 47854 16436 47860 16448
rect 47167 16408 47860 16436
rect 47167 16405 47179 16408
rect 47121 16399 47179 16405
rect 47854 16396 47860 16408
rect 47912 16396 47918 16448
rect 49234 16436 49240 16448
rect 49195 16408 49240 16436
rect 49234 16396 49240 16408
rect 49292 16396 49298 16448
rect 52181 16439 52239 16445
rect 52181 16405 52193 16439
rect 52227 16436 52239 16439
rect 52454 16436 52460 16448
rect 52227 16408 52460 16436
rect 52227 16405 52239 16408
rect 52181 16399 52239 16405
rect 52454 16396 52460 16408
rect 52512 16396 52518 16448
rect 53834 16396 53840 16448
rect 53892 16436 53898 16448
rect 54757 16439 54815 16445
rect 54757 16436 54769 16439
rect 53892 16408 54769 16436
rect 53892 16396 53898 16408
rect 54757 16405 54769 16408
rect 54803 16405 54815 16439
rect 54757 16399 54815 16405
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 2314 16232 2320 16244
rect 2275 16204 2320 16232
rect 2314 16192 2320 16204
rect 2372 16192 2378 16244
rect 2682 16232 2688 16244
rect 2643 16204 2688 16232
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 12345 16235 12403 16241
rect 12345 16201 12357 16235
rect 12391 16232 12403 16235
rect 12434 16232 12440 16244
rect 12391 16204 12440 16232
rect 12391 16201 12403 16204
rect 12345 16195 12403 16201
rect 12434 16192 12440 16204
rect 12492 16192 12498 16244
rect 17954 16232 17960 16244
rect 17915 16204 17960 16232
rect 17954 16192 17960 16204
rect 18012 16192 18018 16244
rect 21818 16232 21824 16244
rect 21779 16204 21824 16232
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 22186 16232 22192 16244
rect 22147 16204 22192 16232
rect 22186 16192 22192 16204
rect 22244 16192 22250 16244
rect 28166 16232 28172 16244
rect 28127 16204 28172 16232
rect 28166 16192 28172 16204
rect 28224 16192 28230 16244
rect 28994 16232 29000 16244
rect 28368 16204 29000 16232
rect 1857 16167 1915 16173
rect 1857 16133 1869 16167
rect 1903 16164 1915 16167
rect 2406 16164 2412 16176
rect 1903 16136 2412 16164
rect 1903 16133 1915 16136
rect 1857 16127 1915 16133
rect 2406 16124 2412 16136
rect 2464 16124 2470 16176
rect 2590 16124 2596 16176
rect 2648 16164 2654 16176
rect 14458 16164 14464 16176
rect 2648 16136 14464 16164
rect 2648 16124 2654 16136
rect 14458 16124 14464 16136
rect 14516 16124 14522 16176
rect 14550 16124 14556 16176
rect 14608 16164 14614 16176
rect 25682 16164 25688 16176
rect 14608 16136 25688 16164
rect 14608 16124 14614 16136
rect 25682 16124 25688 16136
rect 25740 16124 25746 16176
rect 1486 16096 1492 16108
rect 1447 16068 1492 16096
rect 1486 16056 1492 16068
rect 1544 16056 1550 16108
rect 2498 16096 2504 16108
rect 2459 16068 2504 16096
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 2774 16056 2780 16108
rect 2832 16096 2838 16108
rect 4525 16099 4583 16105
rect 2832 16068 2877 16096
rect 2832 16056 2838 16068
rect 4525 16065 4537 16099
rect 4571 16096 4583 16099
rect 4614 16096 4620 16108
rect 4571 16068 4620 16096
rect 4571 16065 4583 16068
rect 4525 16059 4583 16065
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 6822 16056 6828 16108
rect 6880 16096 6886 16108
rect 6989 16099 7047 16105
rect 6989 16096 7001 16099
rect 6880 16068 7001 16096
rect 6880 16056 6886 16068
rect 6989 16065 7001 16068
rect 7035 16065 7047 16099
rect 6989 16059 7047 16065
rect 8938 16056 8944 16108
rect 8996 16096 9002 16108
rect 9490 16096 9496 16108
rect 8996 16068 9496 16096
rect 8996 16056 9002 16068
rect 9490 16056 9496 16068
rect 9548 16096 9554 16108
rect 9585 16099 9643 16105
rect 9585 16096 9597 16099
rect 9548 16068 9597 16096
rect 9548 16056 9554 16068
rect 9585 16065 9597 16068
rect 9631 16065 9643 16099
rect 9585 16059 9643 16065
rect 9852 16099 9910 16105
rect 9852 16065 9864 16099
rect 9898 16096 9910 16099
rect 10594 16096 10600 16108
rect 9898 16068 10600 16096
rect 9898 16065 9910 16068
rect 9852 16059 9910 16065
rect 10594 16056 10600 16068
rect 10652 16056 10658 16108
rect 10962 16056 10968 16108
rect 11020 16096 11026 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11020 16068 11713 16096
rect 11020 16056 11026 16068
rect 11701 16065 11713 16068
rect 11747 16096 11759 16099
rect 11882 16096 11888 16108
rect 11747 16068 11888 16096
rect 11747 16065 11759 16068
rect 11701 16059 11759 16065
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 12526 16096 12532 16108
rect 12487 16068 12532 16096
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16390 16096 16396 16108
rect 15979 16068 16396 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16096 17003 16099
rect 17862 16096 17868 16108
rect 16991 16068 17868 16096
rect 16991 16065 17003 16068
rect 16945 16059 17003 16065
rect 17862 16056 17868 16068
rect 17920 16096 17926 16108
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 17920 16068 18153 16096
rect 17920 16056 17926 16068
rect 18141 16065 18153 16068
rect 18187 16065 18199 16099
rect 18141 16059 18199 16065
rect 18230 16056 18236 16108
rect 18288 16096 18294 16108
rect 18288 16068 18333 16096
rect 18288 16056 18294 16068
rect 18414 16056 18420 16108
rect 18472 16096 18478 16108
rect 22005 16099 22063 16105
rect 18472 16068 18517 16096
rect 18472 16056 18478 16068
rect 22005 16065 22017 16099
rect 22051 16096 22063 16099
rect 22186 16096 22192 16108
rect 22051 16068 22192 16096
rect 22051 16065 22063 16068
rect 22005 16059 22063 16065
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 22281 16099 22339 16105
rect 22281 16065 22293 16099
rect 22327 16096 22339 16099
rect 22370 16096 22376 16108
rect 22327 16068 22376 16096
rect 22327 16065 22339 16068
rect 22281 16059 22339 16065
rect 22370 16056 22376 16068
rect 22428 16096 22434 16108
rect 23014 16096 23020 16108
rect 22428 16068 23020 16096
rect 22428 16056 22434 16068
rect 23014 16056 23020 16068
rect 23072 16056 23078 16108
rect 23198 16096 23204 16108
rect 23159 16068 23204 16096
rect 23198 16056 23204 16068
rect 23256 16056 23262 16108
rect 23468 16099 23526 16105
rect 23468 16065 23480 16099
rect 23514 16096 23526 16099
rect 24394 16096 24400 16108
rect 23514 16068 24400 16096
rect 23514 16065 23526 16068
rect 23468 16059 23526 16065
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 28368 16105 28396 16204
rect 28994 16192 29000 16204
rect 29052 16192 29058 16244
rect 36722 16232 36728 16244
rect 36683 16204 36728 16232
rect 36722 16192 36728 16204
rect 36780 16192 36786 16244
rect 40589 16235 40647 16241
rect 40589 16201 40601 16235
rect 40635 16232 40647 16235
rect 42610 16232 42616 16244
rect 40635 16204 42616 16232
rect 40635 16201 40647 16204
rect 40589 16195 40647 16201
rect 42610 16192 42616 16204
rect 42668 16192 42674 16244
rect 46750 16232 46756 16244
rect 46711 16204 46756 16232
rect 46750 16192 46756 16204
rect 46808 16192 46814 16244
rect 47670 16232 47676 16244
rect 47631 16204 47676 16232
rect 47670 16192 47676 16204
rect 47728 16192 47734 16244
rect 51442 16192 51448 16244
rect 51500 16232 51506 16244
rect 51721 16235 51779 16241
rect 51721 16232 51733 16235
rect 51500 16204 51733 16232
rect 51500 16192 51506 16204
rect 51721 16201 51733 16204
rect 51767 16201 51779 16235
rect 51721 16195 51779 16201
rect 28442 16124 28448 16176
rect 28500 16164 28506 16176
rect 30009 16167 30067 16173
rect 28500 16136 28672 16164
rect 28500 16124 28506 16136
rect 28353 16099 28411 16105
rect 28353 16065 28365 16099
rect 28399 16065 28411 16099
rect 28534 16096 28540 16108
rect 28495 16068 28540 16096
rect 28353 16059 28411 16065
rect 28534 16056 28540 16068
rect 28592 16056 28598 16108
rect 28644 16105 28672 16136
rect 30009 16133 30021 16167
rect 30055 16164 30067 16167
rect 30282 16164 30288 16176
rect 30055 16136 30288 16164
rect 30055 16133 30067 16136
rect 30009 16127 30067 16133
rect 30282 16124 30288 16136
rect 30340 16124 30346 16176
rect 32950 16164 32956 16176
rect 32600 16136 32956 16164
rect 28629 16099 28687 16105
rect 28629 16065 28641 16099
rect 28675 16065 28687 16099
rect 28629 16059 28687 16065
rect 29086 16056 29092 16108
rect 29144 16096 29150 16108
rect 29638 16096 29644 16108
rect 29144 16068 29644 16096
rect 29144 16056 29150 16068
rect 29638 16056 29644 16068
rect 29696 16056 29702 16108
rect 29822 16105 29828 16108
rect 29789 16099 29828 16105
rect 29789 16065 29801 16099
rect 29789 16059 29828 16065
rect 29822 16056 29828 16059
rect 29880 16056 29886 16108
rect 29917 16099 29975 16105
rect 29917 16065 29929 16099
rect 29963 16065 29975 16099
rect 29917 16059 29975 16065
rect 3786 15988 3792 16040
rect 3844 16028 3850 16040
rect 6733 16031 6791 16037
rect 6733 16028 6745 16031
rect 3844 16000 6745 16028
rect 3844 15988 3850 16000
rect 6733 15997 6745 16000
rect 6779 15997 6791 16031
rect 11517 16031 11575 16037
rect 11517 16028 11529 16031
rect 6733 15991 6791 15997
rect 10980 16000 11529 16028
rect 4341 15895 4399 15901
rect 4341 15861 4353 15895
rect 4387 15892 4399 15895
rect 4706 15892 4712 15904
rect 4387 15864 4712 15892
rect 4387 15861 4399 15864
rect 4341 15855 4399 15861
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 6748 15892 6776 15991
rect 10980 15904 11008 16000
rect 11517 15997 11529 16000
rect 11563 15997 11575 16031
rect 11517 15991 11575 15997
rect 16574 15988 16580 16040
rect 16632 16028 16638 16040
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 16632 16000 16681 16028
rect 16632 15988 16638 16000
rect 16669 15997 16681 16000
rect 16715 15997 16727 16031
rect 16669 15991 16727 15997
rect 18325 16031 18383 16037
rect 18325 15997 18337 16031
rect 18371 15997 18383 16031
rect 18325 15991 18383 15997
rect 6914 15892 6920 15904
rect 6748 15864 6920 15892
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 8110 15892 8116 15904
rect 8071 15864 8116 15892
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 10962 15892 10968 15904
rect 10923 15864 10968 15892
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11885 15895 11943 15901
rect 11885 15892 11897 15895
rect 11112 15864 11897 15892
rect 11112 15852 11118 15864
rect 11885 15861 11897 15864
rect 11931 15861 11943 15895
rect 16022 15892 16028 15904
rect 15983 15864 16028 15892
rect 11885 15855 11943 15861
rect 16022 15852 16028 15864
rect 16080 15852 16086 15904
rect 18340 15892 18368 15991
rect 28166 15988 28172 16040
rect 28224 16028 28230 16040
rect 28445 16031 28503 16037
rect 28445 16028 28457 16031
rect 28224 16000 28457 16028
rect 28224 15988 28230 16000
rect 28445 15997 28457 16000
rect 28491 15997 28503 16031
rect 28445 15991 28503 15997
rect 28718 15988 28724 16040
rect 28776 16028 28782 16040
rect 29932 16028 29960 16059
rect 30098 16056 30104 16108
rect 30156 16105 30162 16108
rect 32600 16105 32628 16136
rect 32950 16124 32956 16136
rect 33008 16164 33014 16176
rect 35612 16167 35670 16173
rect 33008 16136 35388 16164
rect 33008 16124 33014 16136
rect 32858 16105 32864 16108
rect 30156 16096 30164 16105
rect 32585 16099 32643 16105
rect 30156 16068 30201 16096
rect 30156 16059 30164 16068
rect 32585 16065 32597 16099
rect 32631 16065 32643 16099
rect 32585 16059 32643 16065
rect 32852 16059 32864 16105
rect 32916 16096 32922 16108
rect 35360 16105 35388 16136
rect 35612 16133 35624 16167
rect 35658 16164 35670 16167
rect 35802 16164 35808 16176
rect 35658 16136 35808 16164
rect 35658 16133 35670 16136
rect 35612 16127 35670 16133
rect 35802 16124 35808 16136
rect 35860 16124 35866 16176
rect 45830 16124 45836 16176
rect 45888 16164 45894 16176
rect 46569 16167 46627 16173
rect 46569 16164 46581 16167
rect 45888 16136 46581 16164
rect 45888 16124 45894 16136
rect 46569 16133 46581 16136
rect 46615 16164 46627 16167
rect 49234 16164 49240 16176
rect 46615 16136 49240 16164
rect 46615 16133 46627 16136
rect 46569 16127 46627 16133
rect 49234 16124 49240 16136
rect 49292 16124 49298 16176
rect 51074 16124 51080 16176
rect 51132 16164 51138 16176
rect 51353 16167 51411 16173
rect 51353 16164 51365 16167
rect 51132 16136 51365 16164
rect 51132 16124 51138 16136
rect 51353 16133 51365 16136
rect 51399 16133 51411 16167
rect 51353 16127 51411 16133
rect 51569 16167 51627 16173
rect 51569 16133 51581 16167
rect 51615 16164 51627 16167
rect 52914 16164 52920 16176
rect 51615 16136 52920 16164
rect 51615 16133 51627 16136
rect 51569 16127 51627 16133
rect 52914 16124 52920 16136
rect 52972 16124 52978 16176
rect 53193 16167 53251 16173
rect 53193 16133 53205 16167
rect 53239 16164 53251 16167
rect 54205 16167 54263 16173
rect 54205 16164 54217 16167
rect 53239 16136 54217 16164
rect 53239 16133 53251 16136
rect 53193 16127 53251 16133
rect 54205 16133 54217 16136
rect 54251 16133 54263 16167
rect 54205 16127 54263 16133
rect 35345 16099 35403 16105
rect 32916 16068 32952 16096
rect 30156 16056 30162 16059
rect 32858 16056 32864 16059
rect 32916 16056 32922 16068
rect 35345 16065 35357 16099
rect 35391 16096 35403 16099
rect 37550 16096 37556 16108
rect 35391 16068 37556 16096
rect 35391 16065 35403 16068
rect 35345 16059 35403 16065
rect 37550 16056 37556 16068
rect 37608 16056 37614 16108
rect 40310 16096 40316 16108
rect 40271 16068 40316 16096
rect 40310 16056 40316 16068
rect 40368 16056 40374 16108
rect 40402 16056 40408 16108
rect 40460 16096 40466 16108
rect 43622 16096 43628 16108
rect 40460 16068 40505 16096
rect 43535 16068 43628 16096
rect 40460 16056 40466 16068
rect 43622 16056 43628 16068
rect 43680 16096 43686 16108
rect 45002 16096 45008 16108
rect 43680 16068 45008 16096
rect 43680 16056 43686 16068
rect 45002 16056 45008 16068
rect 45060 16056 45066 16108
rect 45922 16056 45928 16108
rect 45980 16096 45986 16108
rect 46385 16099 46443 16105
rect 46385 16096 46397 16099
rect 45980 16068 46397 16096
rect 45980 16056 45986 16068
rect 46385 16065 46397 16068
rect 46431 16065 46443 16099
rect 47854 16096 47860 16108
rect 47815 16068 47860 16096
rect 46385 16059 46443 16065
rect 47854 16056 47860 16068
rect 47912 16056 47918 16108
rect 53282 16056 53288 16108
rect 53340 16096 53346 16108
rect 53377 16099 53435 16105
rect 53377 16096 53389 16099
rect 53340 16068 53389 16096
rect 53340 16056 53346 16068
rect 53377 16065 53389 16068
rect 53423 16065 53435 16099
rect 53377 16059 53435 16065
rect 31294 16028 31300 16040
rect 28776 16000 31300 16028
rect 28776 15988 28782 16000
rect 31294 15988 31300 16000
rect 31352 15988 31358 16040
rect 53392 16028 53420 16059
rect 53466 16056 53472 16108
rect 53524 16096 53530 16108
rect 53929 16099 53987 16105
rect 53524 16068 53569 16096
rect 53524 16056 53530 16068
rect 53929 16065 53941 16099
rect 53975 16065 53987 16099
rect 53929 16059 53987 16065
rect 53944 16028 53972 16059
rect 53392 16000 53972 16028
rect 54205 16031 54263 16037
rect 54205 15997 54217 16031
rect 54251 16028 54263 16031
rect 55582 16028 55588 16040
rect 54251 16000 55588 16028
rect 54251 15997 54263 16000
rect 54205 15991 54263 15997
rect 55582 15988 55588 16000
rect 55640 15988 55646 16040
rect 53190 15960 53196 15972
rect 53151 15932 53196 15960
rect 53190 15920 53196 15932
rect 53248 15920 53254 15972
rect 24581 15895 24639 15901
rect 24581 15892 24593 15895
rect 18340 15864 24593 15892
rect 24581 15861 24593 15864
rect 24627 15892 24639 15895
rect 24762 15892 24768 15904
rect 24627 15864 24768 15892
rect 24627 15861 24639 15864
rect 24581 15855 24639 15861
rect 24762 15852 24768 15864
rect 24820 15852 24826 15904
rect 25774 15852 25780 15904
rect 25832 15892 25838 15904
rect 25958 15892 25964 15904
rect 25832 15864 25964 15892
rect 25832 15852 25838 15864
rect 25958 15852 25964 15864
rect 26016 15852 26022 15904
rect 27522 15852 27528 15904
rect 27580 15892 27586 15904
rect 30285 15895 30343 15901
rect 30285 15892 30297 15895
rect 27580 15864 30297 15892
rect 27580 15852 27586 15864
rect 30285 15861 30297 15864
rect 30331 15861 30343 15895
rect 30285 15855 30343 15861
rect 32766 15852 32772 15904
rect 32824 15892 32830 15904
rect 33965 15895 34023 15901
rect 33965 15892 33977 15895
rect 32824 15864 33977 15892
rect 32824 15852 32830 15864
rect 33965 15861 33977 15864
rect 34011 15861 34023 15895
rect 43714 15892 43720 15904
rect 43675 15864 43720 15892
rect 33965 15855 34023 15861
rect 43714 15852 43720 15864
rect 43772 15852 43778 15904
rect 51534 15892 51540 15904
rect 51495 15864 51540 15892
rect 51534 15852 51540 15864
rect 51592 15852 51598 15904
rect 52546 15852 52552 15904
rect 52604 15892 52610 15904
rect 53466 15892 53472 15904
rect 52604 15864 53472 15892
rect 52604 15852 52610 15864
rect 53466 15852 53472 15864
rect 53524 15892 53530 15904
rect 54021 15895 54079 15901
rect 54021 15892 54033 15895
rect 53524 15864 54033 15892
rect 53524 15852 53530 15864
rect 54021 15861 54033 15864
rect 54067 15892 54079 15895
rect 55398 15892 55404 15904
rect 54067 15864 55404 15892
rect 54067 15861 54079 15864
rect 54021 15855 54079 15861
rect 55398 15852 55404 15864
rect 55456 15852 55462 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2222 15648 2228 15700
rect 2280 15688 2286 15700
rect 23017 15691 23075 15697
rect 23017 15688 23029 15691
rect 2280 15660 23029 15688
rect 2280 15648 2286 15660
rect 23017 15657 23029 15660
rect 23063 15688 23075 15691
rect 23569 15691 23627 15697
rect 23569 15688 23581 15691
rect 23063 15660 23581 15688
rect 23063 15657 23075 15660
rect 23017 15651 23075 15657
rect 23569 15657 23581 15660
rect 23615 15657 23627 15691
rect 23750 15688 23756 15700
rect 23711 15660 23756 15688
rect 23569 15651 23627 15657
rect 23750 15648 23756 15660
rect 23808 15648 23814 15700
rect 24394 15688 24400 15700
rect 24355 15660 24400 15688
rect 24394 15648 24400 15660
rect 24452 15648 24458 15700
rect 24486 15648 24492 15700
rect 24544 15688 24550 15700
rect 43165 15691 43223 15697
rect 24544 15660 29868 15688
rect 24544 15648 24550 15660
rect 6546 15620 6552 15632
rect 6507 15592 6552 15620
rect 6546 15580 6552 15592
rect 6604 15580 6610 15632
rect 10594 15620 10600 15632
rect 10555 15592 10600 15620
rect 10594 15580 10600 15592
rect 10652 15580 10658 15632
rect 11882 15620 11888 15632
rect 11843 15592 11888 15620
rect 11882 15580 11888 15592
rect 11940 15580 11946 15632
rect 14458 15580 14464 15632
rect 14516 15620 14522 15632
rect 17405 15623 17463 15629
rect 17405 15620 17417 15623
rect 14516 15592 17417 15620
rect 14516 15580 14522 15592
rect 17405 15589 17417 15592
rect 17451 15589 17463 15623
rect 17770 15620 17776 15632
rect 17405 15583 17463 15589
rect 17604 15592 17776 15620
rect 5902 15512 5908 15564
rect 5960 15552 5966 15564
rect 6730 15552 6736 15564
rect 5960 15524 6736 15552
rect 5960 15512 5966 15524
rect 6730 15512 6736 15524
rect 6788 15552 6794 15564
rect 7101 15555 7159 15561
rect 7101 15552 7113 15555
rect 6788 15524 7113 15552
rect 6788 15512 6794 15524
rect 7101 15521 7113 15524
rect 7147 15521 7159 15555
rect 7101 15515 7159 15521
rect 16393 15555 16451 15561
rect 16393 15521 16405 15555
rect 16439 15552 16451 15555
rect 17034 15552 17040 15564
rect 16439 15524 17040 15552
rect 16439 15521 16451 15524
rect 16393 15515 16451 15521
rect 17034 15512 17040 15524
rect 17092 15552 17098 15564
rect 17218 15552 17224 15564
rect 17092 15524 17224 15552
rect 17092 15512 17098 15524
rect 17218 15512 17224 15524
rect 17276 15552 17282 15564
rect 17604 15552 17632 15592
rect 17770 15580 17776 15592
rect 17828 15580 17834 15632
rect 22066 15592 25084 15620
rect 17276 15524 17632 15552
rect 17681 15555 17739 15561
rect 17276 15512 17282 15524
rect 17681 15521 17693 15555
rect 17727 15552 17739 15555
rect 17727 15524 20300 15552
rect 17727 15521 17739 15524
rect 17681 15515 17739 15521
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15484 1455 15487
rect 1946 15484 1952 15496
rect 1443 15456 1952 15484
rect 1443 15453 1455 15456
rect 1397 15447 1455 15453
rect 1946 15444 1952 15456
rect 2004 15444 2010 15496
rect 2314 15484 2320 15496
rect 2275 15456 2320 15484
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 3844 15456 4077 15484
rect 3844 15444 3850 15456
rect 4065 15453 4077 15456
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 4332 15487 4390 15493
rect 4332 15453 4344 15487
rect 4378 15484 4390 15487
rect 4706 15484 4712 15496
rect 4378 15456 4712 15484
rect 4378 15453 4390 15456
rect 4332 15447 4390 15453
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 10781 15487 10839 15493
rect 10781 15453 10793 15487
rect 10827 15453 10839 15487
rect 10781 15447 10839 15453
rect 7009 15419 7067 15425
rect 7009 15416 7021 15419
rect 2148 15388 7021 15416
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 2148 15357 2176 15388
rect 7009 15385 7021 15388
rect 7055 15385 7067 15419
rect 10796 15416 10824 15447
rect 10870 15444 10876 15496
rect 10928 15484 10934 15496
rect 11054 15484 11060 15496
rect 10928 15456 10973 15484
rect 11015 15456 11060 15484
rect 10928 15444 10934 15456
rect 11054 15444 11060 15456
rect 11112 15444 11118 15496
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 13173 15487 13231 15493
rect 13173 15484 13185 15487
rect 11204 15456 11249 15484
rect 12406 15456 13185 15484
rect 11204 15444 11210 15456
rect 11606 15416 11612 15428
rect 10796 15388 11612 15416
rect 7009 15379 7067 15385
rect 11606 15376 11612 15388
rect 11664 15376 11670 15428
rect 11701 15419 11759 15425
rect 11701 15385 11713 15419
rect 11747 15416 11759 15419
rect 12406 15416 12434 15456
rect 13173 15453 13185 15456
rect 13219 15453 13231 15487
rect 13173 15447 13231 15453
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 13357 15487 13415 15493
rect 13357 15484 13369 15487
rect 13320 15456 13369 15484
rect 13320 15444 13326 15456
rect 13357 15453 13369 15456
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 15804 15456 16129 15484
rect 15804 15444 15810 15456
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 17586 15484 17592 15496
rect 17547 15456 17592 15484
rect 16117 15447 16175 15453
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 17770 15484 17776 15496
rect 17731 15456 17776 15484
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 17865 15487 17923 15493
rect 17865 15453 17877 15487
rect 17911 15453 17923 15487
rect 17865 15447 17923 15453
rect 11747 15388 12434 15416
rect 11747 15385 11759 15388
rect 11701 15379 11759 15385
rect 2133 15351 2191 15357
rect 2133 15317 2145 15351
rect 2179 15317 2191 15351
rect 5442 15348 5448 15360
rect 5403 15320 5448 15348
rect 2133 15311 2191 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 6917 15351 6975 15357
rect 6917 15317 6929 15351
rect 6963 15348 6975 15351
rect 8110 15348 8116 15360
rect 6963 15320 8116 15348
rect 6963 15317 6975 15320
rect 6917 15311 6975 15317
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 10318 15308 10324 15360
rect 10376 15348 10382 15360
rect 11716 15348 11744 15379
rect 17126 15376 17132 15428
rect 17184 15416 17190 15428
rect 17880 15416 17908 15447
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 20162 15484 20168 15496
rect 19484 15456 20168 15484
rect 19484 15444 19490 15456
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 20272 15484 20300 15524
rect 22066 15484 22094 15592
rect 23014 15512 23020 15564
rect 23072 15552 23078 15564
rect 23072 15524 24900 15552
rect 23072 15512 23078 15524
rect 24486 15484 24492 15496
rect 20272 15456 22094 15484
rect 23400 15456 24492 15484
rect 23400 15428 23428 15456
rect 24486 15444 24492 15456
rect 24544 15444 24550 15496
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15484 24639 15487
rect 24670 15484 24676 15496
rect 24627 15456 24676 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 24670 15444 24676 15456
rect 24728 15444 24734 15496
rect 24872 15493 24900 15524
rect 24857 15487 24915 15493
rect 24857 15453 24869 15487
rect 24903 15484 24915 15487
rect 24946 15484 24952 15496
rect 24903 15456 24952 15484
rect 24903 15453 24915 15456
rect 24857 15447 24915 15453
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 17184 15388 17908 15416
rect 20432 15419 20490 15425
rect 17184 15376 17190 15388
rect 20432 15385 20444 15419
rect 20478 15416 20490 15419
rect 21818 15416 21824 15428
rect 20478 15388 21824 15416
rect 20478 15385 20490 15388
rect 20432 15379 20490 15385
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 23382 15416 23388 15428
rect 23295 15388 23388 15416
rect 23382 15376 23388 15388
rect 23440 15376 23446 15428
rect 23569 15419 23627 15425
rect 23569 15385 23581 15419
rect 23615 15416 23627 15419
rect 25056 15416 25084 15592
rect 25406 15512 25412 15564
rect 25464 15552 25470 15564
rect 25961 15555 26019 15561
rect 25961 15552 25973 15555
rect 25464 15524 25973 15552
rect 25464 15512 25470 15524
rect 25961 15521 25973 15524
rect 26007 15521 26019 15555
rect 25961 15515 26019 15521
rect 29288 15524 29776 15552
rect 29288 15496 29316 15524
rect 29270 15484 29276 15496
rect 27356 15456 29276 15484
rect 25958 15416 25964 15428
rect 23615 15388 24900 15416
rect 25056 15388 25964 15416
rect 23615 15385 23627 15388
rect 23569 15379 23627 15385
rect 24872 15360 24900 15388
rect 25958 15376 25964 15388
rect 26016 15376 26022 15428
rect 26234 15425 26240 15428
rect 26228 15379 26240 15425
rect 26292 15416 26298 15428
rect 26292 15388 26328 15416
rect 26234 15376 26240 15379
rect 26292 15376 26298 15388
rect 10376 15320 11744 15348
rect 13265 15351 13323 15357
rect 10376 15308 10382 15320
rect 13265 15317 13277 15351
rect 13311 15348 13323 15351
rect 15194 15348 15200 15360
rect 13311 15320 15200 15348
rect 13311 15317 13323 15320
rect 13265 15311 13323 15317
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 21542 15348 21548 15360
rect 21503 15320 21548 15348
rect 21542 15308 21548 15320
rect 21600 15308 21606 15360
rect 24762 15348 24768 15360
rect 24723 15320 24768 15348
rect 24762 15308 24768 15320
rect 24820 15308 24826 15360
rect 24854 15308 24860 15360
rect 24912 15308 24918 15360
rect 27154 15308 27160 15360
rect 27212 15348 27218 15360
rect 27356 15357 27384 15456
rect 29270 15444 29276 15456
rect 29328 15444 29334 15496
rect 29748 15493 29776 15524
rect 29641 15487 29699 15493
rect 29641 15453 29653 15487
rect 29687 15453 29699 15487
rect 29641 15447 29699 15453
rect 29733 15487 29791 15493
rect 29733 15453 29745 15487
rect 29779 15453 29791 15487
rect 29840 15484 29868 15660
rect 43165 15657 43177 15691
rect 43211 15688 43223 15691
rect 43901 15691 43959 15697
rect 43901 15688 43913 15691
rect 43211 15660 43913 15688
rect 43211 15657 43223 15660
rect 43165 15651 43223 15657
rect 43901 15657 43913 15660
rect 43947 15688 43959 15691
rect 45922 15688 45928 15700
rect 43947 15660 45928 15688
rect 43947 15657 43959 15660
rect 43901 15651 43959 15657
rect 45922 15648 45928 15660
rect 45980 15648 45986 15700
rect 51534 15648 51540 15700
rect 51592 15688 51598 15700
rect 52273 15691 52331 15697
rect 52273 15688 52285 15691
rect 51592 15660 52285 15688
rect 51592 15648 51598 15660
rect 52273 15657 52285 15660
rect 52319 15657 52331 15691
rect 52914 15688 52920 15700
rect 52875 15660 52920 15688
rect 52273 15651 52331 15657
rect 52914 15648 52920 15660
rect 52972 15648 52978 15700
rect 41506 15580 41512 15632
rect 41564 15620 41570 15632
rect 41564 15592 44036 15620
rect 41564 15580 41570 15592
rect 30926 15512 30932 15564
rect 30984 15552 30990 15564
rect 32677 15555 32735 15561
rect 32677 15552 32689 15555
rect 30984 15524 32689 15552
rect 30984 15512 30990 15524
rect 32677 15521 32689 15524
rect 32723 15521 32735 15555
rect 42518 15552 42524 15564
rect 42479 15524 42524 15552
rect 32677 15515 32735 15521
rect 42518 15512 42524 15524
rect 42576 15512 42582 15564
rect 43006 15555 43064 15561
rect 43006 15521 43018 15555
rect 43052 15552 43064 15555
rect 43622 15552 43628 15564
rect 43052 15524 43628 15552
rect 43052 15521 43064 15524
rect 43006 15515 43064 15521
rect 43622 15512 43628 15524
rect 43680 15512 43686 15564
rect 32766 15484 32772 15496
rect 29840 15456 31754 15484
rect 32727 15456 32772 15484
rect 29733 15447 29791 15453
rect 29086 15376 29092 15428
rect 29144 15416 29150 15428
rect 29656 15416 29684 15447
rect 29822 15416 29828 15428
rect 29144 15388 29828 15416
rect 29144 15376 29150 15388
rect 29822 15376 29828 15388
rect 29880 15416 29886 15428
rect 30190 15416 30196 15428
rect 29880 15388 30196 15416
rect 29880 15376 29886 15388
rect 30190 15376 30196 15388
rect 30248 15376 30254 15428
rect 31726 15416 31754 15456
rect 32766 15444 32772 15456
rect 32824 15444 32830 15496
rect 42797 15487 42855 15493
rect 42797 15453 42809 15487
rect 42843 15484 42855 15487
rect 43530 15484 43536 15496
rect 42843 15456 43536 15484
rect 42843 15453 42855 15456
rect 42797 15447 42855 15453
rect 43530 15444 43536 15456
rect 43588 15444 43594 15496
rect 43714 15484 43720 15496
rect 43675 15456 43720 15484
rect 43714 15444 43720 15456
rect 43772 15444 43778 15496
rect 44008 15493 44036 15592
rect 52454 15580 52460 15632
rect 52512 15620 52518 15632
rect 53098 15620 53104 15632
rect 52512 15592 53104 15620
rect 52512 15580 52518 15592
rect 53098 15580 53104 15592
rect 53156 15620 53162 15632
rect 53374 15620 53380 15632
rect 53156 15592 53380 15620
rect 53156 15580 53162 15592
rect 53374 15580 53380 15592
rect 53432 15580 53438 15632
rect 52546 15552 52552 15564
rect 52196 15524 52552 15552
rect 43993 15487 44051 15493
rect 43993 15453 44005 15487
rect 44039 15453 44051 15487
rect 48038 15484 48044 15496
rect 47999 15456 48044 15484
rect 43993 15447 44051 15453
rect 48038 15444 48044 15456
rect 48096 15444 48102 15496
rect 52196 15493 52224 15524
rect 52546 15512 52552 15524
rect 52604 15512 52610 15564
rect 53193 15555 53251 15561
rect 53193 15521 53205 15555
rect 53239 15552 53251 15555
rect 54018 15552 54024 15564
rect 53239 15524 54024 15552
rect 53239 15521 53251 15524
rect 53193 15515 53251 15521
rect 54018 15512 54024 15524
rect 54076 15512 54082 15564
rect 52181 15487 52239 15493
rect 52181 15453 52193 15487
rect 52227 15453 52239 15487
rect 52454 15484 52460 15496
rect 52415 15456 52460 15484
rect 52181 15447 52239 15453
rect 52454 15444 52460 15456
rect 52512 15444 52518 15496
rect 53101 15487 53159 15493
rect 53101 15453 53113 15487
rect 53147 15453 53159 15487
rect 53282 15484 53288 15496
rect 53243 15456 53288 15484
rect 53101 15447 53159 15453
rect 40402 15416 40408 15428
rect 31726 15388 40408 15416
rect 40402 15376 40408 15388
rect 40460 15376 40466 15428
rect 42242 15376 42248 15428
rect 42300 15416 42306 15428
rect 43625 15419 43683 15425
rect 43625 15416 43637 15419
rect 42300 15388 43637 15416
rect 42300 15376 42306 15388
rect 43625 15385 43637 15388
rect 43671 15385 43683 15419
rect 44082 15416 44088 15428
rect 44043 15388 44088 15416
rect 43625 15379 43683 15385
rect 44082 15376 44088 15388
rect 44140 15376 44146 15428
rect 52365 15419 52423 15425
rect 52365 15385 52377 15419
rect 52411 15385 52423 15419
rect 53116 15416 53144 15447
rect 53282 15444 53288 15456
rect 53340 15444 53346 15496
rect 53374 15444 53380 15496
rect 53432 15484 53438 15496
rect 53432 15456 53477 15484
rect 53432 15444 53438 15456
rect 53834 15444 53840 15496
rect 53892 15484 53898 15496
rect 53929 15487 53987 15493
rect 53929 15484 53941 15487
rect 53892 15456 53941 15484
rect 53892 15444 53898 15456
rect 53929 15453 53941 15456
rect 53975 15453 53987 15487
rect 55674 15484 55680 15496
rect 55635 15456 55680 15484
rect 53929 15447 53987 15453
rect 55674 15444 55680 15456
rect 55732 15444 55738 15496
rect 55861 15487 55919 15493
rect 55861 15453 55873 15487
rect 55907 15453 55919 15487
rect 55861 15447 55919 15453
rect 55214 15416 55220 15428
rect 53116 15388 55220 15416
rect 52365 15379 52423 15385
rect 27341 15351 27399 15357
rect 27341 15348 27353 15351
rect 27212 15320 27353 15348
rect 27212 15308 27218 15320
rect 27341 15317 27353 15320
rect 27387 15317 27399 15351
rect 27341 15311 27399 15317
rect 28994 15308 29000 15360
rect 29052 15348 29058 15360
rect 29917 15351 29975 15357
rect 29917 15348 29929 15351
rect 29052 15320 29929 15348
rect 29052 15308 29058 15320
rect 29917 15317 29929 15320
rect 29963 15348 29975 15351
rect 30006 15348 30012 15360
rect 29963 15320 30012 15348
rect 29963 15317 29975 15320
rect 29917 15311 29975 15317
rect 30006 15308 30012 15320
rect 30064 15308 30070 15360
rect 33137 15351 33195 15357
rect 33137 15317 33149 15351
rect 33183 15348 33195 15351
rect 33502 15348 33508 15360
rect 33183 15320 33508 15348
rect 33183 15317 33195 15320
rect 33137 15311 33195 15317
rect 33502 15308 33508 15320
rect 33560 15308 33566 15360
rect 42886 15308 42892 15360
rect 42944 15348 42950 15360
rect 47854 15348 47860 15360
rect 42944 15320 42989 15348
rect 47815 15320 47860 15348
rect 42944 15308 42950 15320
rect 47854 15308 47860 15320
rect 47912 15308 47918 15360
rect 52380 15348 52408 15379
rect 55214 15376 55220 15388
rect 55272 15376 55278 15428
rect 55398 15376 55404 15428
rect 55456 15416 55462 15428
rect 55876 15416 55904 15447
rect 55456 15388 55904 15416
rect 55456 15376 55462 15388
rect 53282 15348 53288 15360
rect 52380 15320 53288 15348
rect 53282 15308 53288 15320
rect 53340 15348 53346 15360
rect 54159 15351 54217 15357
rect 54159 15348 54171 15351
rect 53340 15320 54171 15348
rect 53340 15308 53346 15320
rect 54159 15317 54171 15320
rect 54205 15317 54217 15351
rect 55766 15348 55772 15360
rect 55727 15320 55772 15348
rect 54159 15311 54217 15317
rect 55766 15308 55772 15320
rect 55824 15308 55830 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 4525 15147 4583 15153
rect 4525 15113 4537 15147
rect 4571 15144 4583 15147
rect 4614 15144 4620 15156
rect 4571 15116 4620 15144
rect 4571 15113 4583 15116
rect 4525 15107 4583 15113
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 7006 15104 7012 15156
rect 7064 15144 7070 15156
rect 11517 15147 11575 15153
rect 7064 15116 7972 15144
rect 7064 15104 7070 15116
rect 2498 15036 2504 15088
rect 2556 15076 2562 15088
rect 2556 15048 6132 15076
rect 2556 15036 2562 15048
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 14968 1458 15020
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 15008 2375 15011
rect 2774 15008 2780 15020
rect 2363 14980 2780 15008
rect 2363 14977 2375 14980
rect 2317 14971 2375 14977
rect 2774 14968 2780 14980
rect 2832 14968 2838 15020
rect 4893 15011 4951 15017
rect 4893 14977 4905 15011
rect 4939 15008 4951 15011
rect 5442 15008 5448 15020
rect 4939 14980 5448 15008
rect 4939 14977 4951 14980
rect 4893 14971 4951 14977
rect 5442 14968 5448 14980
rect 5500 14968 5506 15020
rect 4985 14943 5043 14949
rect 4985 14940 4997 14943
rect 2746 14912 4997 14940
rect 2133 14875 2191 14881
rect 2133 14841 2145 14875
rect 2179 14872 2191 14875
rect 2746 14872 2774 14912
rect 4985 14909 4997 14912
rect 5031 14909 5043 14943
rect 4985 14903 5043 14909
rect 5169 14943 5227 14949
rect 5169 14909 5181 14943
rect 5215 14940 5227 14943
rect 5902 14940 5908 14952
rect 5215 14912 5908 14940
rect 5215 14909 5227 14912
rect 5169 14903 5227 14909
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 2179 14844 2774 14872
rect 6104 14872 6132 15048
rect 6178 15036 6184 15088
rect 6236 15076 6242 15088
rect 6236 15048 7880 15076
rect 6236 15036 6242 15048
rect 7466 14968 7472 15020
rect 7524 15008 7530 15020
rect 7852 15017 7880 15048
rect 7944 15017 7972 15116
rect 11517 15113 11529 15147
rect 11563 15144 11575 15147
rect 12526 15144 12532 15156
rect 11563 15116 12532 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 12713 15147 12771 15153
rect 12713 15113 12725 15147
rect 12759 15113 12771 15147
rect 16114 15144 16120 15156
rect 12713 15107 12771 15113
rect 13004 15116 16120 15144
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 12728 15076 12756 15107
rect 11664 15048 12756 15076
rect 11664 15036 11670 15048
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 7524 14980 7573 15008
rect 7524 14968 7530 14980
rect 7561 14977 7573 14980
rect 7607 14977 7619 15011
rect 7561 14971 7619 14977
rect 7653 15011 7711 15017
rect 7653 14977 7665 15011
rect 7699 15008 7711 15011
rect 7837 15011 7895 15017
rect 7699 14980 7788 15008
rect 7699 14977 7711 14980
rect 7653 14971 7711 14977
rect 7760 14872 7788 14980
rect 7837 14977 7849 15011
rect 7883 14977 7895 15011
rect 7837 14971 7895 14977
rect 7929 15011 7987 15017
rect 7929 14977 7941 15011
rect 7975 14977 7987 15011
rect 7929 14971 7987 14977
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 13004 15008 13032 15116
rect 16114 15104 16120 15116
rect 16172 15144 16178 15156
rect 16172 15116 17540 15144
rect 16172 15104 16178 15116
rect 13173 15079 13231 15085
rect 13173 15045 13185 15079
rect 13219 15076 13231 15079
rect 16390 15076 16396 15088
rect 13219 15048 16396 15076
rect 13219 15045 13231 15048
rect 13173 15039 13231 15045
rect 16390 15036 16396 15048
rect 16448 15036 16454 15088
rect 17126 15036 17132 15088
rect 17184 15036 17190 15088
rect 17512 15076 17540 15116
rect 17586 15104 17592 15156
rect 17644 15144 17650 15156
rect 17865 15147 17923 15153
rect 17865 15144 17877 15147
rect 17644 15116 17877 15144
rect 17644 15104 17650 15116
rect 17865 15113 17877 15116
rect 17911 15113 17923 15147
rect 21818 15144 21824 15156
rect 21779 15116 21824 15144
rect 17865 15107 17923 15113
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 23474 15144 23480 15156
rect 23435 15116 23480 15144
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 23934 15144 23940 15156
rect 23895 15116 23940 15144
rect 23934 15104 23940 15116
rect 23992 15104 23998 15156
rect 24670 15144 24676 15156
rect 24583 15116 24676 15144
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 25869 15147 25927 15153
rect 25869 15113 25881 15147
rect 25915 15144 25927 15147
rect 26234 15144 26240 15156
rect 25915 15116 26240 15144
rect 25915 15113 25927 15116
rect 25869 15107 25927 15113
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 29181 15147 29239 15153
rect 29181 15113 29193 15147
rect 29227 15144 29239 15147
rect 29270 15144 29276 15156
rect 29227 15116 29276 15144
rect 29227 15113 29239 15116
rect 29181 15107 29239 15113
rect 29270 15104 29276 15116
rect 29328 15104 29334 15156
rect 30006 15104 30012 15156
rect 30064 15144 30070 15156
rect 30926 15144 30932 15156
rect 30064 15116 30788 15144
rect 30887 15116 30932 15144
rect 30064 15104 30070 15116
rect 17954 15076 17960 15088
rect 17512 15048 17960 15076
rect 17954 15036 17960 15048
rect 18012 15076 18018 15088
rect 22189 15079 22247 15085
rect 22189 15076 22201 15079
rect 18012 15048 18184 15076
rect 18012 15036 18018 15048
rect 11931 14980 13032 15008
rect 13081 15011 13139 15017
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 13081 14977 13093 15011
rect 13127 15008 13139 15011
rect 14090 15008 14096 15020
rect 13127 14980 14096 15008
rect 13127 14977 13139 14980
rect 13081 14971 13139 14977
rect 7852 14940 7880 14971
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 17144 15008 17172 15036
rect 17313 15011 17371 15017
rect 17313 15008 17325 15011
rect 17144 14980 17325 15008
rect 17313 14977 17325 14980
rect 17359 14977 17371 15011
rect 17313 14971 17371 14977
rect 17494 14968 17500 15020
rect 17552 15008 17558 15020
rect 17862 15008 17868 15020
rect 17552 14980 17868 15008
rect 17552 14968 17558 14980
rect 17862 14968 17868 14980
rect 17920 15008 17926 15020
rect 18156 15017 18184 15048
rect 21560 15048 22201 15076
rect 21560 15020 21588 15048
rect 22189 15045 22201 15048
rect 22235 15045 22247 15079
rect 23014 15076 23020 15088
rect 22189 15039 22247 15045
rect 22296 15048 23020 15076
rect 18049 15011 18107 15017
rect 18049 15008 18061 15011
rect 17920 14980 18061 15008
rect 17920 14968 17926 14980
rect 18049 14977 18061 14980
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 18141 15011 18199 15017
rect 18141 14977 18153 15011
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 15008 18291 15011
rect 21542 15008 21548 15020
rect 18279 14980 21548 15008
rect 18279 14977 18291 14980
rect 18233 14971 18291 14977
rect 21542 14968 21548 14980
rect 21600 14968 21606 15020
rect 22296 15017 22324 15048
rect 23014 15036 23020 15048
rect 23072 15036 23078 15088
rect 24302 15076 24308 15088
rect 24263 15048 24308 15076
rect 24302 15036 24308 15048
rect 24360 15036 24366 15088
rect 24688 15076 24716 15104
rect 24535 15045 24593 15051
rect 24688 15048 26372 15076
rect 24535 15042 24547 15045
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22281 15011 22339 15017
rect 22281 14977 22293 15011
rect 22327 14977 22339 15011
rect 22830 15008 22836 15020
rect 22791 14980 22836 15008
rect 22281 14971 22339 14977
rect 8018 14940 8024 14952
rect 7852 14912 8024 14940
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 11977 14943 12035 14949
rect 11977 14940 11989 14943
rect 11900 14912 11989 14940
rect 11900 14884 11928 14912
rect 11977 14909 11989 14912
rect 12023 14909 12035 14943
rect 11977 14903 12035 14909
rect 12066 14900 12072 14952
rect 12124 14940 12130 14952
rect 12124 14912 12169 14940
rect 12124 14900 12130 14912
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 17034 14940 17040 14952
rect 13320 14912 13365 14940
rect 16995 14912 17040 14940
rect 13320 14900 13326 14912
rect 17034 14900 17040 14912
rect 17092 14900 17098 14952
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14909 17187 14943
rect 17129 14903 17187 14909
rect 8478 14872 8484 14884
rect 6104 14844 7604 14872
rect 7760 14844 8484 14872
rect 2179 14841 2191 14844
rect 2133 14835 2191 14841
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 7282 14804 7288 14816
rect 1627 14776 7288 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 7377 14807 7435 14813
rect 7377 14773 7389 14807
rect 7423 14804 7435 14807
rect 7466 14804 7472 14816
rect 7423 14776 7472 14804
rect 7423 14773 7435 14776
rect 7377 14767 7435 14773
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 7576 14804 7604 14844
rect 8478 14832 8484 14844
rect 8536 14832 8542 14884
rect 11882 14832 11888 14884
rect 11940 14832 11946 14884
rect 16853 14875 16911 14881
rect 16853 14872 16865 14875
rect 11992 14844 16865 14872
rect 11992 14804 12020 14844
rect 16853 14841 16865 14844
rect 16899 14841 16911 14875
rect 16853 14835 16911 14841
rect 7576 14776 12020 14804
rect 12066 14764 12072 14816
rect 12124 14804 12130 14816
rect 16666 14804 16672 14816
rect 12124 14776 16672 14804
rect 12124 14764 12130 14776
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 17144 14804 17172 14903
rect 17218 14900 17224 14952
rect 17276 14940 17282 14952
rect 17276 14912 17321 14940
rect 17276 14900 17282 14912
rect 17770 14900 17776 14952
rect 17828 14940 17834 14952
rect 18325 14943 18383 14949
rect 18325 14940 18337 14943
rect 17828 14912 18337 14940
rect 17828 14900 17834 14912
rect 18325 14909 18337 14912
rect 18371 14909 18383 14943
rect 22020 14940 22048 14971
rect 22830 14968 22836 14980
rect 22888 14968 22894 15020
rect 23382 14968 23388 15020
rect 23440 15008 23446 15020
rect 23661 15011 23719 15017
rect 23661 15008 23673 15011
rect 23440 14980 23673 15008
rect 23440 14968 23446 14980
rect 23661 14977 23673 14980
rect 23707 14977 23719 15011
rect 23661 14971 23719 14977
rect 24026 14968 24032 15020
rect 24084 15008 24090 15020
rect 24520 15011 24547 15042
rect 24581 15011 24593 15045
rect 26344 15017 26372 15048
rect 26418 15036 26424 15088
rect 26476 15076 26482 15088
rect 29822 15076 29828 15088
rect 26476 15048 29828 15076
rect 26476 15036 26482 15048
rect 29822 15036 29828 15048
rect 29880 15036 29886 15088
rect 30024 15048 30604 15076
rect 24520 15008 24593 15011
rect 26329 15011 26387 15017
rect 24084 14980 25084 15008
rect 24084 14968 24090 14980
rect 23842 14940 23848 14952
rect 22020 14912 23848 14940
rect 18325 14903 18383 14909
rect 23842 14900 23848 14912
rect 23900 14900 23906 14952
rect 24946 14872 24952 14884
rect 22066 14844 24952 14872
rect 22066 14804 22094 14844
rect 24946 14832 24952 14844
rect 25004 14832 25010 14884
rect 17144 14776 22094 14804
rect 23934 14764 23940 14816
rect 23992 14804 23998 14816
rect 24486 14804 24492 14816
rect 23992 14776 24492 14804
rect 23992 14764 23998 14776
rect 24486 14764 24492 14776
rect 24544 14764 24550 14816
rect 25056 14804 25084 14980
rect 26329 14977 26341 15011
rect 26375 14977 26387 15011
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26329 14971 26387 14977
rect 26896 14980 26985 15008
rect 26896 14952 26924 14980
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 27154 15008 27160 15020
rect 27115 14980 27160 15008
rect 26973 14971 27031 14977
rect 27154 14968 27160 14980
rect 27212 14968 27218 15020
rect 28997 15011 29055 15017
rect 28997 14977 29009 15011
rect 29043 15008 29055 15011
rect 29086 15008 29092 15020
rect 29043 14980 29092 15008
rect 29043 14977 29055 14980
rect 28997 14971 29055 14977
rect 29086 14968 29092 14980
rect 29144 14968 29150 15020
rect 29270 15008 29276 15020
rect 29231 14980 29276 15008
rect 29270 14968 29276 14980
rect 29328 14968 29334 15020
rect 29917 15011 29975 15017
rect 29917 14977 29929 15011
rect 29963 15008 29975 15011
rect 30024 15008 30052 15048
rect 29963 14980 30052 15008
rect 30101 15011 30159 15017
rect 29963 14977 29975 14980
rect 29917 14971 29975 14977
rect 30101 14977 30113 15011
rect 30147 15008 30159 15011
rect 30466 15008 30472 15020
rect 30147 14980 30472 15008
rect 30147 14977 30159 14980
rect 30101 14971 30159 14977
rect 30466 14968 30472 14980
rect 30524 14968 30530 15020
rect 26050 14940 26056 14952
rect 26011 14912 26056 14940
rect 26050 14900 26056 14912
rect 26108 14900 26114 14952
rect 26145 14943 26203 14949
rect 26145 14909 26157 14943
rect 26191 14909 26203 14943
rect 26145 14903 26203 14909
rect 26237 14943 26295 14949
rect 26237 14909 26249 14943
rect 26283 14940 26295 14943
rect 26418 14940 26424 14952
rect 26283 14912 26424 14940
rect 26283 14909 26295 14912
rect 26237 14903 26295 14909
rect 26160 14872 26188 14903
rect 26418 14900 26424 14912
rect 26476 14900 26482 14952
rect 26878 14940 26884 14952
rect 26791 14912 26884 14940
rect 26878 14900 26884 14912
rect 26936 14940 26942 14952
rect 29285 14940 29313 14968
rect 26936 14912 29313 14940
rect 30009 14943 30067 14949
rect 26936 14900 26942 14912
rect 30009 14909 30021 14943
rect 30055 14909 30067 14943
rect 30009 14903 30067 14909
rect 30193 14943 30251 14949
rect 30193 14909 30205 14943
rect 30239 14940 30251 14943
rect 30374 14940 30380 14952
rect 30239 14912 30380 14940
rect 30239 14909 30251 14912
rect 30193 14903 30251 14909
rect 27065 14875 27123 14881
rect 27065 14872 27077 14875
rect 26160 14844 27077 14872
rect 27065 14841 27077 14844
rect 27111 14841 27123 14875
rect 27065 14835 27123 14841
rect 28813 14875 28871 14881
rect 28813 14841 28825 14875
rect 28859 14872 28871 14875
rect 30025 14872 30053 14903
rect 30374 14900 30380 14912
rect 30432 14900 30438 14952
rect 30576 14940 30604 15048
rect 30760 15017 30788 15116
rect 30926 15104 30932 15116
rect 30984 15104 30990 15156
rect 32858 15144 32864 15156
rect 32819 15116 32864 15144
rect 32858 15104 32864 15116
rect 32916 15104 32922 15156
rect 38930 15104 38936 15156
rect 38988 15144 38994 15156
rect 41506 15144 41512 15156
rect 38988 15116 41512 15144
rect 38988 15104 38994 15116
rect 41506 15104 41512 15116
rect 41564 15104 41570 15156
rect 41601 15147 41659 15153
rect 41601 15113 41613 15147
rect 41647 15144 41659 15147
rect 42886 15144 42892 15156
rect 41647 15116 42892 15144
rect 41647 15113 41659 15116
rect 41601 15107 41659 15113
rect 42886 15104 42892 15116
rect 42944 15104 42950 15156
rect 45002 15144 45008 15156
rect 44963 15116 45008 15144
rect 45002 15104 45008 15116
rect 45060 15104 45066 15156
rect 53558 15144 53564 15156
rect 45204 15116 53564 15144
rect 30944 15076 30972 15104
rect 33502 15076 33508 15088
rect 30852 15048 30972 15076
rect 33463 15048 33508 15076
rect 30745 15011 30803 15017
rect 30745 14977 30757 15011
rect 30791 14977 30803 15011
rect 30745 14971 30803 14977
rect 30852 14940 30880 15048
rect 33502 15036 33508 15048
rect 33560 15036 33566 15088
rect 37826 15036 37832 15088
rect 37884 15076 37890 15088
rect 39025 15079 39083 15085
rect 39025 15076 39037 15079
rect 37884 15048 39037 15076
rect 37884 15036 37890 15048
rect 39025 15045 39037 15048
rect 39071 15045 39083 15079
rect 39025 15039 39083 15045
rect 39117 15079 39175 15085
rect 39117 15045 39129 15079
rect 39163 15076 39175 15079
rect 40957 15079 41015 15085
rect 40957 15076 40969 15079
rect 39163 15048 40969 15076
rect 39163 15045 39175 15048
rect 39117 15039 39175 15045
rect 40957 15045 40969 15048
rect 41003 15045 41015 15079
rect 40957 15039 41015 15045
rect 30926 14968 30932 15020
rect 30984 15008 30990 15020
rect 33134 15008 33140 15020
rect 30984 14980 31029 15008
rect 33095 14980 33140 15008
rect 30984 14968 30990 14980
rect 33134 14968 33140 14980
rect 33192 14968 33198 15020
rect 33318 14968 33324 15020
rect 33376 15008 33382 15020
rect 33413 15011 33471 15017
rect 33413 15008 33425 15011
rect 33376 14980 33425 15008
rect 33376 14968 33382 14980
rect 33413 14977 33425 14980
rect 33459 14977 33471 15011
rect 33413 14971 33471 14977
rect 38749 15011 38807 15017
rect 38749 14977 38761 15011
rect 38795 15008 38807 15011
rect 38838 15008 38844 15020
rect 38795 14980 38844 15008
rect 38795 14977 38807 14980
rect 38749 14971 38807 14977
rect 38838 14968 38844 14980
rect 38896 14968 38902 15020
rect 40310 14968 40316 15020
rect 40368 15008 40374 15020
rect 40589 15011 40647 15017
rect 40589 15008 40601 15011
rect 40368 14980 40601 15008
rect 40368 14968 40374 14980
rect 40589 14977 40601 14980
rect 40635 14977 40647 15011
rect 40589 14971 40647 14977
rect 40773 15011 40831 15017
rect 40773 14977 40785 15011
rect 40819 14977 40831 15011
rect 40972 15008 41000 15039
rect 41046 15036 41052 15088
rect 41104 15076 41110 15088
rect 42794 15076 42800 15088
rect 41104 15048 42800 15076
rect 41104 15036 41110 15048
rect 42794 15036 42800 15048
rect 42852 15076 42858 15088
rect 43162 15076 43168 15088
rect 42852 15048 43168 15076
rect 42852 15036 42858 15048
rect 43162 15036 43168 15048
rect 43220 15036 43226 15088
rect 43892 15079 43950 15085
rect 43892 15045 43904 15079
rect 43938 15076 43950 15079
rect 44082 15076 44088 15088
rect 43938 15048 44088 15076
rect 43938 15045 43950 15048
rect 43892 15039 43950 15045
rect 44082 15036 44088 15048
rect 44140 15036 44146 15088
rect 41417 15011 41475 15017
rect 41417 15008 41429 15011
rect 40972 14980 41429 15008
rect 40773 14971 40831 14977
rect 41417 14977 41429 14980
rect 41463 14977 41475 15011
rect 41598 15008 41604 15020
rect 41559 14980 41604 15008
rect 41417 14971 41475 14977
rect 30576 14912 30880 14940
rect 33045 14943 33103 14949
rect 33045 14909 33057 14943
rect 33091 14940 33103 14943
rect 38657 14943 38715 14949
rect 33091 14912 33456 14940
rect 33091 14909 33103 14912
rect 33045 14903 33103 14909
rect 33428 14884 33456 14912
rect 38657 14909 38669 14943
rect 38703 14940 38715 14943
rect 38930 14940 38936 14952
rect 38703 14912 38936 14940
rect 38703 14909 38715 14912
rect 38657 14903 38715 14909
rect 38930 14900 38936 14912
rect 38988 14900 38994 14952
rect 40788 14940 40816 14971
rect 41598 14968 41604 14980
rect 41656 14968 41662 15020
rect 45204 15008 45232 15116
rect 53558 15104 53564 15116
rect 53616 15104 53622 15156
rect 55030 15104 55036 15156
rect 55088 15144 55094 15156
rect 57333 15147 57391 15153
rect 57333 15144 57345 15147
rect 55088 15116 57345 15144
rect 55088 15104 55094 15116
rect 57333 15113 57345 15116
rect 57379 15113 57391 15147
rect 57333 15107 57391 15113
rect 47854 15085 47860 15088
rect 47848 15076 47860 15085
rect 47815 15048 47860 15076
rect 47848 15039 47860 15048
rect 47854 15036 47860 15039
rect 47912 15036 47918 15088
rect 50249 15079 50307 15085
rect 50249 15045 50261 15079
rect 50295 15076 50307 15079
rect 55398 15076 55404 15088
rect 50295 15048 51580 15076
rect 55359 15048 55404 15076
rect 50295 15045 50307 15048
rect 50249 15039 50307 15045
rect 42444 14980 45232 15008
rect 51077 15011 51135 15017
rect 41046 14940 41052 14952
rect 40788 14912 41052 14940
rect 41046 14900 41052 14912
rect 41104 14900 41110 14952
rect 28859 14844 30053 14872
rect 28859 14841 28871 14844
rect 28813 14835 28871 14841
rect 33410 14832 33416 14884
rect 33468 14832 33474 14884
rect 36446 14832 36452 14884
rect 36504 14872 36510 14884
rect 42444 14872 42472 14980
rect 51077 14977 51089 15011
rect 51123 14977 51135 15011
rect 51077 14971 51135 14977
rect 42518 14900 42524 14952
rect 42576 14940 42582 14952
rect 43070 14940 43076 14952
rect 42576 14912 43076 14940
rect 42576 14900 42582 14912
rect 43070 14900 43076 14912
rect 43128 14940 43134 14952
rect 43625 14943 43683 14949
rect 43625 14940 43637 14943
rect 43128 14912 43637 14940
rect 43128 14900 43134 14912
rect 43625 14909 43637 14912
rect 43671 14909 43683 14943
rect 43625 14903 43683 14909
rect 46014 14900 46020 14952
rect 46072 14940 46078 14952
rect 47581 14943 47639 14949
rect 47581 14940 47593 14943
rect 46072 14912 47593 14940
rect 46072 14900 46078 14912
rect 47581 14909 47593 14912
rect 47627 14909 47639 14943
rect 47581 14903 47639 14909
rect 48792 14912 50292 14940
rect 36504 14844 42472 14872
rect 36504 14832 36510 14844
rect 28534 14804 28540 14816
rect 25056 14776 28540 14804
rect 28534 14764 28540 14776
rect 28592 14764 28598 14816
rect 29733 14807 29791 14813
rect 29733 14773 29745 14807
rect 29779 14804 29791 14807
rect 29822 14804 29828 14816
rect 29779 14776 29828 14804
rect 29779 14773 29791 14776
rect 29733 14767 29791 14773
rect 29822 14764 29828 14776
rect 29880 14764 29886 14816
rect 38470 14804 38476 14816
rect 38431 14776 38476 14804
rect 38470 14764 38476 14776
rect 38528 14764 38534 14816
rect 38654 14764 38660 14816
rect 38712 14804 38718 14816
rect 48792 14804 48820 14912
rect 49050 14832 49056 14884
rect 49108 14872 49114 14884
rect 49881 14875 49939 14881
rect 49881 14872 49893 14875
rect 49108 14844 49893 14872
rect 49108 14832 49114 14844
rect 49881 14841 49893 14844
rect 49927 14841 49939 14875
rect 49881 14835 49939 14841
rect 48958 14804 48964 14816
rect 38712 14776 48820 14804
rect 48919 14776 48964 14804
rect 38712 14764 38718 14776
rect 48958 14764 48964 14776
rect 49016 14764 49022 14816
rect 50264 14813 50292 14912
rect 50433 14875 50491 14881
rect 50433 14841 50445 14875
rect 50479 14872 50491 14875
rect 51092 14872 51120 14971
rect 51552 14940 51580 15048
rect 55398 15036 55404 15048
rect 55456 15036 55462 15088
rect 55766 15036 55772 15088
rect 55824 15076 55830 15088
rect 56198 15079 56256 15085
rect 56198 15076 56210 15079
rect 55824 15048 56210 15076
rect 55824 15036 55830 15048
rect 56198 15045 56210 15048
rect 56244 15045 56256 15079
rect 56198 15039 56256 15045
rect 52546 14968 52552 15020
rect 52604 15008 52610 15020
rect 52917 15011 52975 15017
rect 52917 15008 52929 15011
rect 52604 14980 52929 15008
rect 52604 14968 52610 14980
rect 52917 14977 52929 14980
rect 52963 14977 52975 15011
rect 52917 14971 52975 14977
rect 53009 15011 53067 15017
rect 53009 14977 53021 15011
rect 53055 15008 53067 15011
rect 53282 15008 53288 15020
rect 53055 14980 53288 15008
rect 53055 14977 53067 14980
rect 53009 14971 53067 14977
rect 53282 14968 53288 14980
rect 53340 14968 53346 15020
rect 55214 14968 55220 15020
rect 55272 15008 55278 15020
rect 55272 14980 55317 15008
rect 55272 14968 55278 14980
rect 52733 14943 52791 14949
rect 52733 14940 52745 14943
rect 51552 14912 52745 14940
rect 52733 14909 52745 14912
rect 52779 14909 52791 14943
rect 53098 14940 53104 14952
rect 53059 14912 53104 14940
rect 52733 14903 52791 14909
rect 53098 14900 53104 14912
rect 53156 14900 53162 14952
rect 53190 14900 53196 14952
rect 53248 14940 53254 14952
rect 53248 14912 53293 14940
rect 53248 14900 53254 14912
rect 54018 14900 54024 14952
rect 54076 14940 54082 14952
rect 55030 14940 55036 14952
rect 54076 14912 55036 14940
rect 54076 14900 54082 14912
rect 55030 14900 55036 14912
rect 55088 14900 55094 14952
rect 55953 14943 56011 14949
rect 55953 14909 55965 14943
rect 55999 14909 56011 14943
rect 55953 14903 56011 14909
rect 50479 14844 51120 14872
rect 50479 14841 50491 14844
rect 50433 14835 50491 14841
rect 50249 14807 50307 14813
rect 50249 14773 50261 14807
rect 50295 14804 50307 14807
rect 50614 14804 50620 14816
rect 50295 14776 50620 14804
rect 50295 14773 50307 14776
rect 50249 14767 50307 14773
rect 50614 14764 50620 14776
rect 50672 14764 50678 14816
rect 50890 14804 50896 14816
rect 50851 14776 50896 14804
rect 50890 14764 50896 14776
rect 50948 14764 50954 14816
rect 55968 14804 55996 14903
rect 56318 14804 56324 14816
rect 55968 14776 56324 14804
rect 56318 14764 56324 14776
rect 56376 14764 56382 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2682 14600 2688 14612
rect 2004 14572 2688 14600
rect 2004 14560 2010 14572
rect 2682 14560 2688 14572
rect 2740 14600 2746 14612
rect 2961 14603 3019 14609
rect 2961 14600 2973 14603
rect 2740 14572 2973 14600
rect 2740 14560 2746 14572
rect 2961 14569 2973 14572
rect 3007 14569 3019 14603
rect 2961 14563 3019 14569
rect 5442 14560 5448 14612
rect 5500 14600 5506 14612
rect 7834 14600 7840 14612
rect 5500 14572 7840 14600
rect 5500 14560 5506 14572
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 8021 14603 8079 14609
rect 8021 14569 8033 14603
rect 8067 14600 8079 14603
rect 8110 14600 8116 14612
rect 8067 14572 8116 14600
rect 8067 14569 8079 14572
rect 8021 14563 8079 14569
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 14090 14600 14096 14612
rect 14051 14572 14096 14600
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 14461 14603 14519 14609
rect 14461 14569 14473 14603
rect 14507 14600 14519 14603
rect 16022 14600 16028 14612
rect 14507 14572 16028 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 16022 14560 16028 14572
rect 16080 14560 16086 14612
rect 17034 14560 17040 14612
rect 17092 14600 17098 14612
rect 17313 14603 17371 14609
rect 17313 14600 17325 14603
rect 17092 14572 17325 14600
rect 17092 14560 17098 14572
rect 17313 14569 17325 14572
rect 17359 14569 17371 14603
rect 17313 14563 17371 14569
rect 17586 14560 17592 14612
rect 17644 14600 17650 14612
rect 17954 14600 17960 14612
rect 17644 14572 17960 14600
rect 17644 14560 17650 14572
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 23382 14600 23388 14612
rect 19352 14572 23388 14600
rect 14550 14532 14556 14544
rect 2746 14504 14556 14532
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 2590 14396 2596 14408
rect 1627 14368 2596 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 1848 14331 1906 14337
rect 1848 14297 1860 14331
rect 1894 14328 1906 14331
rect 2314 14328 2320 14340
rect 1894 14300 2320 14328
rect 1894 14297 1906 14300
rect 1848 14291 1906 14297
rect 2314 14288 2320 14300
rect 2372 14288 2378 14340
rect 2746 14328 2774 14504
rect 14550 14492 14556 14504
rect 14608 14492 14614 14544
rect 19352 14532 19380 14572
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 26050 14560 26056 14612
rect 26108 14600 26114 14612
rect 26329 14603 26387 14609
rect 26329 14600 26341 14603
rect 26108 14572 26341 14600
rect 26108 14560 26114 14572
rect 26329 14569 26341 14572
rect 26375 14569 26387 14603
rect 26329 14563 26387 14569
rect 28399 14603 28457 14609
rect 28399 14569 28411 14603
rect 28445 14600 28457 14603
rect 29270 14600 29276 14612
rect 28445 14572 29276 14600
rect 28445 14569 28457 14572
rect 28399 14563 28457 14569
rect 29270 14560 29276 14572
rect 29328 14560 29334 14612
rect 30190 14560 30196 14612
rect 30248 14600 30254 14612
rect 30929 14603 30987 14609
rect 30929 14600 30941 14603
rect 30248 14572 30941 14600
rect 30248 14560 30254 14572
rect 30929 14569 30941 14572
rect 30975 14569 30987 14603
rect 30929 14563 30987 14569
rect 36630 14560 36636 14612
rect 36688 14600 36694 14612
rect 38654 14600 38660 14612
rect 36688 14572 38660 14600
rect 36688 14560 36694 14572
rect 38654 14560 38660 14572
rect 38712 14560 38718 14612
rect 39022 14560 39028 14612
rect 39080 14600 39086 14612
rect 47581 14603 47639 14609
rect 39080 14572 47440 14600
rect 39080 14560 39086 14572
rect 24578 14532 24584 14544
rect 17420 14504 19380 14532
rect 19444 14504 24584 14532
rect 7926 14464 7932 14476
rect 7887 14436 7932 14464
rect 7926 14424 7932 14436
rect 7984 14424 7990 14476
rect 10594 14464 10600 14476
rect 8036 14436 10600 14464
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14396 6883 14399
rect 7006 14396 7012 14408
rect 6871 14368 7012 14396
rect 6871 14365 6883 14368
rect 6825 14359 6883 14365
rect 7006 14356 7012 14368
rect 7064 14356 7070 14408
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14396 7159 14399
rect 7374 14396 7380 14408
rect 7147 14368 7380 14396
rect 7147 14365 7159 14368
rect 7101 14359 7159 14365
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 7834 14356 7840 14408
rect 7892 14396 7898 14408
rect 8036 14405 8064 14436
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 16577 14467 16635 14473
rect 16577 14433 16589 14467
rect 16623 14464 16635 14467
rect 17420 14464 17448 14504
rect 17586 14464 17592 14476
rect 16623 14436 17448 14464
rect 17547 14436 17592 14464
rect 16623 14433 16635 14436
rect 16577 14427 16635 14433
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 17770 14464 17776 14476
rect 17731 14436 17776 14464
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 17862 14424 17868 14476
rect 17920 14464 17926 14476
rect 19444 14464 19472 14504
rect 24578 14492 24584 14504
rect 24636 14492 24642 14544
rect 24688 14504 28994 14532
rect 17920 14436 19472 14464
rect 17920 14424 17926 14436
rect 21174 14424 21180 14476
rect 21232 14464 21238 14476
rect 24302 14464 24308 14476
rect 21232 14436 24308 14464
rect 21232 14424 21238 14436
rect 24302 14424 24308 14436
rect 24360 14424 24366 14476
rect 8021 14399 8079 14405
rect 8021 14396 8033 14399
rect 7892 14368 8033 14396
rect 7892 14356 7898 14368
rect 8021 14365 8033 14368
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8168 14368 8953 14396
rect 8168 14356 8174 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 2424 14300 2774 14328
rect 1762 14220 1768 14272
rect 1820 14260 1826 14272
rect 2424 14260 2452 14300
rect 7190 14288 7196 14340
rect 7248 14328 7254 14340
rect 7561 14331 7619 14337
rect 7561 14328 7573 14331
rect 7248 14300 7573 14328
rect 7248 14288 7254 14300
rect 7561 14297 7573 14300
rect 7607 14297 7619 14331
rect 8478 14328 8484 14340
rect 7561 14291 7619 14297
rect 7668 14300 8484 14328
rect 6638 14260 6644 14272
rect 1820 14232 2452 14260
rect 6599 14232 6644 14260
rect 1820 14220 1826 14232
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 7009 14263 7067 14269
rect 7009 14229 7021 14263
rect 7055 14260 7067 14263
rect 7668 14260 7696 14300
rect 8478 14288 8484 14300
rect 8536 14328 8542 14340
rect 9140 14328 9168 14359
rect 13538 14356 13544 14408
rect 13596 14396 13602 14408
rect 14277 14399 14335 14405
rect 14277 14396 14289 14399
rect 13596 14368 14289 14396
rect 13596 14356 13602 14368
rect 14277 14365 14289 14368
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 14550 14356 14556 14408
rect 14608 14396 14614 14408
rect 16482 14396 16488 14408
rect 14608 14368 14653 14396
rect 16443 14368 16488 14396
rect 14608 14356 14614 14368
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 16669 14399 16727 14405
rect 16669 14365 16681 14399
rect 16715 14365 16727 14399
rect 16669 14359 16727 14365
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14396 16819 14399
rect 17126 14396 17132 14408
rect 16807 14368 17132 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 16684 14328 16712 14359
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 17494 14396 17500 14408
rect 17455 14368 17500 14396
rect 17494 14356 17500 14368
rect 17552 14356 17558 14408
rect 17682 14399 17740 14405
rect 17682 14365 17694 14399
rect 17728 14396 17740 14399
rect 17728 14368 17816 14396
rect 17728 14365 17740 14368
rect 17682 14359 17740 14365
rect 17218 14328 17224 14340
rect 8536 14300 9168 14328
rect 14016 14300 16344 14328
rect 16684 14300 17224 14328
rect 8536 14288 8542 14300
rect 7055 14232 7696 14260
rect 7055 14229 7067 14232
rect 7009 14223 7067 14229
rect 7742 14220 7748 14272
rect 7800 14260 7806 14272
rect 8205 14263 8263 14269
rect 8205 14260 8217 14263
rect 7800 14232 8217 14260
rect 7800 14220 7806 14232
rect 8205 14229 8217 14232
rect 8251 14229 8263 14263
rect 8205 14223 8263 14229
rect 9309 14263 9367 14269
rect 9309 14229 9321 14263
rect 9355 14260 9367 14263
rect 9766 14260 9772 14272
rect 9355 14232 9772 14260
rect 9355 14229 9367 14232
rect 9309 14223 9367 14229
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 9950 14220 9956 14272
rect 10008 14260 10014 14272
rect 14016 14260 14044 14300
rect 16316 14269 16344 14300
rect 17218 14288 17224 14300
rect 17276 14288 17282 14340
rect 17788 14328 17816 14368
rect 22830 14356 22836 14408
rect 22888 14396 22894 14408
rect 24688 14396 24716 14504
rect 28966 14464 28994 14504
rect 34698 14492 34704 14544
rect 34756 14532 34762 14544
rect 35526 14532 35532 14544
rect 34756 14504 35532 14532
rect 34756 14492 34762 14504
rect 35526 14492 35532 14504
rect 35584 14492 35590 14544
rect 36817 14535 36875 14541
rect 36817 14501 36829 14535
rect 36863 14532 36875 14535
rect 37734 14532 37740 14544
rect 36863 14504 37740 14532
rect 36863 14501 36875 14504
rect 36817 14495 36875 14501
rect 37734 14492 37740 14504
rect 37792 14492 37798 14544
rect 41690 14532 41696 14544
rect 41651 14504 41696 14532
rect 41690 14492 41696 14504
rect 41748 14492 41754 14544
rect 28966 14436 29685 14464
rect 22888 14368 24716 14396
rect 22888 14356 22894 14368
rect 25682 14356 25688 14408
rect 25740 14396 25746 14408
rect 25961 14399 26019 14405
rect 25961 14396 25973 14399
rect 25740 14368 25973 14396
rect 25740 14356 25746 14368
rect 25961 14365 25973 14368
rect 26007 14396 26019 14399
rect 26878 14396 26884 14408
rect 26007 14368 26884 14396
rect 26007 14365 26019 14368
rect 25961 14359 26019 14365
rect 26878 14356 26884 14368
rect 26936 14356 26942 14408
rect 28166 14396 28172 14408
rect 28127 14368 28172 14396
rect 28166 14356 28172 14368
rect 28224 14356 28230 14408
rect 29454 14356 29460 14408
rect 29512 14396 29518 14408
rect 29549 14399 29607 14405
rect 29549 14396 29561 14399
rect 29512 14368 29561 14396
rect 29512 14356 29518 14368
rect 29549 14365 29561 14368
rect 29595 14365 29607 14399
rect 29549 14359 29607 14365
rect 20622 14328 20628 14340
rect 17788 14300 20628 14328
rect 20622 14288 20628 14300
rect 20680 14288 20686 14340
rect 24394 14288 24400 14340
rect 24452 14328 24458 14340
rect 26145 14331 26203 14337
rect 26145 14328 26157 14331
rect 24452 14300 26157 14328
rect 24452 14288 24458 14300
rect 26145 14297 26157 14300
rect 26191 14328 26203 14331
rect 27154 14328 27160 14340
rect 26191 14300 27160 14328
rect 26191 14297 26203 14300
rect 26145 14291 26203 14297
rect 27154 14288 27160 14300
rect 27212 14288 27218 14340
rect 10008 14232 14044 14260
rect 16301 14263 16359 14269
rect 10008 14220 10014 14232
rect 16301 14229 16313 14263
rect 16347 14229 16359 14263
rect 16301 14223 16359 14229
rect 16758 14220 16764 14272
rect 16816 14260 16822 14272
rect 20070 14260 20076 14272
rect 16816 14232 20076 14260
rect 16816 14220 16822 14232
rect 20070 14220 20076 14232
rect 20128 14220 20134 14272
rect 29564 14260 29592 14359
rect 29657 14328 29685 14436
rect 37550 14424 37556 14476
rect 37608 14464 37614 14476
rect 37921 14467 37979 14473
rect 37921 14464 37933 14467
rect 37608 14436 37933 14464
rect 37608 14424 37614 14436
rect 37921 14433 37933 14436
rect 37967 14433 37979 14467
rect 41598 14464 41604 14476
rect 37921 14427 37979 14433
rect 38948 14436 41604 14464
rect 29822 14405 29828 14408
rect 29816 14396 29828 14405
rect 29783 14368 29828 14396
rect 29816 14359 29828 14368
rect 29822 14356 29828 14359
rect 29880 14356 29886 14408
rect 33318 14356 33324 14408
rect 33376 14396 33382 14408
rect 37826 14396 37832 14408
rect 33376 14368 37832 14396
rect 33376 14356 33382 14368
rect 37826 14356 37832 14368
rect 37884 14356 37890 14408
rect 38188 14399 38246 14405
rect 38188 14365 38200 14399
rect 38234 14396 38246 14399
rect 38470 14396 38476 14408
rect 38234 14368 38476 14396
rect 38234 14365 38246 14368
rect 38188 14359 38246 14365
rect 38470 14356 38476 14368
rect 38528 14356 38534 14408
rect 35345 14331 35403 14337
rect 35345 14328 35357 14331
rect 29657 14300 35357 14328
rect 35345 14297 35357 14300
rect 35391 14328 35403 14331
rect 36354 14328 36360 14340
rect 35391 14300 36360 14328
rect 35391 14297 35403 14300
rect 35345 14291 35403 14297
rect 36354 14288 36360 14300
rect 36412 14288 36418 14340
rect 36538 14328 36544 14340
rect 36499 14300 36544 14328
rect 36538 14288 36544 14300
rect 36596 14288 36602 14340
rect 36722 14288 36728 14340
rect 36780 14328 36786 14340
rect 38948 14328 38976 14436
rect 41598 14424 41604 14436
rect 41656 14464 41662 14476
rect 42705 14467 42763 14473
rect 42705 14464 42717 14467
rect 41656 14436 42717 14464
rect 41656 14424 41662 14436
rect 42705 14433 42717 14436
rect 42751 14433 42763 14467
rect 42705 14427 42763 14433
rect 47412 14464 47440 14572
rect 47581 14569 47593 14603
rect 47627 14569 47639 14603
rect 47581 14563 47639 14569
rect 47765 14603 47823 14609
rect 47765 14569 47777 14603
rect 47811 14600 47823 14603
rect 48038 14600 48044 14612
rect 47811 14572 48044 14600
rect 47811 14569 47823 14572
rect 47765 14563 47823 14569
rect 47596 14532 47624 14563
rect 48038 14560 48044 14572
rect 48096 14560 48102 14612
rect 51074 14600 51080 14612
rect 48700 14572 51080 14600
rect 48593 14535 48651 14541
rect 48593 14532 48605 14535
rect 47596 14504 48605 14532
rect 48593 14501 48605 14504
rect 48639 14501 48651 14535
rect 48593 14495 48651 14501
rect 48700 14464 48728 14572
rect 51074 14560 51080 14572
rect 51132 14560 51138 14612
rect 52181 14603 52239 14609
rect 52181 14569 52193 14603
rect 52227 14600 52239 14603
rect 53190 14600 53196 14612
rect 52227 14572 53196 14600
rect 52227 14569 52239 14572
rect 52181 14563 52239 14569
rect 53190 14560 53196 14572
rect 53248 14560 53254 14612
rect 55214 14560 55220 14612
rect 55272 14600 55278 14612
rect 55401 14603 55459 14609
rect 55401 14600 55413 14603
rect 55272 14572 55413 14600
rect 55272 14560 55278 14572
rect 55401 14569 55413 14572
rect 55447 14569 55459 14603
rect 55401 14563 55459 14569
rect 55493 14603 55551 14609
rect 55493 14569 55505 14603
rect 55539 14600 55551 14603
rect 55674 14600 55680 14612
rect 55539 14572 55680 14600
rect 55539 14569 55551 14572
rect 55493 14563 55551 14569
rect 55674 14560 55680 14572
rect 55732 14560 55738 14612
rect 50798 14464 50804 14476
rect 47412 14436 48728 14464
rect 50759 14436 50804 14464
rect 41506 14356 41512 14408
rect 41564 14396 41570 14408
rect 41693 14399 41751 14405
rect 41693 14396 41705 14399
rect 41564 14368 41705 14396
rect 41564 14356 41570 14368
rect 41693 14365 41705 14368
rect 41739 14365 41751 14399
rect 41693 14359 41751 14365
rect 41969 14399 42027 14405
rect 41969 14365 41981 14399
rect 42015 14396 42027 14399
rect 42242 14396 42248 14408
rect 42015 14368 42248 14396
rect 42015 14365 42027 14368
rect 41969 14359 42027 14365
rect 42242 14356 42248 14368
rect 42300 14356 42306 14408
rect 36780 14300 38976 14328
rect 42521 14331 42579 14337
rect 36780 14288 36786 14300
rect 42521 14297 42533 14331
rect 42567 14328 42579 14331
rect 42794 14328 42800 14340
rect 42567 14300 42800 14328
rect 42567 14297 42579 14300
rect 42521 14291 42579 14297
rect 42794 14288 42800 14300
rect 42852 14288 42858 14340
rect 47412 14337 47440 14436
rect 50798 14424 50804 14436
rect 50856 14424 50862 14476
rect 55582 14464 55588 14476
rect 55543 14436 55588 14464
rect 55582 14424 55588 14436
rect 55640 14424 55646 14476
rect 48225 14399 48283 14405
rect 48225 14365 48237 14399
rect 48271 14396 48283 14399
rect 49050 14396 49056 14408
rect 48271 14368 49056 14396
rect 48271 14365 48283 14368
rect 48225 14359 48283 14365
rect 49050 14356 49056 14368
rect 49108 14356 49114 14408
rect 49237 14399 49295 14405
rect 49237 14365 49249 14399
rect 49283 14365 49295 14399
rect 49237 14359 49295 14365
rect 47397 14331 47455 14337
rect 47397 14297 47409 14331
rect 47443 14297 47455 14331
rect 47397 14291 47455 14297
rect 48409 14331 48467 14337
rect 48409 14297 48421 14331
rect 48455 14328 48467 14331
rect 48498 14328 48504 14340
rect 48455 14300 48504 14328
rect 48455 14297 48467 14300
rect 48409 14291 48467 14297
rect 48498 14288 48504 14300
rect 48556 14328 48562 14340
rect 48958 14328 48964 14340
rect 48556 14300 48964 14328
rect 48556 14288 48562 14300
rect 48958 14288 48964 14300
rect 49016 14328 49022 14340
rect 49252 14328 49280 14359
rect 50890 14356 50896 14408
rect 50948 14396 50954 14408
rect 51057 14399 51115 14405
rect 51057 14396 51069 14399
rect 50948 14368 51069 14396
rect 50948 14356 50954 14368
rect 51057 14365 51069 14368
rect 51103 14365 51115 14399
rect 51057 14359 51115 14365
rect 55030 14356 55036 14408
rect 55088 14396 55094 14408
rect 55309 14399 55367 14405
rect 55309 14396 55321 14399
rect 55088 14368 55321 14396
rect 55088 14356 55094 14368
rect 55309 14365 55321 14368
rect 55355 14365 55367 14399
rect 55309 14359 55367 14365
rect 49016 14300 49280 14328
rect 49016 14288 49022 14300
rect 32122 14260 32128 14272
rect 29564 14232 32128 14260
rect 32122 14220 32128 14232
rect 32180 14260 32186 14272
rect 32950 14260 32956 14272
rect 32180 14232 32956 14260
rect 32180 14220 32186 14232
rect 32950 14220 32956 14232
rect 33008 14220 33014 14272
rect 37734 14220 37740 14272
rect 37792 14260 37798 14272
rect 39022 14260 39028 14272
rect 37792 14232 39028 14260
rect 37792 14220 37798 14232
rect 39022 14220 39028 14232
rect 39080 14220 39086 14272
rect 39301 14263 39359 14269
rect 39301 14229 39313 14263
rect 39347 14260 39359 14263
rect 40402 14260 40408 14272
rect 39347 14232 40408 14260
rect 39347 14229 39359 14232
rect 39301 14223 39359 14229
rect 40402 14220 40408 14232
rect 40460 14220 40466 14272
rect 41874 14260 41880 14272
rect 41835 14232 41880 14260
rect 41874 14220 41880 14232
rect 41932 14220 41938 14272
rect 47607 14263 47665 14269
rect 47607 14229 47619 14263
rect 47653 14260 47665 14263
rect 47854 14260 47860 14272
rect 47653 14232 47860 14260
rect 47653 14229 47665 14232
rect 47607 14223 47665 14229
rect 47854 14220 47860 14232
rect 47912 14260 47918 14272
rect 49145 14263 49203 14269
rect 49145 14260 49157 14263
rect 47912 14232 49157 14260
rect 47912 14220 47918 14232
rect 49145 14229 49157 14232
rect 49191 14229 49203 14263
rect 49145 14223 49203 14229
rect 51902 14220 51908 14272
rect 51960 14260 51966 14272
rect 54202 14260 54208 14272
rect 51960 14232 54208 14260
rect 51960 14220 51966 14232
rect 54202 14220 54208 14232
rect 54260 14220 54266 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 2314 14056 2320 14068
rect 2275 14028 2320 14056
rect 2314 14016 2320 14028
rect 2372 14016 2378 14068
rect 2682 14056 2688 14068
rect 2643 14028 2688 14056
rect 2682 14016 2688 14028
rect 2740 14016 2746 14068
rect 7282 14016 7288 14068
rect 7340 14056 7346 14068
rect 14461 14059 14519 14065
rect 7340 14028 14412 14056
rect 7340 14016 7346 14028
rect 7742 13988 7748 14000
rect 2516 13960 7604 13988
rect 7703 13960 7748 13988
rect 2516 13929 2544 13960
rect 1397 13923 1455 13929
rect 1397 13889 1409 13923
rect 1443 13889 1455 13923
rect 1397 13883 1455 13889
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13889 2559 13923
rect 2501 13883 2559 13889
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13920 2835 13923
rect 2866 13920 2872 13932
rect 2823 13892 2872 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 1412 13852 1440 13883
rect 2866 13880 2872 13892
rect 2924 13920 2930 13932
rect 3970 13920 3976 13932
rect 2924 13892 3976 13920
rect 2924 13880 2930 13892
rect 3970 13880 3976 13892
rect 4028 13880 4034 13932
rect 7576 13920 7604 13960
rect 7742 13948 7748 13960
rect 7800 13948 7806 14000
rect 7926 13948 7932 14000
rect 7984 13988 7990 14000
rect 8202 13988 8208 14000
rect 7984 13960 8208 13988
rect 7984 13948 7990 13960
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 9766 13988 9772 14000
rect 9727 13960 9772 13988
rect 9766 13948 9772 13960
rect 9824 13948 9830 14000
rect 12066 13988 12072 14000
rect 9876 13960 12072 13988
rect 9876 13920 9904 13960
rect 12066 13948 12072 13960
rect 12124 13948 12130 14000
rect 14093 13991 14151 13997
rect 14093 13957 14105 13991
rect 14139 13957 14151 13991
rect 14093 13951 14151 13957
rect 7576 13892 9904 13920
rect 10042 13880 10048 13932
rect 10100 13920 10106 13932
rect 10686 13920 10692 13932
rect 10100 13892 10692 13920
rect 10100 13880 10106 13892
rect 10686 13880 10692 13892
rect 10744 13920 10750 13932
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 10744 13892 10793 13920
rect 10744 13880 10750 13892
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 14108 13920 14136 13951
rect 14274 13948 14280 14000
rect 14332 13997 14338 14000
rect 14332 13991 14351 13997
rect 14339 13957 14351 13991
rect 14384 13988 14412 14028
rect 14461 14025 14473 14059
rect 14507 14056 14519 14059
rect 14550 14056 14556 14068
rect 14507 14028 14556 14056
rect 14507 14025 14519 14028
rect 14461 14019 14519 14025
rect 14550 14016 14556 14028
rect 14608 14016 14614 14068
rect 16482 14016 16488 14068
rect 16540 14056 16546 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 16540 14028 17693 14056
rect 16540 14016 16546 14028
rect 17681 14025 17693 14028
rect 17727 14025 17739 14059
rect 17681 14019 17739 14025
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 20809 14059 20867 14065
rect 20809 14056 20821 14059
rect 20680 14028 20821 14056
rect 20680 14016 20686 14028
rect 20809 14025 20821 14028
rect 20855 14025 20867 14059
rect 20809 14019 20867 14025
rect 23293 14059 23351 14065
rect 23293 14025 23305 14059
rect 23339 14056 23351 14059
rect 23658 14056 23664 14068
rect 23339 14028 23664 14056
rect 23339 14025 23351 14028
rect 23293 14019 23351 14025
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 23779 14059 23837 14065
rect 23779 14025 23791 14059
rect 23825 14056 23837 14059
rect 24597 14059 24655 14065
rect 24597 14056 24609 14059
rect 23825 14028 24609 14056
rect 23825 14025 23837 14028
rect 23779 14019 23837 14025
rect 24597 14025 24609 14028
rect 24643 14056 24655 14059
rect 24762 14056 24768 14068
rect 24643 14028 24768 14056
rect 24643 14025 24655 14028
rect 24597 14019 24655 14025
rect 24762 14016 24768 14028
rect 24820 14016 24826 14068
rect 25314 14016 25320 14068
rect 25372 14056 25378 14068
rect 26053 14059 26111 14065
rect 26053 14056 26065 14059
rect 25372 14028 26065 14056
rect 25372 14016 25378 14028
rect 26053 14025 26065 14028
rect 26099 14025 26111 14059
rect 26053 14019 26111 14025
rect 26418 14016 26424 14068
rect 26476 14056 26482 14068
rect 30466 14056 30472 14068
rect 26476 14028 30472 14056
rect 26476 14016 26482 14028
rect 30466 14016 30472 14028
rect 30524 14016 30530 14068
rect 34054 14016 34060 14068
rect 34112 14056 34118 14068
rect 35529 14059 35587 14065
rect 35529 14056 35541 14059
rect 34112 14028 35541 14056
rect 34112 14016 34118 14028
rect 35529 14025 35541 14028
rect 35575 14025 35587 14059
rect 36446 14056 36452 14068
rect 36407 14028 36452 14056
rect 35529 14019 35587 14025
rect 36446 14016 36452 14028
rect 36504 14016 36510 14068
rect 37826 14056 37832 14068
rect 37787 14028 37832 14056
rect 37826 14016 37832 14028
rect 37884 14016 37890 14068
rect 38562 14016 38568 14068
rect 38620 14056 38626 14068
rect 38838 14056 38844 14068
rect 38620 14028 38844 14056
rect 38620 14016 38626 14028
rect 38838 14016 38844 14028
rect 38896 14056 38902 14068
rect 41414 14056 41420 14068
rect 38896 14028 41420 14056
rect 38896 14016 38902 14028
rect 41414 14016 41420 14028
rect 41472 14056 41478 14068
rect 41874 14056 41880 14068
rect 41472 14028 41880 14056
rect 41472 14016 41478 14028
rect 41874 14016 41880 14028
rect 41932 14016 41938 14068
rect 52178 14016 52184 14068
rect 52236 14056 52242 14068
rect 53101 14059 53159 14065
rect 53101 14056 53113 14059
rect 52236 14028 53113 14056
rect 52236 14016 52242 14028
rect 53101 14025 53113 14028
rect 53147 14025 53159 14059
rect 54018 14056 54024 14068
rect 53979 14028 54024 14056
rect 53101 14019 53159 14025
rect 54018 14016 54024 14028
rect 54076 14016 54082 14068
rect 54202 14056 54208 14068
rect 54163 14028 54208 14056
rect 54202 14016 54208 14028
rect 54260 14016 54266 14068
rect 16758 13988 16764 14000
rect 14384 13960 16764 13988
rect 14332 13951 14351 13957
rect 14332 13948 14338 13951
rect 16758 13948 16764 13960
rect 16816 13948 16822 14000
rect 22462 13988 22468 14000
rect 16960 13960 22468 13988
rect 14550 13920 14556 13932
rect 14108 13892 14556 13920
rect 10781 13883 10839 13889
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 16960 13929 16988 13960
rect 22462 13948 22468 13960
rect 22520 13948 22526 14000
rect 23474 13948 23480 14000
rect 23532 13988 23538 14000
rect 23569 13991 23627 13997
rect 23569 13988 23581 13991
rect 23532 13960 23581 13988
rect 23532 13948 23538 13960
rect 23569 13957 23581 13960
rect 23615 13988 23627 13991
rect 24397 13991 24455 13997
rect 24397 13988 24409 13991
rect 23615 13960 24409 13988
rect 23615 13957 23627 13960
rect 23569 13951 23627 13957
rect 24397 13957 24409 13960
rect 24443 13957 24455 13991
rect 24397 13951 24455 13957
rect 16945 13923 17003 13929
rect 16945 13889 16957 13923
rect 16991 13889 17003 13923
rect 16945 13883 17003 13889
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17218 13920 17224 13932
rect 17083 13892 17224 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 17494 13880 17500 13932
rect 17552 13920 17558 13932
rect 17865 13923 17923 13929
rect 17865 13920 17877 13923
rect 17552 13892 17877 13920
rect 17552 13880 17558 13892
rect 17865 13889 17877 13892
rect 17911 13889 17923 13923
rect 17865 13883 17923 13889
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 18506 13920 18512 13932
rect 18095 13892 18512 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 18506 13880 18512 13892
rect 18564 13880 18570 13932
rect 19426 13920 19432 13932
rect 19387 13892 19432 13920
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 19696 13923 19754 13929
rect 19696 13889 19708 13923
rect 19742 13920 19754 13923
rect 19978 13920 19984 13932
rect 19742 13892 19984 13920
rect 19742 13889 19754 13892
rect 19696 13883 19754 13889
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 22186 13880 22192 13932
rect 22244 13920 22250 13932
rect 22244 13892 24256 13920
rect 22244 13880 22250 13892
rect 4614 13852 4620 13864
rect 1412 13824 4620 13852
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 6696 13824 8125 13852
rect 6696 13812 6702 13824
rect 8113 13821 8125 13824
rect 8159 13821 8171 13855
rect 8113 13815 8171 13821
rect 8481 13855 8539 13861
rect 8481 13821 8493 13855
rect 8527 13852 8539 13855
rect 8527 13824 10548 13852
rect 8527 13821 8539 13824
rect 8481 13815 8539 13821
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 7742 13784 7748 13796
rect 7340 13756 7748 13784
rect 7340 13744 7346 13756
rect 7742 13744 7748 13756
rect 7800 13744 7806 13796
rect 8018 13784 8024 13796
rect 7979 13756 8024 13784
rect 8018 13744 8024 13756
rect 8076 13744 8082 13796
rect 9950 13784 9956 13796
rect 9911 13756 9956 13784
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 10520 13784 10548 13824
rect 10594 13812 10600 13864
rect 10652 13852 10658 13864
rect 10965 13855 11023 13861
rect 10652 13824 10697 13852
rect 10652 13812 10658 13824
rect 10965 13821 10977 13855
rect 11011 13852 11023 13855
rect 11422 13852 11428 13864
rect 11011 13824 11428 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 12158 13852 12164 13864
rect 11532 13824 12164 13852
rect 11532 13784 11560 13824
rect 12158 13812 12164 13824
rect 12216 13812 12222 13864
rect 16666 13852 16672 13864
rect 16627 13824 16672 13852
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 16850 13852 16856 13864
rect 16811 13824 16856 13852
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 17126 13812 17132 13864
rect 17184 13852 17190 13864
rect 17954 13852 17960 13864
rect 17184 13824 17229 13852
rect 17915 13824 17960 13852
rect 17184 13812 17190 13824
rect 17954 13812 17960 13824
rect 18012 13812 18018 13864
rect 18141 13855 18199 13861
rect 18141 13821 18153 13855
rect 18187 13821 18199 13855
rect 18141 13815 18199 13821
rect 10520 13756 11560 13784
rect 16758 13744 16764 13796
rect 16816 13784 16822 13796
rect 16942 13784 16948 13796
rect 16816 13756 16948 13784
rect 16816 13744 16822 13756
rect 16942 13744 16948 13756
rect 17000 13744 17006 13796
rect 17770 13744 17776 13796
rect 17828 13784 17834 13796
rect 18046 13784 18052 13796
rect 17828 13756 18052 13784
rect 17828 13744 17834 13756
rect 18046 13744 18052 13756
rect 18104 13784 18110 13796
rect 18156 13784 18184 13815
rect 20990 13812 20996 13864
rect 21048 13852 21054 13864
rect 23014 13852 23020 13864
rect 21048 13824 23020 13852
rect 21048 13812 21054 13824
rect 23014 13812 23020 13824
rect 23072 13812 23078 13864
rect 23842 13812 23848 13864
rect 23900 13852 23906 13864
rect 24118 13852 24124 13864
rect 23900 13824 24124 13852
rect 23900 13812 23906 13824
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 18104 13756 18184 13784
rect 23860 13784 23888 13812
rect 23937 13787 23995 13793
rect 23937 13784 23949 13787
rect 23860 13756 23949 13784
rect 18104 13744 18110 13756
rect 23937 13753 23949 13756
rect 23983 13753 23995 13787
rect 24228 13784 24256 13892
rect 24670 13880 24676 13932
rect 24728 13920 24734 13932
rect 25332 13920 25360 14016
rect 31570 13948 31576 14000
rect 31628 13988 31634 14000
rect 31628 13960 36308 13988
rect 31628 13948 31634 13960
rect 25682 13920 25688 13932
rect 24728 13892 25360 13920
rect 25643 13892 25688 13920
rect 24728 13880 24734 13892
rect 25682 13880 25688 13892
rect 25740 13880 25746 13932
rect 32950 13880 32956 13932
rect 33008 13920 33014 13932
rect 33229 13923 33287 13929
rect 33229 13920 33241 13923
rect 33008 13892 33241 13920
rect 33008 13880 33014 13892
rect 33229 13889 33241 13892
rect 33275 13889 33287 13923
rect 33229 13883 33287 13889
rect 33318 13880 33324 13932
rect 33376 13920 33382 13932
rect 36280 13929 36308 13960
rect 36354 13948 36360 14000
rect 36412 13988 36418 14000
rect 37737 13991 37795 13997
rect 37737 13988 37749 13991
rect 36412 13960 37749 13988
rect 36412 13948 36418 13960
rect 37737 13957 37749 13960
rect 37783 13988 37795 13991
rect 38378 13988 38384 14000
rect 37783 13960 38384 13988
rect 37783 13957 37795 13960
rect 37737 13951 37795 13957
rect 38378 13948 38384 13960
rect 38436 13948 38442 14000
rect 38470 13948 38476 14000
rect 38528 13988 38534 14000
rect 52733 13991 52791 13997
rect 38528 13960 45692 13988
rect 38528 13948 38534 13960
rect 33485 13923 33543 13929
rect 33485 13920 33497 13923
rect 33376 13892 33497 13920
rect 33376 13880 33382 13892
rect 33485 13889 33497 13892
rect 33531 13889 33543 13923
rect 33485 13883 33543 13889
rect 35345 13923 35403 13929
rect 35345 13889 35357 13923
rect 35391 13920 35403 13923
rect 36265 13923 36323 13929
rect 35391 13892 36032 13920
rect 35391 13889 35403 13892
rect 35345 13883 35403 13889
rect 24765 13787 24823 13793
rect 24765 13784 24777 13787
rect 24228 13756 24777 13784
rect 23937 13747 23995 13753
rect 24765 13753 24777 13756
rect 24811 13784 24823 13787
rect 25682 13784 25688 13796
rect 24811 13756 25688 13784
rect 24811 13753 24823 13756
rect 24765 13747 24823 13753
rect 25682 13744 25688 13756
rect 25740 13744 25746 13796
rect 34606 13784 34612 13796
rect 34567 13756 34612 13784
rect 34606 13744 34612 13756
rect 34664 13744 34670 13796
rect 36004 13784 36032 13892
rect 36265 13889 36277 13923
rect 36311 13889 36323 13923
rect 38562 13920 38568 13932
rect 38523 13892 38568 13920
rect 36265 13883 36323 13889
rect 38562 13880 38568 13892
rect 38620 13880 38626 13932
rect 38746 13880 38752 13932
rect 38804 13920 38810 13932
rect 40402 13920 40408 13932
rect 38804 13892 38849 13920
rect 40363 13892 40408 13920
rect 38804 13880 38810 13892
rect 40402 13880 40408 13892
rect 40460 13880 40466 13932
rect 41690 13880 41696 13932
rect 41748 13920 41754 13932
rect 45664 13929 45692 13960
rect 52733 13957 52745 13991
rect 52779 13988 52791 13991
rect 53190 13988 53196 14000
rect 52779 13960 53196 13988
rect 52779 13957 52791 13960
rect 52733 13951 52791 13957
rect 53190 13948 53196 13960
rect 53248 13948 53254 14000
rect 53834 13988 53840 14000
rect 53795 13960 53840 13988
rect 53834 13948 53840 13960
rect 53892 13948 53898 14000
rect 42869 13923 42927 13929
rect 42869 13920 42881 13923
rect 41748 13892 42881 13920
rect 41748 13880 41754 13892
rect 42869 13889 42881 13892
rect 42915 13889 42927 13923
rect 42869 13883 42927 13889
rect 45649 13923 45707 13929
rect 45649 13889 45661 13923
rect 45695 13889 45707 13923
rect 45649 13883 45707 13889
rect 45833 13923 45891 13929
rect 45833 13889 45845 13923
rect 45879 13920 45891 13923
rect 45879 13892 46980 13920
rect 45879 13889 45891 13892
rect 45833 13883 45891 13889
rect 36081 13855 36139 13861
rect 36081 13821 36093 13855
rect 36127 13852 36139 13855
rect 36170 13852 36176 13864
rect 36127 13824 36176 13852
rect 36127 13821 36139 13824
rect 36081 13815 36139 13821
rect 36170 13812 36176 13824
rect 36228 13852 36234 13864
rect 36722 13852 36728 13864
rect 36228 13824 36728 13852
rect 36228 13812 36234 13824
rect 36722 13812 36728 13824
rect 36780 13812 36786 13864
rect 36906 13812 36912 13864
rect 36964 13852 36970 13864
rect 38657 13855 38715 13861
rect 38657 13852 38669 13855
rect 36964 13824 38669 13852
rect 36964 13812 36970 13824
rect 38657 13821 38669 13824
rect 38703 13821 38715 13855
rect 38657 13815 38715 13821
rect 40310 13812 40316 13864
rect 40368 13852 40374 13864
rect 40681 13855 40739 13861
rect 40681 13852 40693 13855
rect 40368 13824 40693 13852
rect 40368 13812 40374 13824
rect 40681 13821 40693 13824
rect 40727 13852 40739 13855
rect 40770 13852 40776 13864
rect 40727 13824 40776 13852
rect 40727 13821 40739 13824
rect 40681 13815 40739 13821
rect 40770 13812 40776 13824
rect 40828 13812 40834 13864
rect 42518 13812 42524 13864
rect 42576 13852 42582 13864
rect 42613 13855 42671 13861
rect 42613 13852 42625 13855
rect 42576 13824 42625 13852
rect 42576 13812 42582 13824
rect 42613 13821 42625 13824
rect 42659 13821 42671 13855
rect 42613 13815 42671 13821
rect 36630 13784 36636 13796
rect 36004 13756 36636 13784
rect 36630 13744 36636 13756
rect 36688 13744 36694 13796
rect 46952 13784 46980 13892
rect 47394 13880 47400 13932
rect 47452 13920 47458 13932
rect 47765 13923 47823 13929
rect 47765 13920 47777 13923
rect 47452 13892 47777 13920
rect 47452 13880 47458 13892
rect 47765 13889 47777 13892
rect 47811 13889 47823 13923
rect 47765 13883 47823 13889
rect 52917 13923 52975 13929
rect 52917 13889 52929 13923
rect 52963 13889 52975 13923
rect 52917 13883 52975 13889
rect 53009 13923 53067 13929
rect 53009 13889 53021 13923
rect 53055 13920 53067 13923
rect 54110 13920 54116 13932
rect 53055 13892 53972 13920
rect 54071 13892 54116 13920
rect 53055 13889 53067 13892
rect 53009 13883 53067 13889
rect 47854 13852 47860 13864
rect 47815 13824 47860 13852
rect 47854 13812 47860 13824
rect 47912 13812 47918 13864
rect 52932 13852 52960 13883
rect 53098 13852 53104 13864
rect 52932 13824 53104 13852
rect 53098 13812 53104 13824
rect 53156 13812 53162 13864
rect 53944 13852 53972 13892
rect 54110 13880 54116 13892
rect 54168 13880 54174 13932
rect 54570 13852 54576 13864
rect 53944 13824 54576 13852
rect 54570 13812 54576 13824
rect 54628 13812 54634 13864
rect 48133 13787 48191 13793
rect 48133 13784 48145 13787
rect 46952 13756 48145 13784
rect 48133 13753 48145 13756
rect 48179 13753 48191 13787
rect 48133 13747 48191 13753
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 7910 13719 7968 13725
rect 7910 13716 7922 13719
rect 6972 13688 7922 13716
rect 6972 13676 6978 13688
rect 7910 13685 7922 13688
rect 7956 13716 7968 13719
rect 10134 13716 10140 13728
rect 7956 13688 10140 13716
rect 7956 13685 7968 13688
rect 7910 13679 7968 13685
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 14277 13719 14335 13725
rect 14277 13685 14289 13719
rect 14323 13716 14335 13719
rect 14734 13716 14740 13728
rect 14323 13688 14740 13716
rect 14323 13685 14335 13688
rect 14277 13679 14335 13685
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 18138 13676 18144 13728
rect 18196 13716 18202 13728
rect 19426 13716 19432 13728
rect 18196 13688 19432 13716
rect 18196 13676 18202 13688
rect 19426 13676 19432 13688
rect 19484 13676 19490 13728
rect 23658 13676 23664 13728
rect 23716 13716 23722 13728
rect 23753 13719 23811 13725
rect 23753 13716 23765 13719
rect 23716 13688 23765 13716
rect 23716 13676 23722 13688
rect 23753 13685 23765 13688
rect 23799 13685 23811 13719
rect 23753 13679 23811 13685
rect 24302 13676 24308 13728
rect 24360 13716 24366 13728
rect 24578 13716 24584 13728
rect 24360 13688 24584 13716
rect 24360 13676 24366 13688
rect 24578 13676 24584 13688
rect 24636 13676 24642 13728
rect 25590 13676 25596 13728
rect 25648 13716 25654 13728
rect 26053 13719 26111 13725
rect 26053 13716 26065 13719
rect 25648 13688 26065 13716
rect 25648 13676 25654 13688
rect 26053 13685 26065 13688
rect 26099 13685 26111 13719
rect 26234 13716 26240 13728
rect 26195 13688 26240 13716
rect 26053 13679 26111 13685
rect 26234 13676 26240 13688
rect 26292 13676 26298 13728
rect 30374 13676 30380 13728
rect 30432 13716 30438 13728
rect 37918 13716 37924 13728
rect 30432 13688 37924 13716
rect 30432 13676 30438 13688
rect 37918 13676 37924 13688
rect 37976 13676 37982 13728
rect 42794 13676 42800 13728
rect 42852 13716 42858 13728
rect 43993 13719 44051 13725
rect 43993 13716 44005 13719
rect 42852 13688 44005 13716
rect 42852 13676 42858 13688
rect 43993 13685 44005 13688
rect 44039 13685 44051 13719
rect 43993 13679 44051 13685
rect 46017 13719 46075 13725
rect 46017 13685 46029 13719
rect 46063 13716 46075 13719
rect 46198 13716 46204 13728
rect 46063 13688 46204 13716
rect 46063 13685 46075 13688
rect 46017 13679 46075 13685
rect 46198 13676 46204 13688
rect 46256 13676 46262 13728
rect 53282 13716 53288 13728
rect 53243 13688 53288 13716
rect 53282 13676 53288 13688
rect 53340 13676 53346 13728
rect 53926 13676 53932 13728
rect 53984 13716 53990 13728
rect 54389 13719 54447 13725
rect 54389 13716 54401 13719
rect 53984 13688 54401 13716
rect 53984 13676 53990 13688
rect 54389 13685 54401 13688
rect 54435 13685 54447 13719
rect 54389 13679 54447 13685
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 6914 13512 6920 13524
rect 6875 13484 6920 13512
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7193 13515 7251 13521
rect 7193 13512 7205 13515
rect 7156 13484 7205 13512
rect 7156 13472 7162 13484
rect 7193 13481 7205 13484
rect 7239 13512 7251 13515
rect 7650 13512 7656 13524
rect 7239 13484 7656 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 8018 13472 8024 13524
rect 8076 13512 8082 13524
rect 10042 13512 10048 13524
rect 8076 13484 10048 13512
rect 8076 13472 8082 13484
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10226 13512 10232 13524
rect 10187 13484 10232 13512
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 19978 13512 19984 13524
rect 12406 13484 15056 13512
rect 19939 13484 19984 13512
rect 6638 13404 6644 13456
rect 6696 13444 6702 13456
rect 7377 13447 7435 13453
rect 7377 13444 7389 13447
rect 6696 13416 7389 13444
rect 6696 13404 6702 13416
rect 7377 13413 7389 13416
rect 7423 13413 7435 13447
rect 7377 13407 7435 13413
rect 7742 13404 7748 13456
rect 7800 13444 7806 13456
rect 8110 13444 8116 13456
rect 7800 13416 8116 13444
rect 7800 13404 7806 13416
rect 8110 13404 8116 13416
rect 8168 13444 8174 13456
rect 8205 13447 8263 13453
rect 8205 13444 8217 13447
rect 8168 13416 8217 13444
rect 8168 13404 8174 13416
rect 8205 13413 8217 13416
rect 8251 13413 8263 13447
rect 8205 13407 8263 13413
rect 9950 13404 9956 13456
rect 10008 13444 10014 13456
rect 10594 13444 10600 13456
rect 10008 13416 10600 13444
rect 10008 13404 10014 13416
rect 2590 13336 2596 13388
rect 2648 13376 2654 13388
rect 3786 13376 3792 13388
rect 2648 13348 3792 13376
rect 2648 13336 2654 13348
rect 3786 13336 3792 13348
rect 3844 13336 3850 13388
rect 7190 13336 7196 13388
rect 7248 13376 7254 13388
rect 10244 13385 10272 13416
rect 10594 13404 10600 13416
rect 10652 13444 10658 13456
rect 12406 13444 12434 13484
rect 10652 13416 12434 13444
rect 15028 13444 15056 13484
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 22094 13472 22100 13524
rect 22152 13512 22158 13524
rect 22830 13512 22836 13524
rect 22152 13484 22836 13512
rect 22152 13472 22158 13484
rect 22830 13472 22836 13484
rect 22888 13472 22894 13524
rect 23106 13512 23112 13524
rect 23019 13484 23112 13512
rect 23106 13472 23112 13484
rect 23164 13512 23170 13524
rect 23569 13515 23627 13521
rect 23569 13512 23581 13515
rect 23164 13484 23581 13512
rect 23164 13472 23170 13484
rect 23569 13481 23581 13484
rect 23615 13512 23627 13515
rect 30374 13512 30380 13524
rect 23615 13484 30380 13512
rect 23615 13481 23627 13484
rect 23569 13475 23627 13481
rect 30374 13472 30380 13484
rect 30432 13472 30438 13524
rect 30466 13472 30472 13524
rect 30524 13512 30530 13524
rect 30561 13515 30619 13521
rect 30561 13512 30573 13515
rect 30524 13484 30573 13512
rect 30524 13472 30530 13484
rect 30561 13481 30573 13484
rect 30607 13481 30619 13515
rect 33318 13512 33324 13524
rect 33279 13484 33324 13512
rect 30561 13475 30619 13481
rect 33318 13472 33324 13484
rect 33376 13472 33382 13524
rect 36541 13515 36599 13521
rect 36541 13481 36553 13515
rect 36587 13512 36599 13515
rect 36630 13512 36636 13524
rect 36587 13484 36636 13512
rect 36587 13481 36599 13484
rect 36541 13475 36599 13481
rect 36630 13472 36636 13484
rect 36688 13472 36694 13524
rect 37277 13515 37335 13521
rect 37277 13481 37289 13515
rect 37323 13512 37335 13515
rect 38010 13512 38016 13524
rect 37323 13484 38016 13512
rect 37323 13481 37335 13484
rect 37277 13475 37335 13481
rect 38010 13472 38016 13484
rect 38068 13512 38074 13524
rect 38470 13512 38476 13524
rect 38068 13484 38476 13512
rect 38068 13472 38074 13484
rect 38470 13472 38476 13484
rect 38528 13472 38534 13524
rect 41414 13512 41420 13524
rect 41375 13484 41420 13512
rect 41414 13472 41420 13484
rect 41472 13472 41478 13524
rect 42794 13512 42800 13524
rect 42755 13484 42800 13512
rect 42794 13472 42800 13484
rect 42852 13472 42858 13524
rect 50614 13472 50620 13524
rect 50672 13512 50678 13524
rect 51169 13515 51227 13521
rect 51169 13512 51181 13515
rect 50672 13484 51181 13512
rect 50672 13472 50678 13484
rect 51169 13481 51181 13484
rect 51215 13512 51227 13515
rect 54570 13512 54576 13524
rect 51215 13484 53604 13512
rect 54531 13484 54576 13512
rect 51215 13481 51227 13484
rect 51169 13475 51227 13481
rect 20438 13444 20444 13456
rect 15028 13416 20444 13444
rect 10652 13404 10658 13416
rect 20438 13404 20444 13416
rect 20496 13404 20502 13456
rect 23290 13444 23296 13456
rect 22066 13416 23296 13444
rect 10229 13379 10287 13385
rect 7248 13348 8340 13376
rect 7248 13336 7254 13348
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13308 2375 13311
rect 2774 13308 2780 13320
rect 2363 13280 2780 13308
rect 2363 13277 2375 13280
rect 2317 13271 2375 13277
rect 2774 13268 2780 13280
rect 2832 13268 2838 13320
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13308 7343 13311
rect 7558 13308 7564 13320
rect 7331 13280 7564 13308
rect 7331 13277 7343 13280
rect 7285 13271 7343 13277
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13308 7711 13311
rect 7926 13308 7932 13320
rect 7699 13280 7932 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 8018 13268 8024 13320
rect 8076 13308 8082 13320
rect 8312 13317 8340 13348
rect 10229 13345 10241 13379
rect 10275 13345 10287 13379
rect 11422 13376 11428 13388
rect 11383 13348 11428 13376
rect 10229 13339 10287 13345
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 22066 13376 22094 13416
rect 23290 13404 23296 13416
rect 23348 13444 23354 13456
rect 23753 13447 23811 13453
rect 23753 13444 23765 13447
rect 23348 13416 23765 13444
rect 23348 13404 23354 13416
rect 23753 13413 23765 13416
rect 23799 13413 23811 13447
rect 34514 13444 34520 13456
rect 23753 13407 23811 13413
rect 23860 13416 34520 13444
rect 20180 13348 22094 13376
rect 8113 13311 8171 13317
rect 8113 13308 8125 13311
rect 8076 13280 8125 13308
rect 8076 13268 8082 13280
rect 8113 13277 8125 13280
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13277 8355 13311
rect 10134 13308 10140 13320
rect 10095 13280 10140 13308
rect 8297 13271 8355 13277
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13308 11759 13311
rect 11790 13308 11796 13320
rect 11747 13280 11796 13308
rect 11747 13277 11759 13280
rect 11701 13271 11759 13277
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 12250 13268 12256 13320
rect 12308 13308 12314 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 12308 13280 14105 13308
rect 12308 13268 12314 13280
rect 14093 13277 14105 13280
rect 14139 13308 14151 13311
rect 18138 13308 18144 13320
rect 14139 13280 18144 13308
rect 14139 13277 14151 13280
rect 14093 13271 14151 13277
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 20180 13317 20208 13348
rect 22646 13336 22652 13388
rect 22704 13376 22710 13388
rect 23860 13376 23888 13416
rect 34514 13404 34520 13416
rect 34572 13404 34578 13456
rect 51353 13447 51411 13453
rect 51353 13413 51365 13447
rect 51399 13413 51411 13447
rect 51353 13407 51411 13413
rect 22704 13348 23888 13376
rect 22704 13336 22710 13348
rect 25038 13336 25044 13388
rect 25096 13376 25102 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 25096 13348 25145 13376
rect 25096 13336 25102 13348
rect 25133 13345 25145 13348
rect 25179 13376 25191 13379
rect 25406 13376 25412 13388
rect 25179 13348 25412 13376
rect 25179 13345 25191 13348
rect 25133 13339 25191 13345
rect 25406 13336 25412 13348
rect 25464 13336 25470 13388
rect 28353 13379 28411 13385
rect 28353 13345 28365 13379
rect 28399 13376 28411 13379
rect 33134 13376 33140 13388
rect 28399 13348 33140 13376
rect 28399 13345 28411 13348
rect 28353 13339 28411 13345
rect 33134 13336 33140 13348
rect 33192 13376 33198 13388
rect 33965 13379 34023 13385
rect 33192 13348 33640 13376
rect 33192 13336 33198 13348
rect 20165 13311 20223 13317
rect 20165 13277 20177 13311
rect 20211 13277 20223 13311
rect 20165 13271 20223 13277
rect 20441 13311 20499 13317
rect 20441 13277 20453 13311
rect 20487 13308 20499 13311
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 20487 13280 21281 13308
rect 20487 13277 20499 13280
rect 20441 13271 20499 13277
rect 21269 13277 21281 13280
rect 21315 13277 21327 13311
rect 21910 13308 21916 13320
rect 21871 13280 21916 13308
rect 21269 13271 21327 13277
rect 4062 13249 4068 13252
rect 4056 13203 4068 13249
rect 4120 13240 4126 13252
rect 4120 13212 4156 13240
rect 4062 13200 4068 13203
rect 4120 13200 4126 13212
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 9766 13240 9772 13252
rect 8444 13212 9772 13240
rect 8444 13200 8450 13212
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 10410 13200 10416 13252
rect 10468 13240 10474 13252
rect 10686 13240 10692 13252
rect 10468 13212 10692 13240
rect 10468 13200 10474 13212
rect 10686 13200 10692 13212
rect 10744 13200 10750 13252
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14338 13243 14396 13249
rect 14338 13240 14350 13243
rect 14240 13212 14350 13240
rect 14240 13200 14246 13212
rect 14338 13209 14350 13212
rect 14384 13209 14396 13243
rect 14338 13203 14396 13209
rect 19426 13200 19432 13252
rect 19484 13240 19490 13252
rect 20456 13240 20484 13271
rect 21910 13268 21916 13280
rect 21968 13268 21974 13320
rect 22465 13311 22523 13317
rect 22465 13277 22477 13311
rect 22511 13308 22523 13311
rect 22830 13308 22836 13320
rect 22511 13280 22836 13308
rect 22511 13277 22523 13280
rect 22465 13271 22523 13277
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 24762 13268 24768 13320
rect 24820 13308 24826 13320
rect 24857 13311 24915 13317
rect 24857 13308 24869 13311
rect 24820 13280 24869 13308
rect 24820 13268 24826 13280
rect 24857 13277 24869 13280
rect 24903 13277 24915 13311
rect 24857 13271 24915 13277
rect 25682 13268 25688 13320
rect 25740 13308 25746 13320
rect 25777 13311 25835 13317
rect 25777 13308 25789 13311
rect 25740 13280 25789 13308
rect 25740 13268 25746 13280
rect 25777 13277 25789 13280
rect 25823 13277 25835 13311
rect 25777 13271 25835 13277
rect 26145 13311 26203 13317
rect 26145 13277 26157 13311
rect 26191 13308 26203 13311
rect 26789 13311 26847 13317
rect 26789 13308 26801 13311
rect 26191 13280 26801 13308
rect 26191 13277 26203 13280
rect 26145 13271 26203 13277
rect 26789 13277 26801 13280
rect 26835 13277 26847 13311
rect 26789 13271 26847 13277
rect 27890 13268 27896 13320
rect 27948 13308 27954 13320
rect 28261 13311 28319 13317
rect 28261 13308 28273 13311
rect 27948 13280 28273 13308
rect 27948 13268 27954 13280
rect 28261 13277 28273 13280
rect 28307 13277 28319 13311
rect 28442 13308 28448 13320
rect 28403 13280 28448 13308
rect 28261 13271 28319 13277
rect 28442 13268 28448 13280
rect 28500 13268 28506 13320
rect 30374 13308 30380 13320
rect 30335 13280 30380 13308
rect 30374 13268 30380 13280
rect 30432 13308 30438 13320
rect 31846 13308 31852 13320
rect 30432 13280 31754 13308
rect 31807 13280 31852 13308
rect 30432 13268 30438 13280
rect 19484 13212 20484 13240
rect 21085 13243 21143 13249
rect 19484 13200 19490 13212
rect 21085 13209 21097 13243
rect 21131 13240 21143 13243
rect 22094 13240 22100 13252
rect 21131 13212 22100 13240
rect 21131 13209 21143 13212
rect 21085 13203 21143 13209
rect 22094 13200 22100 13212
rect 22152 13200 22158 13252
rect 23385 13243 23443 13249
rect 23385 13209 23397 13243
rect 23431 13240 23443 13243
rect 23474 13240 23480 13252
rect 23431 13212 23480 13240
rect 23431 13209 23443 13212
rect 23385 13203 23443 13209
rect 23474 13200 23480 13212
rect 23532 13200 23538 13252
rect 23601 13243 23659 13249
rect 23601 13209 23613 13243
rect 23647 13240 23659 13243
rect 24780 13240 24808 13268
rect 23647 13212 24808 13240
rect 25961 13243 26019 13249
rect 23647 13209 23659 13212
rect 23601 13203 23659 13209
rect 25961 13209 25973 13243
rect 26007 13240 26019 13243
rect 26234 13240 26240 13252
rect 26007 13212 26240 13240
rect 26007 13209 26019 13212
rect 25961 13203 26019 13209
rect 26234 13200 26240 13212
rect 26292 13200 26298 13252
rect 31726 13240 31754 13280
rect 31846 13268 31852 13280
rect 31904 13268 31910 13320
rect 33318 13268 33324 13320
rect 33376 13308 33382 13320
rect 33612 13317 33640 13348
rect 33965 13345 33977 13379
rect 34011 13376 34023 13379
rect 34054 13376 34060 13388
rect 34011 13348 34060 13376
rect 34011 13345 34023 13348
rect 33965 13339 34023 13345
rect 34054 13336 34060 13348
rect 34112 13336 34118 13388
rect 46014 13376 46020 13388
rect 45975 13348 46020 13376
rect 46014 13336 46020 13348
rect 46072 13336 46078 13388
rect 33505 13311 33563 13317
rect 33505 13308 33517 13311
rect 33376 13280 33517 13308
rect 33376 13268 33382 13280
rect 33505 13277 33517 13280
rect 33551 13277 33563 13311
rect 33505 13271 33563 13277
rect 33597 13311 33655 13317
rect 33597 13277 33609 13311
rect 33643 13277 33655 13311
rect 36357 13311 36415 13317
rect 36357 13308 36369 13311
rect 33597 13271 33655 13277
rect 33797 13280 36369 13308
rect 33797 13240 33825 13280
rect 36357 13277 36369 13280
rect 36403 13308 36415 13311
rect 36538 13308 36544 13320
rect 36403 13280 36544 13308
rect 36403 13277 36415 13280
rect 36357 13271 36415 13277
rect 36538 13268 36544 13280
rect 36596 13308 36602 13320
rect 37093 13311 37151 13317
rect 37093 13308 37105 13311
rect 36596 13280 37105 13308
rect 36596 13268 36602 13280
rect 37093 13277 37105 13280
rect 37139 13277 37151 13311
rect 37093 13271 37151 13277
rect 38654 13268 38660 13320
rect 38712 13308 38718 13320
rect 38749 13311 38807 13317
rect 38749 13308 38761 13311
rect 38712 13280 38761 13308
rect 38712 13268 38718 13280
rect 38749 13277 38761 13280
rect 38795 13277 38807 13311
rect 39022 13308 39028 13320
rect 38983 13280 39028 13308
rect 38749 13271 38807 13277
rect 39022 13268 39028 13280
rect 39080 13268 39086 13320
rect 40402 13268 40408 13320
rect 40460 13308 40466 13320
rect 41233 13311 41291 13317
rect 41233 13308 41245 13311
rect 40460 13280 41245 13308
rect 40460 13268 40466 13280
rect 41233 13277 41245 13280
rect 41279 13308 41291 13311
rect 42426 13308 42432 13320
rect 41279 13280 42432 13308
rect 41279 13277 41291 13280
rect 41233 13271 41291 13277
rect 42426 13268 42432 13280
rect 42484 13268 42490 13320
rect 42797 13311 42855 13317
rect 42797 13277 42809 13311
rect 42843 13308 42855 13311
rect 42886 13308 42892 13320
rect 42843 13280 42892 13308
rect 42843 13277 42855 13280
rect 42797 13271 42855 13277
rect 42886 13268 42892 13280
rect 42944 13268 42950 13320
rect 48498 13308 48504 13320
rect 48459 13280 48504 13308
rect 48498 13268 48504 13280
rect 48556 13268 48562 13320
rect 50801 13311 50859 13317
rect 50801 13277 50813 13311
rect 50847 13308 50859 13311
rect 51258 13308 51264 13320
rect 50847 13280 51264 13308
rect 50847 13277 50859 13280
rect 50801 13271 50859 13277
rect 51258 13268 51264 13280
rect 51316 13268 51322 13320
rect 51368 13308 51396 13407
rect 53576 13376 53604 13484
rect 54570 13472 54576 13484
rect 54628 13472 54634 13524
rect 55030 13472 55036 13524
rect 55088 13512 55094 13524
rect 55677 13515 55735 13521
rect 55677 13512 55689 13515
rect 55088 13484 55689 13512
rect 55088 13472 55094 13484
rect 55677 13481 55689 13484
rect 55723 13481 55735 13515
rect 57701 13515 57759 13521
rect 57701 13512 57713 13515
rect 55677 13475 55735 13481
rect 56336 13484 57713 13512
rect 54757 13447 54815 13453
rect 54757 13413 54769 13447
rect 54803 13413 54815 13447
rect 54757 13407 54815 13413
rect 54772 13376 54800 13407
rect 54846 13404 54852 13456
rect 54904 13444 54910 13456
rect 56336 13444 56364 13484
rect 57701 13481 57713 13484
rect 57747 13481 57759 13515
rect 57701 13475 57759 13481
rect 54904 13416 56364 13444
rect 54904 13404 54910 13416
rect 55214 13376 55220 13388
rect 53576 13348 54064 13376
rect 54772 13348 55220 13376
rect 51997 13311 52055 13317
rect 51997 13308 52009 13311
rect 51368 13280 52009 13308
rect 51997 13277 52009 13280
rect 52043 13277 52055 13311
rect 53282 13308 53288 13320
rect 53243 13280 53288 13308
rect 51997 13271 52055 13277
rect 53282 13268 53288 13280
rect 53340 13268 53346 13320
rect 53469 13311 53527 13317
rect 53469 13277 53481 13311
rect 53515 13308 53527 13311
rect 53926 13308 53932 13320
rect 53515 13280 53932 13308
rect 53515 13277 53527 13280
rect 53469 13271 53527 13277
rect 53926 13268 53932 13280
rect 53984 13268 53990 13320
rect 54036 13308 54064 13348
rect 55214 13336 55220 13348
rect 55272 13376 55278 13388
rect 55309 13379 55367 13385
rect 55309 13376 55321 13379
rect 55272 13348 55321 13376
rect 55272 13336 55278 13348
rect 55309 13345 55321 13348
rect 55355 13345 55367 13379
rect 55309 13339 55367 13345
rect 56318 13308 56324 13320
rect 54036 13280 55260 13308
rect 56279 13280 56324 13308
rect 31726 13212 33825 13240
rect 33873 13243 33931 13249
rect 33873 13209 33885 13243
rect 33919 13240 33931 13243
rect 34606 13240 34612 13252
rect 33919 13212 34612 13240
rect 33919 13209 33931 13212
rect 33873 13203 33931 13209
rect 34606 13200 34612 13212
rect 34664 13200 34670 13252
rect 38672 13240 38700 13268
rect 41046 13240 41052 13252
rect 34716 13212 38700 13240
rect 41007 13212 41052 13240
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 2130 13172 2136 13184
rect 2091 13144 2136 13172
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 5169 13175 5227 13181
rect 5169 13172 5181 13175
rect 4672 13144 5181 13172
rect 4672 13132 4678 13144
rect 5169 13141 5181 13144
rect 5215 13141 5227 13175
rect 5169 13135 5227 13141
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 7558 13172 7564 13184
rect 7248 13144 7564 13172
rect 7248 13132 7254 13144
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 7926 13132 7932 13184
rect 7984 13172 7990 13184
rect 8478 13172 8484 13184
rect 7984 13144 8484 13172
rect 7984 13132 7990 13144
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 10505 13175 10563 13181
rect 10505 13141 10517 13175
rect 10551 13172 10563 13175
rect 11514 13172 11520 13184
rect 10551 13144 11520 13172
rect 10551 13141 10563 13144
rect 10505 13135 10563 13141
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 15473 13175 15531 13181
rect 15473 13172 15485 13175
rect 14608 13144 15485 13172
rect 14608 13132 14614 13144
rect 15473 13141 15485 13144
rect 15519 13141 15531 13175
rect 15473 13135 15531 13141
rect 20349 13175 20407 13181
rect 20349 13141 20361 13175
rect 20395 13172 20407 13175
rect 20622 13172 20628 13184
rect 20395 13144 20628 13172
rect 20395 13141 20407 13144
rect 20349 13135 20407 13141
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 21726 13132 21732 13184
rect 21784 13172 21790 13184
rect 22186 13172 22192 13184
rect 21784 13144 22192 13172
rect 21784 13132 21790 13144
rect 22186 13132 22192 13144
rect 22244 13172 22250 13184
rect 22649 13175 22707 13181
rect 22649 13172 22661 13175
rect 22244 13144 22661 13172
rect 22244 13132 22250 13144
rect 22649 13141 22661 13144
rect 22695 13172 22707 13175
rect 24026 13172 24032 13184
rect 22695 13144 24032 13172
rect 22695 13141 22707 13144
rect 22649 13135 22707 13141
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 26602 13172 26608 13184
rect 26563 13144 26608 13172
rect 26602 13132 26608 13144
rect 26660 13132 26666 13184
rect 31662 13172 31668 13184
rect 31623 13144 31668 13172
rect 31662 13132 31668 13144
rect 31720 13132 31726 13184
rect 33318 13132 33324 13184
rect 33376 13172 33382 13184
rect 34716 13172 34744 13212
rect 41046 13200 41052 13212
rect 41104 13200 41110 13252
rect 46106 13200 46112 13252
rect 46164 13240 46170 13252
rect 46262 13243 46320 13249
rect 46262 13240 46274 13243
rect 46164 13212 46274 13240
rect 46164 13200 46170 13212
rect 46262 13209 46274 13212
rect 46308 13209 46320 13243
rect 46262 13203 46320 13209
rect 48682 13200 48688 13252
rect 48740 13240 48746 13252
rect 53377 13243 53435 13249
rect 53377 13240 53389 13243
rect 48740 13212 53389 13240
rect 48740 13200 48746 13212
rect 53377 13209 53389 13212
rect 53423 13209 53435 13243
rect 53377 13203 53435 13209
rect 54110 13200 54116 13252
rect 54168 13240 54174 13252
rect 54389 13243 54447 13249
rect 54389 13240 54401 13243
rect 54168 13212 54401 13240
rect 54168 13200 54174 13212
rect 54389 13209 54401 13212
rect 54435 13240 54447 13243
rect 54846 13240 54852 13252
rect 54435 13212 54852 13240
rect 54435 13209 54447 13212
rect 54389 13203 54447 13209
rect 54846 13200 54852 13212
rect 54904 13200 54910 13252
rect 55232 13240 55260 13280
rect 56318 13268 56324 13280
rect 56376 13268 56382 13320
rect 55677 13243 55735 13249
rect 55677 13240 55689 13243
rect 55232 13212 55689 13240
rect 55677 13209 55689 13212
rect 55723 13209 55735 13243
rect 55677 13203 55735 13209
rect 56042 13200 56048 13252
rect 56100 13240 56106 13252
rect 56566 13243 56624 13249
rect 56566 13240 56578 13243
rect 56100 13212 56578 13240
rect 56100 13200 56106 13212
rect 56566 13209 56578 13212
rect 56612 13209 56624 13243
rect 56566 13203 56624 13209
rect 38562 13172 38568 13184
rect 33376 13144 34744 13172
rect 38523 13144 38568 13172
rect 33376 13132 33382 13144
rect 38562 13132 38568 13144
rect 38620 13132 38626 13184
rect 38933 13175 38991 13181
rect 38933 13141 38945 13175
rect 38979 13172 38991 13175
rect 39114 13172 39120 13184
rect 38979 13144 39120 13172
rect 38979 13141 38991 13144
rect 38933 13135 38991 13141
rect 39114 13132 39120 13144
rect 39172 13132 39178 13184
rect 42242 13132 42248 13184
rect 42300 13172 42306 13184
rect 42613 13175 42671 13181
rect 42613 13172 42625 13175
rect 42300 13144 42625 13172
rect 42300 13132 42306 13144
rect 42613 13141 42625 13144
rect 42659 13141 42671 13175
rect 47394 13172 47400 13184
rect 47355 13144 47400 13172
rect 42613 13135 42671 13141
rect 47394 13132 47400 13144
rect 47452 13132 47458 13184
rect 48590 13172 48596 13184
rect 48551 13144 48596 13172
rect 48590 13132 48596 13144
rect 48648 13132 48654 13184
rect 51166 13172 51172 13184
rect 51127 13144 51172 13172
rect 51166 13132 51172 13144
rect 51224 13132 51230 13184
rect 51810 13172 51816 13184
rect 51771 13144 51816 13172
rect 51810 13132 51816 13144
rect 51868 13132 51874 13184
rect 51994 13132 52000 13184
rect 52052 13172 52058 13184
rect 54589 13175 54647 13181
rect 54589 13172 54601 13175
rect 52052 13144 54601 13172
rect 52052 13132 52058 13144
rect 54589 13141 54601 13144
rect 54635 13141 54647 13175
rect 54589 13135 54647 13141
rect 55861 13175 55919 13181
rect 55861 13141 55873 13175
rect 55907 13172 55919 13175
rect 56226 13172 56232 13184
rect 55907 13144 56232 13172
rect 55907 13141 55919 13144
rect 55861 13135 55919 13141
rect 56226 13132 56232 13144
rect 56284 13132 56290 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 4062 12968 4068 12980
rect 4023 12940 4068 12968
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 4433 12971 4491 12977
rect 4433 12937 4445 12971
rect 4479 12968 4491 12971
rect 4614 12968 4620 12980
rect 4479 12940 4620 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 7374 12968 7380 12980
rect 7156 12940 7380 12968
rect 7156 12928 7162 12940
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 10410 12968 10416 12980
rect 7800 12940 10416 12968
rect 7800 12928 7806 12940
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 14182 12968 14188 12980
rect 10520 12940 12434 12968
rect 14143 12940 14188 12968
rect 2225 12903 2283 12909
rect 2225 12869 2237 12903
rect 2271 12900 2283 12903
rect 10520 12900 10548 12940
rect 10778 12900 10784 12912
rect 2271 12872 10548 12900
rect 10704 12872 10784 12900
rect 2271 12869 2283 12872
rect 2225 12863 2283 12869
rect 1854 12832 1860 12844
rect 1815 12804 1860 12832
rect 1854 12792 1860 12804
rect 1912 12792 1918 12844
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12801 2743 12835
rect 3602 12832 3608 12844
rect 3563 12804 3608 12832
rect 2685 12795 2743 12801
rect 2700 12764 2728 12795
rect 3602 12792 3608 12804
rect 3660 12792 3666 12844
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12801 4307 12835
rect 4249 12795 4307 12801
rect 2700 12736 4108 12764
rect 2866 12628 2872 12640
rect 2827 12600 2872 12628
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 3418 12628 3424 12640
rect 3379 12600 3424 12628
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 4080 12628 4108 12736
rect 4264 12696 4292 12795
rect 4338 12792 4344 12844
rect 4396 12832 4402 12844
rect 4525 12835 4583 12841
rect 4525 12832 4537 12835
rect 4396 12804 4537 12832
rect 4396 12792 4402 12804
rect 4525 12801 4537 12804
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 6638 12832 6644 12844
rect 5316 12804 6644 12832
rect 5316 12792 5322 12804
rect 6638 12792 6644 12804
rect 6696 12832 6702 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 6696 12804 7205 12832
rect 6696 12792 6702 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 7432 12804 7481 12832
rect 7432 12792 7438 12804
rect 7469 12801 7481 12804
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 7616 12804 8217 12832
rect 7616 12792 7622 12804
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 8389 12835 8447 12841
rect 8389 12801 8401 12835
rect 8435 12832 8447 12835
rect 8478 12832 8484 12844
rect 8435 12804 8484 12832
rect 8435 12801 8447 12804
rect 8389 12795 8447 12801
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12832 10655 12835
rect 10704 12832 10732 12872
rect 10778 12860 10784 12872
rect 10836 12860 10842 12912
rect 12406 12900 12434 12940
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 14550 12968 14556 12980
rect 14511 12940 14556 12968
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 24026 12968 24032 12980
rect 17236 12940 24032 12968
rect 17236 12900 17264 12940
rect 24026 12928 24032 12940
rect 24084 12928 24090 12980
rect 24121 12971 24179 12977
rect 24121 12937 24133 12971
rect 24167 12968 24179 12971
rect 24486 12968 24492 12980
rect 24167 12940 24492 12968
rect 24167 12937 24179 12940
rect 24121 12931 24179 12937
rect 24486 12928 24492 12940
rect 24544 12968 24550 12980
rect 24670 12968 24676 12980
rect 24544 12940 24676 12968
rect 24544 12928 24550 12940
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 24762 12928 24768 12980
rect 24820 12968 24826 12980
rect 25409 12971 25467 12977
rect 25409 12968 25421 12971
rect 24820 12940 25421 12968
rect 24820 12928 24826 12940
rect 25409 12937 25421 12940
rect 25455 12937 25467 12971
rect 31478 12968 31484 12980
rect 25409 12931 25467 12937
rect 30668 12940 31484 12968
rect 18138 12900 18144 12912
rect 12406 12872 17264 12900
rect 17328 12872 18144 12900
rect 11238 12832 11244 12844
rect 10643 12804 10732 12832
rect 10796 12804 11244 12832
rect 10643 12801 10655 12804
rect 10597 12795 10655 12801
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12764 7343 12767
rect 7742 12764 7748 12776
rect 7331 12736 7748 12764
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 8110 12724 8116 12776
rect 8168 12764 8174 12776
rect 10428 12764 10456 12795
rect 10796 12764 10824 12804
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11514 12832 11520 12844
rect 11475 12804 11520 12832
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 11790 12832 11796 12844
rect 11751 12804 11796 12832
rect 11790 12792 11796 12804
rect 11848 12832 11854 12844
rect 13814 12832 13820 12844
rect 11848 12804 13820 12832
rect 11848 12792 11854 12804
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14369 12835 14427 12841
rect 14369 12801 14381 12835
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12832 14703 12835
rect 15102 12832 15108 12844
rect 14691 12804 15108 12832
rect 14691 12801 14703 12804
rect 14645 12795 14703 12801
rect 8168 12736 10824 12764
rect 8168 12724 8174 12736
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 10928 12736 11621 12764
rect 10928 12724 10934 12736
rect 11609 12733 11621 12736
rect 11655 12733 11667 12767
rect 14384 12764 14412 12795
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 17129 12835 17187 12841
rect 17129 12801 17141 12835
rect 17175 12832 17187 12835
rect 17328 12832 17356 12872
rect 18138 12860 18144 12872
rect 18196 12860 18202 12912
rect 18506 12860 18512 12912
rect 18564 12900 18570 12912
rect 19337 12903 19395 12909
rect 19337 12900 19349 12903
rect 18564 12872 19349 12900
rect 18564 12860 18570 12872
rect 19337 12869 19349 12872
rect 19383 12869 19395 12903
rect 30558 12900 30564 12912
rect 19337 12863 19395 12869
rect 19536 12872 30564 12900
rect 17175 12804 17356 12832
rect 17396 12835 17454 12841
rect 17175 12801 17187 12804
rect 17129 12795 17187 12801
rect 17396 12801 17408 12835
rect 17442 12832 17454 12835
rect 18969 12835 19027 12841
rect 18969 12832 18981 12835
rect 17442 12804 18981 12832
rect 17442 12801 17454 12804
rect 17396 12795 17454 12801
rect 18969 12801 18981 12804
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 19153 12835 19211 12841
rect 19153 12801 19165 12835
rect 19199 12801 19211 12835
rect 19426 12832 19432 12844
rect 19387 12804 19432 12832
rect 19153 12795 19211 12801
rect 19168 12764 19196 12795
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 19334 12764 19340 12776
rect 14384 12736 16160 12764
rect 19168 12736 19340 12764
rect 11609 12727 11667 12733
rect 7006 12696 7012 12708
rect 4264 12668 7012 12696
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 7653 12699 7711 12705
rect 7653 12665 7665 12699
rect 7699 12696 7711 12699
rect 9582 12696 9588 12708
rect 7699 12668 9588 12696
rect 7699 12665 7711 12668
rect 7653 12659 7711 12665
rect 9582 12656 9588 12668
rect 9640 12656 9646 12708
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 16022 12696 16028 12708
rect 9824 12668 16028 12696
rect 9824 12656 9830 12668
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 5442 12628 5448 12640
rect 4080 12600 5448 12628
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 7469 12631 7527 12637
rect 7469 12597 7481 12631
rect 7515 12628 7527 12631
rect 7834 12628 7840 12640
rect 7515 12600 7840 12628
rect 7515 12597 7527 12600
rect 7469 12591 7527 12597
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 8570 12628 8576 12640
rect 8531 12600 8576 12628
rect 8570 12588 8576 12600
rect 8628 12588 8634 12640
rect 10594 12628 10600 12640
rect 10555 12600 10600 12628
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 10781 12631 10839 12637
rect 10781 12597 10793 12631
rect 10827 12628 10839 12631
rect 11054 12628 11060 12640
rect 10827 12600 11060 12628
rect 10827 12597 10839 12600
rect 10781 12591 10839 12597
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 11296 12600 11529 12628
rect 11296 12588 11302 12600
rect 11517 12597 11529 12600
rect 11563 12597 11575 12631
rect 11517 12591 11575 12597
rect 11977 12631 12035 12637
rect 11977 12597 11989 12631
rect 12023 12628 12035 12631
rect 12802 12628 12808 12640
rect 12023 12600 12808 12628
rect 12023 12597 12035 12600
rect 11977 12591 12035 12597
rect 12802 12588 12808 12600
rect 12860 12588 12866 12640
rect 16132 12628 16160 12736
rect 19334 12724 19340 12736
rect 19392 12724 19398 12776
rect 18506 12696 18512 12708
rect 18467 12668 18512 12696
rect 18506 12656 18512 12668
rect 18564 12656 18570 12708
rect 19536 12628 19564 12872
rect 30558 12860 30564 12872
rect 30616 12860 30622 12912
rect 30668 12909 30696 12940
rect 31478 12928 31484 12940
rect 31536 12928 31542 12980
rect 46017 12971 46075 12977
rect 31588 12940 44772 12968
rect 30653 12903 30711 12909
rect 30653 12869 30665 12903
rect 30699 12869 30711 12903
rect 30853 12903 30911 12909
rect 30853 12900 30865 12903
rect 30653 12863 30711 12869
rect 30760 12872 30865 12900
rect 21910 12832 21916 12844
rect 21823 12804 21916 12832
rect 21910 12792 21916 12804
rect 21968 12832 21974 12844
rect 24029 12835 24087 12841
rect 24029 12832 24041 12835
rect 21968 12804 24041 12832
rect 21968 12792 21974 12804
rect 24029 12801 24041 12804
rect 24075 12801 24087 12835
rect 24029 12795 24087 12801
rect 24765 12835 24823 12841
rect 24765 12801 24777 12835
rect 24811 12832 24823 12835
rect 25593 12835 25651 12841
rect 25593 12832 25605 12835
rect 24811 12804 25605 12832
rect 24811 12801 24823 12804
rect 24765 12795 24823 12801
rect 25593 12801 25605 12804
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 22186 12724 22192 12776
rect 22244 12764 22250 12776
rect 22646 12764 22652 12776
rect 22244 12736 22652 12764
rect 22244 12724 22250 12736
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 22830 12724 22836 12776
rect 22888 12764 22894 12776
rect 22925 12767 22983 12773
rect 22925 12764 22937 12767
rect 22888 12736 22937 12764
rect 22888 12724 22894 12736
rect 22925 12733 22937 12736
rect 22971 12764 22983 12767
rect 24780 12764 24808 12795
rect 22971 12736 24808 12764
rect 22971 12733 22983 12736
rect 22925 12727 22983 12733
rect 25406 12724 25412 12776
rect 25464 12764 25470 12776
rect 30760 12764 30788 12872
rect 30853 12869 30865 12872
rect 30899 12900 30911 12903
rect 31588 12900 31616 12940
rect 30899 12872 31616 12900
rect 30899 12869 30911 12872
rect 30853 12863 30911 12869
rect 31662 12860 31668 12912
rect 31720 12900 31726 12912
rect 32370 12903 32428 12909
rect 32370 12900 32382 12903
rect 31720 12872 32382 12900
rect 31720 12860 31726 12872
rect 32370 12869 32382 12872
rect 32416 12869 32428 12903
rect 32370 12863 32428 12869
rect 35434 12860 35440 12912
rect 35492 12900 35498 12912
rect 35805 12903 35863 12909
rect 35805 12900 35817 12903
rect 35492 12872 35817 12900
rect 35492 12860 35498 12872
rect 35805 12869 35817 12872
rect 35851 12869 35863 12903
rect 35805 12863 35863 12869
rect 38372 12903 38430 12909
rect 38372 12869 38384 12903
rect 38418 12900 38430 12903
rect 38562 12900 38568 12912
rect 38418 12872 38568 12900
rect 38418 12869 38430 12872
rect 38372 12863 38430 12869
rect 38562 12860 38568 12872
rect 38620 12860 38626 12912
rect 39022 12860 39028 12912
rect 39080 12900 39086 12912
rect 40681 12903 40739 12909
rect 40681 12900 40693 12903
rect 39080 12872 40693 12900
rect 39080 12860 39086 12872
rect 32122 12832 32128 12844
rect 32083 12804 32128 12832
rect 32122 12792 32128 12804
rect 32180 12832 32186 12844
rect 32674 12832 32680 12844
rect 32180 12804 32680 12832
rect 32180 12792 32186 12804
rect 32674 12792 32680 12804
rect 32732 12792 32738 12844
rect 35621 12835 35679 12841
rect 35621 12801 35633 12835
rect 35667 12832 35679 12835
rect 35986 12832 35992 12844
rect 35667 12804 35992 12832
rect 35667 12801 35679 12804
rect 35621 12795 35679 12801
rect 35986 12792 35992 12804
rect 36044 12792 36050 12844
rect 37550 12792 37556 12844
rect 37608 12832 37614 12844
rect 38105 12835 38163 12841
rect 38105 12832 38117 12835
rect 37608 12804 38117 12832
rect 37608 12792 37614 12804
rect 38105 12801 38117 12804
rect 38151 12801 38163 12835
rect 38105 12795 38163 12801
rect 25464 12736 30788 12764
rect 35437 12767 35495 12773
rect 25464 12724 25470 12736
rect 35437 12733 35449 12767
rect 35483 12764 35495 12767
rect 35894 12764 35900 12776
rect 35483 12736 35900 12764
rect 35483 12733 35495 12736
rect 35437 12727 35495 12733
rect 35894 12724 35900 12736
rect 35952 12724 35958 12776
rect 21450 12656 21456 12708
rect 21508 12696 21514 12708
rect 22097 12699 22155 12705
rect 22097 12696 22109 12699
rect 21508 12668 22109 12696
rect 21508 12656 21514 12668
rect 22097 12665 22109 12668
rect 22143 12696 22155 12699
rect 30374 12696 30380 12708
rect 22143 12668 30380 12696
rect 22143 12665 22155 12668
rect 22097 12659 22155 12665
rect 30374 12656 30380 12668
rect 30432 12656 30438 12708
rect 30558 12656 30564 12708
rect 30616 12696 30622 12708
rect 31021 12699 31079 12705
rect 31021 12696 31033 12699
rect 30616 12668 31033 12696
rect 30616 12656 30622 12668
rect 31021 12665 31033 12668
rect 31067 12665 31079 12699
rect 40512 12696 40540 12872
rect 40681 12869 40693 12872
rect 40727 12869 40739 12903
rect 40681 12863 40739 12869
rect 41046 12860 41052 12912
rect 41104 12900 41110 12912
rect 41785 12903 41843 12909
rect 41785 12900 41797 12903
rect 41104 12872 41797 12900
rect 41104 12860 41110 12872
rect 41785 12869 41797 12872
rect 41831 12869 41843 12903
rect 41785 12863 41843 12869
rect 42426 12860 42432 12912
rect 42484 12900 42490 12912
rect 42797 12903 42855 12909
rect 42797 12900 42809 12903
rect 42484 12872 42809 12900
rect 42484 12860 42490 12872
rect 42797 12869 42809 12872
rect 42843 12869 42855 12903
rect 44744 12900 44772 12940
rect 46017 12937 46029 12971
rect 46063 12968 46075 12971
rect 46106 12968 46112 12980
rect 46063 12940 46112 12968
rect 46063 12937 46075 12940
rect 46017 12931 46075 12937
rect 46106 12928 46112 12940
rect 46164 12928 46170 12980
rect 48777 12971 48835 12977
rect 48777 12937 48789 12971
rect 48823 12968 48835 12971
rect 49050 12968 49056 12980
rect 48823 12940 49056 12968
rect 48823 12937 48835 12940
rect 48777 12931 48835 12937
rect 49050 12928 49056 12940
rect 49108 12928 49114 12980
rect 52178 12968 52184 12980
rect 52139 12940 52184 12968
rect 52178 12928 52184 12940
rect 52236 12928 52242 12980
rect 55030 12968 55036 12980
rect 54991 12940 55036 12968
rect 55030 12928 55036 12940
rect 55088 12928 55094 12980
rect 56042 12968 56048 12980
rect 56003 12940 56048 12968
rect 56042 12928 56048 12940
rect 56100 12928 56106 12980
rect 48038 12900 48044 12912
rect 44744 12872 48044 12900
rect 42797 12863 42855 12869
rect 48038 12860 48044 12872
rect 48096 12860 48102 12912
rect 51068 12903 51126 12909
rect 51068 12869 51080 12903
rect 51114 12900 51126 12903
rect 51810 12900 51816 12912
rect 51114 12872 51816 12900
rect 51114 12869 51126 12872
rect 51068 12863 51126 12869
rect 51810 12860 51816 12872
rect 51868 12860 51874 12912
rect 54570 12860 54576 12912
rect 54628 12900 54634 12912
rect 55122 12900 55128 12912
rect 54628 12872 55128 12900
rect 54628 12860 54634 12872
rect 55122 12860 55128 12872
rect 55180 12900 55186 12912
rect 55401 12903 55459 12909
rect 55401 12900 55413 12903
rect 55180 12872 55413 12900
rect 55180 12860 55186 12872
rect 55401 12869 55413 12872
rect 55447 12869 55459 12903
rect 55401 12863 55459 12869
rect 40589 12835 40647 12841
rect 40589 12801 40601 12835
rect 40635 12801 40647 12835
rect 40770 12832 40776 12844
rect 40731 12804 40776 12832
rect 40589 12795 40647 12801
rect 40604 12764 40632 12795
rect 40770 12792 40776 12804
rect 40828 12792 40834 12844
rect 41693 12835 41751 12841
rect 41693 12801 41705 12835
rect 41739 12801 41751 12835
rect 42610 12832 42616 12844
rect 42571 12804 42616 12832
rect 41693 12795 41751 12801
rect 41046 12764 41052 12776
rect 40604 12736 41052 12764
rect 41046 12724 41052 12736
rect 41104 12764 41110 12776
rect 41708 12764 41736 12795
rect 42610 12792 42616 12804
rect 42668 12792 42674 12844
rect 43441 12835 43499 12841
rect 43441 12801 43453 12835
rect 43487 12832 43499 12835
rect 44450 12832 44456 12844
rect 43487 12804 44456 12832
rect 43487 12801 43499 12804
rect 43441 12795 43499 12801
rect 44450 12792 44456 12804
rect 44508 12792 44514 12844
rect 46198 12832 46204 12844
rect 46159 12804 46204 12832
rect 46198 12792 46204 12804
rect 46256 12792 46262 12844
rect 48682 12832 48688 12844
rect 48643 12804 48688 12832
rect 48682 12792 48688 12804
rect 48740 12792 48746 12844
rect 48866 12832 48872 12844
rect 48827 12804 48872 12832
rect 48866 12792 48872 12804
rect 48924 12792 48930 12844
rect 50798 12832 50804 12844
rect 50759 12804 50804 12832
rect 50798 12792 50804 12804
rect 50856 12792 50862 12844
rect 54846 12792 54852 12844
rect 54904 12832 54910 12844
rect 55217 12835 55275 12841
rect 55217 12832 55229 12835
rect 54904 12804 55229 12832
rect 54904 12792 54910 12804
rect 55217 12801 55229 12804
rect 55263 12801 55275 12835
rect 55493 12835 55551 12841
rect 55493 12832 55505 12835
rect 55217 12795 55275 12801
rect 55416 12804 55505 12832
rect 55416 12776 55444 12804
rect 55493 12801 55505 12804
rect 55539 12801 55551 12835
rect 56226 12832 56232 12844
rect 56187 12804 56232 12832
rect 55493 12795 55551 12801
rect 56226 12792 56232 12804
rect 56284 12792 56290 12844
rect 42886 12764 42892 12776
rect 41104 12736 42892 12764
rect 41104 12724 41110 12736
rect 42886 12724 42892 12736
rect 42944 12724 42950 12776
rect 43530 12764 43536 12776
rect 43491 12736 43536 12764
rect 43530 12724 43536 12736
rect 43588 12724 43594 12776
rect 43714 12764 43720 12776
rect 43675 12736 43720 12764
rect 43714 12724 43720 12736
rect 43772 12724 43778 12776
rect 55398 12724 55404 12776
rect 55456 12724 55462 12776
rect 42981 12699 43039 12705
rect 40512 12668 41414 12696
rect 31021 12659 31079 12665
rect 16132 12600 19564 12628
rect 22922 12588 22928 12640
rect 22980 12628 22986 12640
rect 23106 12628 23112 12640
rect 22980 12600 23112 12628
rect 22980 12588 22986 12600
rect 23106 12588 23112 12600
rect 23164 12588 23170 12640
rect 24854 12628 24860 12640
rect 24767 12600 24860 12628
rect 24854 12588 24860 12600
rect 24912 12628 24918 12640
rect 25682 12628 25688 12640
rect 24912 12600 25688 12628
rect 24912 12588 24918 12600
rect 25682 12588 25688 12600
rect 25740 12588 25746 12640
rect 30834 12628 30840 12640
rect 30795 12600 30840 12628
rect 30834 12588 30840 12600
rect 30892 12588 30898 12640
rect 33502 12628 33508 12640
rect 33415 12600 33508 12628
rect 33502 12588 33508 12600
rect 33560 12628 33566 12640
rect 38838 12628 38844 12640
rect 33560 12600 38844 12628
rect 33560 12588 33566 12600
rect 38838 12588 38844 12600
rect 38896 12588 38902 12640
rect 39114 12588 39120 12640
rect 39172 12628 39178 12640
rect 39485 12631 39543 12637
rect 39485 12628 39497 12631
rect 39172 12600 39497 12628
rect 39172 12588 39178 12600
rect 39485 12597 39497 12600
rect 39531 12597 39543 12631
rect 41386 12628 41414 12668
rect 42981 12665 42993 12699
rect 43027 12696 43039 12699
rect 43990 12696 43996 12708
rect 43027 12668 43996 12696
rect 43027 12665 43039 12668
rect 42981 12659 43039 12665
rect 43990 12656 43996 12668
rect 44048 12656 44054 12708
rect 43530 12628 43536 12640
rect 41386 12600 43536 12628
rect 39485 12591 39543 12597
rect 43530 12588 43536 12600
rect 43588 12588 43594 12640
rect 43622 12588 43628 12640
rect 43680 12628 43686 12640
rect 43680 12600 43725 12628
rect 43680 12588 43686 12600
rect 51074 12588 51080 12640
rect 51132 12628 51138 12640
rect 54662 12628 54668 12640
rect 51132 12600 54668 12628
rect 51132 12588 51138 12600
rect 54662 12588 54668 12600
rect 54720 12628 54726 12640
rect 56318 12628 56324 12640
rect 54720 12600 56324 12628
rect 54720 12588 54726 12600
rect 56318 12588 56324 12600
rect 56376 12588 56382 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 6638 12424 6644 12436
rect 6599 12396 6644 12424
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 6825 12427 6883 12433
rect 6825 12393 6837 12427
rect 6871 12424 6883 12427
rect 7377 12427 7435 12433
rect 7377 12424 7389 12427
rect 6871 12396 7389 12424
rect 6871 12393 6883 12396
rect 6825 12387 6883 12393
rect 7377 12393 7389 12396
rect 7423 12393 7435 12427
rect 7377 12387 7435 12393
rect 14967 12427 15025 12433
rect 14967 12393 14979 12427
rect 15013 12424 15025 12427
rect 15838 12424 15844 12436
rect 15013 12396 15844 12424
rect 15013 12393 15025 12396
rect 14967 12387 15025 12393
rect 15838 12384 15844 12396
rect 15896 12424 15902 12436
rect 16209 12427 16267 12433
rect 16209 12424 16221 12427
rect 15896 12396 16221 12424
rect 15896 12384 15902 12396
rect 16209 12393 16221 12396
rect 16255 12393 16267 12427
rect 16390 12424 16396 12436
rect 16351 12396 16396 12424
rect 16209 12387 16267 12393
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 20806 12424 20812 12436
rect 20719 12396 20812 12424
rect 20806 12384 20812 12396
rect 20864 12424 20870 12436
rect 21269 12427 21327 12433
rect 21269 12424 21281 12427
rect 20864 12396 21281 12424
rect 20864 12384 20870 12396
rect 21269 12393 21281 12396
rect 21315 12424 21327 12427
rect 21358 12424 21364 12436
rect 21315 12396 21364 12424
rect 21315 12393 21327 12396
rect 21269 12387 21327 12393
rect 21358 12384 21364 12396
rect 21416 12424 21422 12436
rect 21729 12427 21787 12433
rect 21729 12424 21741 12427
rect 21416 12396 21741 12424
rect 21416 12384 21422 12396
rect 21729 12393 21741 12396
rect 21775 12393 21787 12427
rect 21910 12424 21916 12436
rect 21871 12396 21916 12424
rect 21729 12387 21787 12393
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 22278 12424 22284 12436
rect 22046 12396 22284 12424
rect 3234 12356 3240 12368
rect 3147 12328 3240 12356
rect 3234 12316 3240 12328
rect 3292 12356 3298 12368
rect 7190 12356 7196 12368
rect 3292 12328 7196 12356
rect 3292 12316 3298 12328
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 10778 12356 10784 12368
rect 9232 12328 10784 12356
rect 5994 12248 6000 12300
rect 6052 12288 6058 12300
rect 6549 12291 6607 12297
rect 6549 12288 6561 12291
rect 6052 12260 6561 12288
rect 6052 12248 6058 12260
rect 6549 12257 6561 12260
rect 6595 12257 6607 12291
rect 8294 12288 8300 12300
rect 6549 12251 6607 12257
rect 7116 12260 8300 12288
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12189 1915 12223
rect 1857 12183 1915 12189
rect 2124 12223 2182 12229
rect 2124 12189 2136 12223
rect 2170 12220 2182 12223
rect 3418 12220 3424 12232
rect 2170 12192 3424 12220
rect 2170 12189 2182 12192
rect 2124 12183 2182 12189
rect 1872 12152 1900 12183
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 6457 12223 6515 12229
rect 6457 12189 6469 12223
rect 6503 12220 6515 12223
rect 7116 12220 7144 12260
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 9232 12297 9260 12328
rect 10778 12316 10784 12328
rect 10836 12356 10842 12368
rect 15194 12356 15200 12368
rect 10836 12328 15200 12356
rect 10836 12316 10842 12328
rect 15194 12316 15200 12328
rect 15252 12316 15258 12368
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 21453 12359 21511 12365
rect 21453 12356 21465 12359
rect 19392 12328 21465 12356
rect 19392 12316 19398 12328
rect 21453 12325 21465 12328
rect 21499 12356 21511 12359
rect 22046 12356 22074 12396
rect 22278 12384 22284 12396
rect 22336 12384 22342 12436
rect 23106 12384 23112 12436
rect 23164 12424 23170 12436
rect 23164 12396 23209 12424
rect 23164 12384 23170 12396
rect 24026 12384 24032 12436
rect 24084 12424 24090 12436
rect 24581 12427 24639 12433
rect 24581 12424 24593 12427
rect 24084 12396 24593 12424
rect 24084 12384 24090 12396
rect 24581 12393 24593 12396
rect 24627 12424 24639 12427
rect 24670 12424 24676 12436
rect 24627 12396 24676 12424
rect 24627 12393 24639 12396
rect 24581 12387 24639 12393
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 25590 12424 25596 12436
rect 25551 12396 25596 12424
rect 25590 12384 25596 12396
rect 25648 12384 25654 12436
rect 27430 12424 27436 12436
rect 26068 12396 27436 12424
rect 21499 12328 22074 12356
rect 21499 12325 21511 12328
rect 21453 12319 21511 12325
rect 8941 12291 8999 12297
rect 8941 12288 8953 12291
rect 8628 12260 8953 12288
rect 8628 12248 8634 12260
rect 8941 12257 8953 12260
rect 8987 12257 8999 12291
rect 8941 12251 8999 12257
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12257 9275 12291
rect 9217 12251 9275 12257
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 11701 12291 11759 12297
rect 9640 12260 10732 12288
rect 9640 12248 9646 12260
rect 7282 12220 7288 12232
rect 6503 12192 7144 12220
rect 7243 12192 7288 12220
rect 6503 12189 6515 12192
rect 6457 12183 6515 12189
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 7524 12192 7665 12220
rect 7524 12180 7530 12192
rect 7653 12189 7665 12192
rect 7699 12189 7711 12223
rect 10226 12220 10232 12232
rect 10187 12192 10232 12220
rect 7653 12183 7711 12189
rect 2590 12152 2596 12164
rect 1872 12124 2596 12152
rect 2590 12112 2596 12124
rect 2648 12112 2654 12164
rect 7668 12152 7696 12183
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10704 12229 10732 12260
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 16022 12288 16028 12300
rect 11747 12260 16028 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 16390 12248 16396 12300
rect 16448 12288 16454 12300
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 16448 12260 17233 12288
rect 16448 12248 16454 12260
rect 17221 12257 17233 12260
rect 17267 12288 17279 12291
rect 17402 12288 17408 12300
rect 17267 12260 17408 12288
rect 17267 12257 17279 12260
rect 17221 12251 17279 12257
rect 17402 12248 17408 12260
rect 17460 12248 17466 12300
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12288 17555 12291
rect 18046 12288 18052 12300
rect 17543 12260 18052 12288
rect 17543 12257 17555 12260
rect 17497 12251 17555 12257
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 18966 12248 18972 12300
rect 19024 12288 19030 12300
rect 21542 12288 21548 12300
rect 19024 12260 21548 12288
rect 19024 12248 19030 12260
rect 21542 12248 21548 12260
rect 21600 12248 21606 12300
rect 23106 12248 23112 12300
rect 23164 12288 23170 12300
rect 26068 12297 26096 12396
rect 27430 12384 27436 12396
rect 27488 12424 27494 12436
rect 29454 12424 29460 12436
rect 27488 12396 29460 12424
rect 27488 12384 27494 12396
rect 29454 12384 29460 12396
rect 29512 12384 29518 12436
rect 29822 12384 29828 12436
rect 29880 12424 29886 12436
rect 30929 12427 30987 12433
rect 30929 12424 30941 12427
rect 29880 12396 30941 12424
rect 29880 12384 29886 12396
rect 30929 12393 30941 12396
rect 30975 12393 30987 12427
rect 31846 12424 31852 12436
rect 31807 12396 31852 12424
rect 30929 12387 30987 12393
rect 31846 12384 31852 12396
rect 31904 12384 31910 12436
rect 38746 12384 38752 12436
rect 38804 12424 38810 12436
rect 39853 12427 39911 12433
rect 39853 12424 39865 12427
rect 38804 12396 39865 12424
rect 38804 12384 38810 12396
rect 39853 12393 39865 12396
rect 39899 12393 39911 12427
rect 39853 12387 39911 12393
rect 39942 12384 39948 12436
rect 40000 12424 40006 12436
rect 40000 12396 42472 12424
rect 40000 12384 40006 12396
rect 34977 12359 35035 12365
rect 34977 12325 34989 12359
rect 35023 12356 35035 12359
rect 37274 12356 37280 12368
rect 35023 12328 37280 12356
rect 35023 12325 35035 12328
rect 34977 12319 35035 12325
rect 37274 12316 37280 12328
rect 37332 12316 37338 12368
rect 38657 12359 38715 12365
rect 38657 12325 38669 12359
rect 38703 12325 38715 12359
rect 38657 12319 38715 12325
rect 42245 12359 42303 12365
rect 42245 12325 42257 12359
rect 42291 12356 42303 12359
rect 42334 12356 42340 12368
rect 42291 12328 42340 12356
rect 42291 12325 42303 12328
rect 42245 12319 42303 12325
rect 26053 12291 26111 12297
rect 23164 12260 25268 12288
rect 23164 12248 23170 12260
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12189 10747 12223
rect 11054 12220 11060 12232
rect 11015 12192 11060 12220
rect 10689 12183 10747 12189
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11422 12220 11428 12232
rect 11383 12192 11428 12220
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12621 12223 12679 12229
rect 12621 12220 12633 12223
rect 12492 12192 12633 12220
rect 12492 12180 12498 12192
rect 12621 12189 12633 12192
rect 12667 12189 12679 12223
rect 12802 12220 12808 12232
rect 12763 12192 12808 12220
rect 12621 12183 12679 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 14734 12220 14740 12232
rect 14695 12192 14740 12220
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 15930 12180 15936 12232
rect 15988 12220 15994 12232
rect 16298 12220 16304 12232
rect 15988 12192 16304 12220
rect 15988 12180 15994 12192
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 21818 12220 21824 12232
rect 17880 12192 21824 12220
rect 10244 12152 10272 12180
rect 7668 12124 10272 12152
rect 12989 12155 13047 12161
rect 12989 12121 13001 12155
rect 13035 12152 13047 12155
rect 13722 12152 13728 12164
rect 13035 12124 13728 12152
rect 13035 12121 13047 12124
rect 12989 12115 13047 12121
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 15562 12112 15568 12164
rect 15620 12152 15626 12164
rect 16025 12155 16083 12161
rect 16025 12152 16037 12155
rect 15620 12124 16037 12152
rect 15620 12112 15626 12124
rect 16025 12121 16037 12124
rect 16071 12152 16083 12155
rect 17880 12152 17908 12192
rect 21818 12180 21824 12192
rect 21876 12180 21882 12232
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12220 22155 12223
rect 22370 12220 22376 12232
rect 22143 12192 22376 12220
rect 22143 12189 22155 12192
rect 22097 12183 22155 12189
rect 21082 12152 21088 12164
rect 16071 12124 17908 12152
rect 21043 12124 21088 12152
rect 16071 12121 16083 12124
rect 16025 12115 16083 12121
rect 21082 12112 21088 12124
rect 21140 12112 21146 12164
rect 21301 12155 21359 12161
rect 21301 12121 21313 12155
rect 21347 12152 21359 12155
rect 21726 12152 21732 12164
rect 21347 12124 21732 12152
rect 21347 12121 21359 12124
rect 21301 12115 21359 12121
rect 21726 12112 21732 12124
rect 21784 12112 21790 12164
rect 21928 12152 21956 12183
rect 22370 12180 22376 12192
rect 22428 12180 22434 12232
rect 22830 12180 22836 12232
rect 22888 12220 22894 12232
rect 25240 12229 25268 12260
rect 26053 12257 26065 12291
rect 26099 12257 26111 12291
rect 26053 12251 26111 12257
rect 29454 12248 29460 12300
rect 29512 12288 29518 12300
rect 29549 12291 29607 12297
rect 29549 12288 29561 12291
rect 29512 12260 29561 12288
rect 29512 12248 29518 12260
rect 29549 12257 29561 12260
rect 29595 12257 29607 12291
rect 36630 12288 36636 12300
rect 29549 12251 29607 12257
rect 31312 12260 36636 12288
rect 22999 12223 23057 12229
rect 22999 12220 23011 12223
rect 22888 12192 23011 12220
rect 22888 12180 22894 12192
rect 22999 12189 23011 12192
rect 23045 12189 23057 12223
rect 22999 12183 23057 12189
rect 25225 12223 25283 12229
rect 25225 12189 25237 12223
rect 25271 12189 25283 12223
rect 25225 12183 25283 12189
rect 28534 12180 28540 12232
rect 28592 12220 28598 12232
rect 28813 12223 28871 12229
rect 28813 12220 28825 12223
rect 28592 12192 28825 12220
rect 28592 12180 28598 12192
rect 28813 12189 28825 12192
rect 28859 12189 28871 12223
rect 28813 12183 28871 12189
rect 28902 12180 28908 12232
rect 28960 12220 28966 12232
rect 31312 12220 31340 12260
rect 36630 12248 36636 12260
rect 36688 12288 36694 12300
rect 38010 12288 38016 12300
rect 36688 12260 38016 12288
rect 36688 12248 36694 12260
rect 38010 12248 38016 12260
rect 38068 12248 38074 12300
rect 38672 12288 38700 12319
rect 42334 12316 42340 12328
rect 42392 12316 42398 12368
rect 42444 12356 42472 12396
rect 42518 12384 42524 12436
rect 42576 12424 42582 12436
rect 43070 12424 43076 12436
rect 42576 12396 43076 12424
rect 42576 12384 42582 12396
rect 43070 12384 43076 12396
rect 43128 12384 43134 12436
rect 43180 12396 43668 12424
rect 43180 12356 43208 12396
rect 42444 12328 43208 12356
rect 43254 12316 43260 12368
rect 43312 12356 43318 12368
rect 43312 12328 43484 12356
rect 43312 12316 43318 12328
rect 42352 12288 42380 12316
rect 38672 12260 39160 12288
rect 42352 12260 43208 12288
rect 39132 12232 39160 12260
rect 31478 12220 31484 12232
rect 28960 12192 31340 12220
rect 31439 12192 31484 12220
rect 28960 12180 28966 12192
rect 31478 12180 31484 12192
rect 31536 12180 31542 12232
rect 31665 12223 31723 12229
rect 31665 12189 31677 12223
rect 31711 12189 31723 12223
rect 31665 12183 31723 12189
rect 22848 12152 22876 12180
rect 21928 12124 22876 12152
rect 23474 12112 23480 12164
rect 23532 12152 23538 12164
rect 24397 12155 24455 12161
rect 24397 12152 24409 12155
rect 23532 12124 24409 12152
rect 23532 12112 23538 12124
rect 24397 12121 24409 12124
rect 24443 12121 24455 12155
rect 24397 12115 24455 12121
rect 24613 12155 24671 12161
rect 24613 12121 24625 12155
rect 24659 12152 24671 12155
rect 24854 12152 24860 12164
rect 24659 12124 24860 12152
rect 24659 12121 24671 12124
rect 24613 12115 24671 12121
rect 24854 12112 24860 12124
rect 24912 12112 24918 12164
rect 25409 12155 25467 12161
rect 25409 12121 25421 12155
rect 25455 12152 25467 12155
rect 25590 12152 25596 12164
rect 25455 12124 25596 12152
rect 25455 12121 25467 12124
rect 25409 12115 25467 12121
rect 25590 12112 25596 12124
rect 25648 12112 25654 12164
rect 26320 12155 26378 12161
rect 26320 12121 26332 12155
rect 26366 12152 26378 12155
rect 26602 12152 26608 12164
rect 26366 12124 26608 12152
rect 26366 12121 26378 12124
rect 26320 12115 26378 12121
rect 26602 12112 26608 12124
rect 26660 12112 26666 12164
rect 29794 12155 29852 12161
rect 29794 12152 29806 12155
rect 28644 12124 29806 12152
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 7837 12087 7895 12093
rect 7837 12084 7849 12087
rect 7524 12056 7849 12084
rect 7524 12044 7530 12056
rect 7837 12053 7849 12056
rect 7883 12053 7895 12087
rect 7837 12047 7895 12053
rect 7926 12044 7932 12096
rect 7984 12084 7990 12096
rect 12618 12084 12624 12096
rect 7984 12056 12624 12084
rect 7984 12044 7990 12056
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 13630 12084 13636 12096
rect 13136 12056 13636 12084
rect 13136 12044 13142 12056
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 16235 12087 16293 12093
rect 16235 12053 16247 12087
rect 16281 12084 16293 12087
rect 16574 12084 16580 12096
rect 16281 12056 16580 12084
rect 16281 12053 16293 12056
rect 16235 12047 16293 12053
rect 16574 12044 16580 12056
rect 16632 12044 16638 12096
rect 22738 12044 22744 12096
rect 22796 12084 22802 12096
rect 24765 12087 24823 12093
rect 24765 12084 24777 12087
rect 22796 12056 24777 12084
rect 22796 12044 22802 12056
rect 24765 12053 24777 12056
rect 24811 12084 24823 12087
rect 25222 12084 25228 12096
rect 24811 12056 25228 12084
rect 24811 12053 24823 12056
rect 24765 12047 24823 12053
rect 25222 12044 25228 12056
rect 25280 12044 25286 12096
rect 25608 12084 25636 12112
rect 28644 12093 28672 12124
rect 29794 12121 29806 12124
rect 29840 12121 29852 12155
rect 31680 12152 31708 12183
rect 34514 12180 34520 12232
rect 34572 12220 34578 12232
rect 35253 12223 35311 12229
rect 35253 12220 35265 12223
rect 34572 12192 35265 12220
rect 34572 12180 34578 12192
rect 35253 12189 35265 12192
rect 35299 12189 35311 12223
rect 35253 12183 35311 12189
rect 35986 12180 35992 12232
rect 36044 12220 36050 12232
rect 36173 12223 36231 12229
rect 36173 12220 36185 12223
rect 36044 12192 36185 12220
rect 36044 12180 36050 12192
rect 36173 12189 36185 12192
rect 36219 12220 36231 12223
rect 36722 12220 36728 12232
rect 36219 12192 36728 12220
rect 36219 12189 36231 12192
rect 36173 12183 36231 12189
rect 36722 12180 36728 12192
rect 36780 12180 36786 12232
rect 38562 12229 38568 12232
rect 38555 12223 38568 12229
rect 38555 12220 38567 12223
rect 38523 12192 38567 12220
rect 38555 12189 38567 12192
rect 38555 12183 38568 12189
rect 38562 12180 38568 12183
rect 38620 12180 38626 12232
rect 38746 12220 38752 12232
rect 38707 12192 38752 12220
rect 38746 12180 38752 12192
rect 38804 12180 38810 12232
rect 38838 12180 38844 12232
rect 38896 12220 38902 12232
rect 38896 12192 38941 12220
rect 38896 12180 38902 12192
rect 39114 12180 39120 12232
rect 39172 12220 39178 12232
rect 39853 12223 39911 12229
rect 39853 12220 39865 12223
rect 39172 12192 39865 12220
rect 39172 12180 39178 12192
rect 39853 12189 39865 12192
rect 39899 12189 39911 12223
rect 39853 12183 39911 12189
rect 40037 12223 40095 12229
rect 40037 12189 40049 12223
rect 40083 12220 40095 12223
rect 40770 12220 40776 12232
rect 40083 12192 40776 12220
rect 40083 12189 40095 12192
rect 40037 12183 40095 12189
rect 40770 12180 40776 12192
rect 40828 12180 40834 12232
rect 42518 12180 42524 12232
rect 42576 12220 42582 12232
rect 43053 12223 43111 12229
rect 43180 12226 43208 12260
rect 43053 12220 43065 12223
rect 42576 12217 42912 12220
rect 42996 12217 43065 12220
rect 42576 12192 43065 12217
rect 42576 12180 42582 12192
rect 42884 12189 43024 12192
rect 43053 12189 43065 12192
rect 43099 12189 43111 12223
rect 42884 12186 42932 12189
rect 43053 12183 43111 12189
rect 43162 12220 43220 12226
rect 43162 12186 43174 12220
rect 43208 12186 43220 12220
rect 43162 12180 43220 12186
rect 43254 12180 43260 12232
rect 43312 12220 43318 12232
rect 43456 12229 43484 12328
rect 43640 12288 43668 12396
rect 43714 12384 43720 12436
rect 43772 12424 43778 12436
rect 44085 12427 44143 12433
rect 44085 12424 44097 12427
rect 43772 12396 44097 12424
rect 43772 12384 43778 12396
rect 44085 12393 44097 12396
rect 44131 12393 44143 12427
rect 44085 12387 44143 12393
rect 48317 12427 48375 12433
rect 48317 12393 48329 12427
rect 48363 12424 48375 12427
rect 48590 12424 48596 12436
rect 48363 12396 48596 12424
rect 48363 12393 48375 12396
rect 48317 12387 48375 12393
rect 48590 12384 48596 12396
rect 48648 12384 48654 12436
rect 50617 12427 50675 12433
rect 50617 12393 50629 12427
rect 50663 12424 50675 12427
rect 51166 12424 51172 12436
rect 50663 12396 51172 12424
rect 50663 12393 50675 12396
rect 50617 12387 50675 12393
rect 51166 12384 51172 12396
rect 51224 12384 51230 12436
rect 51442 12384 51448 12436
rect 51500 12424 51506 12436
rect 51813 12427 51871 12433
rect 51813 12424 51825 12427
rect 51500 12396 51825 12424
rect 51500 12384 51506 12396
rect 51813 12393 51825 12396
rect 51859 12424 51871 12427
rect 51902 12424 51908 12436
rect 51859 12396 51908 12424
rect 51859 12393 51871 12396
rect 51813 12387 51871 12393
rect 51902 12384 51908 12396
rect 51960 12384 51966 12436
rect 48225 12359 48283 12365
rect 48225 12325 48237 12359
rect 48271 12356 48283 12359
rect 48682 12356 48688 12368
rect 48271 12328 48688 12356
rect 48271 12325 48283 12328
rect 48225 12319 48283 12325
rect 48682 12316 48688 12328
rect 48740 12316 48746 12368
rect 51258 12316 51264 12368
rect 51316 12356 51322 12368
rect 51994 12356 52000 12368
rect 51316 12328 52000 12356
rect 51316 12316 51322 12328
rect 51994 12316 52000 12328
rect 52052 12316 52058 12368
rect 43640 12260 47348 12288
rect 43441 12223 43499 12229
rect 43312 12192 43357 12220
rect 43312 12180 43318 12192
rect 43441 12189 43453 12223
rect 43487 12189 43499 12223
rect 43990 12220 43996 12232
rect 43951 12192 43996 12220
rect 43441 12183 43499 12189
rect 43990 12180 43996 12192
rect 44048 12180 44054 12232
rect 47320 12220 47348 12260
rect 47394 12248 47400 12300
rect 47452 12288 47458 12300
rect 48409 12291 48467 12297
rect 48409 12288 48421 12291
rect 47452 12260 48421 12288
rect 47452 12248 47458 12260
rect 48409 12257 48421 12260
rect 48455 12257 48467 12291
rect 50801 12291 50859 12297
rect 50801 12288 50813 12291
rect 48409 12251 48467 12257
rect 48516 12260 50813 12288
rect 47670 12220 47676 12232
rect 47320 12192 47676 12220
rect 47670 12180 47676 12192
rect 47728 12220 47734 12232
rect 48133 12223 48191 12229
rect 48133 12220 48145 12223
rect 47728 12192 48145 12220
rect 47728 12180 47734 12192
rect 48133 12189 48145 12192
rect 48179 12220 48191 12223
rect 48314 12220 48320 12232
rect 48179 12192 48320 12220
rect 48179 12189 48191 12192
rect 48133 12183 48191 12189
rect 48314 12180 48320 12192
rect 48372 12220 48378 12232
rect 48516 12220 48544 12260
rect 50801 12257 50813 12260
rect 50847 12257 50859 12291
rect 50801 12251 50859 12257
rect 50893 12291 50951 12297
rect 50893 12257 50905 12291
rect 50939 12288 50951 12291
rect 51442 12288 51448 12300
rect 50939 12260 51448 12288
rect 50939 12257 50951 12260
rect 50893 12251 50951 12257
rect 51442 12248 51448 12260
rect 51500 12248 51506 12300
rect 55582 12288 55588 12300
rect 55543 12260 55588 12288
rect 55582 12248 55588 12260
rect 55640 12248 55646 12300
rect 48372 12192 48544 12220
rect 48593 12223 48651 12229
rect 48372 12180 48378 12192
rect 48593 12189 48605 12223
rect 48639 12220 48651 12223
rect 48682 12220 48688 12232
rect 48639 12192 48688 12220
rect 48639 12189 48651 12192
rect 48593 12183 48651 12189
rect 48682 12180 48688 12192
rect 48740 12180 48746 12232
rect 48774 12180 48780 12232
rect 48832 12220 48838 12232
rect 50985 12223 51043 12229
rect 50985 12220 50997 12223
rect 48832 12192 50997 12220
rect 48832 12180 48838 12192
rect 50985 12189 50997 12192
rect 51031 12189 51043 12223
rect 50985 12183 51043 12189
rect 51077 12223 51135 12229
rect 51077 12189 51089 12223
rect 51123 12189 51135 12223
rect 51077 12183 51135 12189
rect 29794 12115 29852 12121
rect 29932 12124 31708 12152
rect 34977 12155 35035 12161
rect 27433 12087 27491 12093
rect 27433 12084 27445 12087
rect 25608 12056 27445 12084
rect 27433 12053 27445 12056
rect 27479 12053 27491 12087
rect 27433 12047 27491 12053
rect 28629 12087 28687 12093
rect 28629 12053 28641 12087
rect 28675 12053 28687 12087
rect 28629 12047 28687 12053
rect 28810 12044 28816 12096
rect 28868 12084 28874 12096
rect 29932 12084 29960 12124
rect 34977 12121 34989 12155
rect 35023 12152 35035 12155
rect 36446 12152 36452 12164
rect 35023 12124 36452 12152
rect 35023 12121 35035 12124
rect 34977 12115 35035 12121
rect 36446 12112 36452 12124
rect 36504 12152 36510 12164
rect 36906 12152 36912 12164
rect 36504 12124 36912 12152
rect 36504 12112 36510 12124
rect 36906 12112 36912 12124
rect 36964 12112 36970 12164
rect 41690 12152 41696 12164
rect 38626 12124 41696 12152
rect 28868 12056 29960 12084
rect 28868 12044 28874 12056
rect 34790 12044 34796 12096
rect 34848 12084 34854 12096
rect 35161 12087 35219 12093
rect 35161 12084 35173 12087
rect 34848 12056 35173 12084
rect 34848 12044 34854 12056
rect 35161 12053 35173 12056
rect 35207 12084 35219 12087
rect 35618 12084 35624 12096
rect 35207 12056 35624 12084
rect 35207 12053 35219 12056
rect 35161 12047 35219 12053
rect 35618 12044 35624 12056
rect 35676 12084 35682 12096
rect 35897 12087 35955 12093
rect 35897 12084 35909 12087
rect 35676 12056 35909 12084
rect 35676 12044 35682 12056
rect 35897 12053 35909 12056
rect 35943 12084 35955 12087
rect 36538 12084 36544 12096
rect 35943 12056 36544 12084
rect 35943 12053 35955 12056
rect 35897 12047 35955 12053
rect 36538 12044 36544 12056
rect 36596 12044 36602 12096
rect 38378 12084 38384 12096
rect 38339 12056 38384 12084
rect 38378 12044 38384 12056
rect 38436 12044 38442 12096
rect 38470 12044 38476 12096
rect 38528 12084 38534 12096
rect 38626 12084 38654 12124
rect 41690 12112 41696 12124
rect 41748 12112 41754 12164
rect 41874 12152 41880 12164
rect 41835 12124 41880 12152
rect 41874 12112 41880 12124
rect 41932 12112 41938 12164
rect 51092 12152 51120 12183
rect 55122 12180 55128 12232
rect 55180 12220 55186 12232
rect 55309 12223 55367 12229
rect 55309 12220 55321 12223
rect 55180 12192 55321 12220
rect 55180 12180 55186 12192
rect 55309 12189 55321 12192
rect 55355 12189 55367 12223
rect 55309 12183 55367 12189
rect 55398 12180 55404 12232
rect 55456 12220 55462 12232
rect 55456 12192 55501 12220
rect 55456 12180 55462 12192
rect 51629 12155 51687 12161
rect 51629 12152 51641 12155
rect 51092 12124 51641 12152
rect 51629 12121 51641 12124
rect 51675 12152 51687 12155
rect 52178 12152 52184 12164
rect 51675 12124 52184 12152
rect 51675 12121 51687 12124
rect 51629 12115 51687 12121
rect 52178 12112 52184 12124
rect 52236 12112 52242 12164
rect 38528 12056 38654 12084
rect 42337 12087 42395 12093
rect 38528 12044 38534 12056
rect 42337 12053 42349 12087
rect 42383 12084 42395 12087
rect 42702 12084 42708 12096
rect 42383 12056 42708 12084
rect 42383 12053 42395 12056
rect 42337 12047 42395 12053
rect 42702 12044 42708 12056
rect 42760 12044 42766 12096
rect 42797 12087 42855 12093
rect 42797 12053 42809 12087
rect 42843 12084 42855 12087
rect 43990 12084 43996 12096
rect 42843 12056 43996 12084
rect 42843 12053 42855 12056
rect 42797 12047 42855 12053
rect 43990 12044 43996 12056
rect 44048 12044 44054 12096
rect 47854 12084 47860 12096
rect 47815 12056 47860 12084
rect 47854 12044 47860 12056
rect 47912 12044 47918 12096
rect 51534 12044 51540 12096
rect 51592 12084 51598 12096
rect 51829 12087 51887 12093
rect 51829 12084 51841 12087
rect 51592 12056 51841 12084
rect 51592 12044 51598 12056
rect 51829 12053 51841 12056
rect 51875 12053 51887 12087
rect 51829 12047 51887 12053
rect 53926 12044 53932 12096
rect 53984 12084 53990 12096
rect 55585 12087 55643 12093
rect 55585 12084 55597 12087
rect 53984 12056 55597 12084
rect 53984 12044 53990 12056
rect 55585 12053 55597 12056
rect 55631 12053 55643 12087
rect 55585 12047 55643 12053
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 2593 11883 2651 11889
rect 2593 11880 2605 11883
rect 2188 11852 2605 11880
rect 2188 11840 2194 11852
rect 2593 11849 2605 11852
rect 2639 11849 2651 11883
rect 2593 11843 2651 11849
rect 10965 11883 11023 11889
rect 10965 11849 10977 11883
rect 11011 11880 11023 11883
rect 11422 11880 11428 11892
rect 11011 11852 11428 11880
rect 11011 11849 11023 11852
rect 10965 11843 11023 11849
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 26878 11880 26884 11892
rect 11572 11852 26884 11880
rect 11572 11840 11578 11852
rect 26878 11840 26884 11852
rect 26936 11840 26942 11892
rect 26970 11840 26976 11892
rect 27028 11880 27034 11892
rect 33502 11880 33508 11892
rect 27028 11852 33508 11880
rect 27028 11840 27034 11852
rect 33502 11840 33508 11852
rect 33560 11840 33566 11892
rect 33594 11840 33600 11892
rect 33652 11880 33658 11892
rect 37090 11880 37096 11892
rect 33652 11852 37096 11880
rect 33652 11840 33658 11852
rect 37090 11840 37096 11852
rect 37148 11840 37154 11892
rect 41690 11840 41696 11892
rect 41748 11880 41754 11892
rect 46566 11880 46572 11892
rect 41748 11852 45600 11880
rect 46527 11852 46572 11880
rect 41748 11840 41754 11852
rect 5626 11812 5632 11824
rect 1412 11784 5488 11812
rect 5587 11784 5632 11812
rect 1412 11753 1440 11784
rect 1397 11747 1455 11753
rect 1397 11713 1409 11747
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11744 2559 11747
rect 3234 11744 3240 11756
rect 2547 11716 3240 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 3234 11704 3240 11716
rect 3292 11704 3298 11756
rect 3510 11744 3516 11756
rect 3471 11716 3516 11744
rect 3510 11704 3516 11716
rect 3568 11704 3574 11756
rect 5460 11744 5488 11784
rect 5626 11772 5632 11784
rect 5684 11772 5690 11824
rect 7466 11812 7472 11824
rect 7427 11784 7472 11812
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 10781 11815 10839 11821
rect 10781 11781 10793 11815
rect 10827 11812 10839 11815
rect 12434 11812 12440 11824
rect 10827 11784 12440 11812
rect 10827 11781 10839 11784
rect 10781 11775 10839 11781
rect 12434 11772 12440 11784
rect 12492 11772 12498 11824
rect 12618 11772 12624 11824
rect 12676 11812 12682 11824
rect 15562 11812 15568 11824
rect 12676 11784 14872 11812
rect 15523 11784 15568 11812
rect 12676 11772 12682 11784
rect 5902 11744 5908 11756
rect 5460 11716 5908 11744
rect 5902 11704 5908 11716
rect 5960 11704 5966 11756
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8665 11747 8723 11753
rect 8665 11744 8677 11747
rect 8536 11716 8677 11744
rect 8536 11704 8542 11716
rect 8665 11713 8677 11716
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 10100 11716 10609 11744
rect 10100 11704 10106 11716
rect 10597 11713 10609 11716
rect 10643 11744 10655 11747
rect 10870 11744 10876 11756
rect 10643 11716 10876 11744
rect 10643 11713 10655 11716
rect 10597 11707 10655 11713
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 2682 11676 2688 11688
rect 2643 11648 2688 11676
rect 2682 11636 2688 11648
rect 2740 11636 2746 11688
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 9398 11676 9404 11688
rect 8435 11648 9404 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 2133 11611 2191 11617
rect 2133 11577 2145 11611
rect 2179 11608 2191 11611
rect 3602 11608 3608 11620
rect 2179 11580 3608 11608
rect 2179 11577 2191 11580
rect 2133 11571 2191 11577
rect 3602 11568 3608 11580
rect 3660 11568 3666 11620
rect 8294 11568 8300 11620
rect 8352 11608 8358 11620
rect 12176 11608 12204 11707
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12308 11716 13001 11744
rect 12308 11704 12314 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 13170 11744 13176 11756
rect 13131 11716 13176 11744
rect 12989 11707 13047 11713
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 14844 11753 14872 11784
rect 15562 11772 15568 11784
rect 15620 11772 15626 11824
rect 16022 11772 16028 11824
rect 16080 11812 16086 11824
rect 22186 11812 22192 11824
rect 16080 11784 22192 11812
rect 16080 11772 16086 11784
rect 22186 11772 22192 11784
rect 22244 11772 22250 11824
rect 24118 11812 24124 11824
rect 24079 11784 24124 11812
rect 24118 11772 24124 11784
rect 24176 11772 24182 11824
rect 24486 11772 24492 11824
rect 24544 11812 24550 11824
rect 28445 11815 28503 11821
rect 28445 11812 28457 11815
rect 24544 11784 28457 11812
rect 24544 11772 24550 11784
rect 28445 11781 28457 11784
rect 28491 11781 28503 11815
rect 28445 11775 28503 11781
rect 28626 11772 28632 11824
rect 28684 11812 28690 11824
rect 41874 11812 41880 11824
rect 28684 11784 41880 11812
rect 28684 11772 28690 11784
rect 41874 11772 41880 11784
rect 41932 11772 41938 11824
rect 42886 11812 42892 11824
rect 42847 11784 42892 11812
rect 42886 11772 42892 11784
rect 42944 11772 42950 11824
rect 43070 11772 43076 11824
rect 43128 11812 43134 11824
rect 43128 11784 43760 11812
rect 43128 11772 43134 11784
rect 14829 11747 14887 11753
rect 14829 11713 14841 11747
rect 14875 11744 14887 11747
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 14875 11716 15485 11744
rect 14875 11713 14887 11716
rect 14829 11707 14887 11713
rect 15473 11713 15485 11716
rect 15519 11744 15531 11747
rect 15930 11744 15936 11756
rect 15519 11716 15936 11744
rect 15519 11713 15531 11716
rect 15473 11707 15531 11713
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 16758 11704 16764 11756
rect 16816 11744 16822 11756
rect 17126 11744 17132 11756
rect 16816 11716 17132 11744
rect 16816 11704 16822 11716
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 18966 11744 18972 11756
rect 18927 11716 18972 11744
rect 18966 11704 18972 11716
rect 19024 11704 19030 11756
rect 19150 11744 19156 11756
rect 19111 11716 19156 11744
rect 19150 11704 19156 11716
rect 19208 11704 19214 11756
rect 19245 11747 19303 11753
rect 19245 11713 19257 11747
rect 19291 11744 19303 11747
rect 19426 11744 19432 11756
rect 19291 11716 19432 11744
rect 19291 11713 19303 11716
rect 19245 11707 19303 11713
rect 19426 11704 19432 11716
rect 19484 11744 19490 11756
rect 19978 11744 19984 11756
rect 19484 11716 19984 11744
rect 19484 11704 19490 11716
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 22094 11704 22100 11756
rect 22152 11744 22158 11756
rect 22278 11744 22284 11756
rect 22152 11716 22197 11744
rect 22239 11716 22284 11744
rect 22152 11704 22158 11716
rect 22278 11704 22284 11716
rect 22336 11704 22342 11756
rect 23566 11704 23572 11756
rect 23624 11744 23630 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23624 11716 23949 11744
rect 23624 11704 23630 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 26418 11744 26424 11756
rect 23937 11707 23995 11713
rect 24136 11716 26424 11744
rect 13354 11676 13360 11688
rect 13096 11648 13360 11676
rect 13096 11620 13124 11648
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 15712 11648 15757 11676
rect 15712 11636 15718 11648
rect 16666 11636 16672 11688
rect 16724 11676 16730 11688
rect 16853 11679 16911 11685
rect 16853 11676 16865 11679
rect 16724 11648 16865 11676
rect 16724 11636 16730 11648
rect 16853 11645 16865 11648
rect 16899 11676 16911 11679
rect 16942 11676 16948 11688
rect 16899 11648 16948 11676
rect 16899 11645 16911 11648
rect 16853 11639 16911 11645
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 17034 11636 17040 11688
rect 17092 11676 17098 11688
rect 21266 11676 21272 11688
rect 17092 11648 21272 11676
rect 17092 11636 17098 11648
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 21542 11636 21548 11688
rect 21600 11676 21606 11688
rect 22005 11679 22063 11685
rect 22005 11676 22017 11679
rect 21600 11648 22017 11676
rect 21600 11636 21606 11648
rect 22005 11645 22017 11648
rect 22051 11645 22063 11679
rect 22005 11639 22063 11645
rect 22189 11679 22247 11685
rect 22189 11645 22201 11679
rect 22235 11676 22247 11679
rect 24136 11676 24164 11716
rect 26418 11704 26424 11716
rect 26476 11704 26482 11756
rect 26510 11704 26516 11756
rect 26568 11744 26574 11756
rect 28077 11747 28135 11753
rect 28077 11744 28089 11747
rect 26568 11716 28089 11744
rect 26568 11704 26574 11716
rect 28077 11713 28089 11716
rect 28123 11744 28135 11747
rect 29365 11747 29423 11753
rect 28123 11716 29224 11744
rect 28123 11713 28135 11716
rect 28077 11707 28135 11713
rect 22235 11648 24164 11676
rect 22235 11645 22247 11648
rect 22189 11639 22247 11645
rect 24210 11636 24216 11688
rect 24268 11676 24274 11688
rect 28810 11676 28816 11688
rect 24268 11648 28816 11676
rect 24268 11636 24274 11648
rect 28810 11636 28816 11648
rect 28868 11636 28874 11688
rect 13078 11608 13084 11620
rect 8352 11580 12434 11608
rect 13039 11580 13084 11608
rect 8352 11568 8358 11580
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 3326 11540 3332 11552
rect 3287 11512 3332 11540
rect 3326 11500 3332 11512
rect 3384 11500 3390 11552
rect 5718 11540 5724 11552
rect 5679 11512 5724 11540
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 7561 11543 7619 11549
rect 7561 11509 7573 11543
rect 7607 11540 7619 11543
rect 9950 11540 9956 11552
rect 7607 11512 9956 11540
rect 7607 11509 7619 11512
rect 7561 11503 7619 11509
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 12406 11540 12434 11580
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 15105 11611 15163 11617
rect 15105 11577 15117 11611
rect 15151 11608 15163 11611
rect 29089 11611 29147 11617
rect 29089 11608 29101 11611
rect 15151 11580 21956 11608
rect 15151 11577 15163 11580
rect 15105 11571 15163 11577
rect 12526 11540 12532 11552
rect 12406 11512 12532 11540
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 14274 11540 14280 11552
rect 13780 11512 14280 11540
rect 13780 11500 13786 11512
rect 14274 11500 14280 11512
rect 14332 11540 14338 11552
rect 17034 11540 17040 11552
rect 14332 11512 17040 11540
rect 14332 11500 14338 11512
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 18782 11540 18788 11552
rect 18743 11512 18788 11540
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 21818 11540 21824 11552
rect 21779 11512 21824 11540
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 21928 11540 21956 11580
rect 28460 11580 29101 11608
rect 24210 11540 24216 11552
rect 21928 11512 24216 11540
rect 24210 11500 24216 11512
rect 24268 11500 24274 11552
rect 24305 11543 24363 11549
rect 24305 11509 24317 11543
rect 24351 11540 24363 11543
rect 24946 11540 24952 11552
rect 24351 11512 24952 11540
rect 24351 11509 24363 11512
rect 24305 11503 24363 11509
rect 24946 11500 24952 11512
rect 25004 11500 25010 11552
rect 28460 11549 28488 11580
rect 29089 11577 29101 11580
rect 29135 11577 29147 11611
rect 29196 11608 29224 11716
rect 29365 11713 29377 11747
rect 29411 11744 29423 11747
rect 29914 11744 29920 11756
rect 29411 11716 29920 11744
rect 29411 11713 29423 11716
rect 29365 11707 29423 11713
rect 29914 11704 29920 11716
rect 29972 11704 29978 11756
rect 31110 11704 31116 11756
rect 31168 11744 31174 11756
rect 31478 11744 31484 11756
rect 31168 11716 31484 11744
rect 31168 11704 31174 11716
rect 31478 11704 31484 11716
rect 31536 11744 31542 11756
rect 32493 11747 32551 11753
rect 32493 11744 32505 11747
rect 31536 11716 32505 11744
rect 31536 11704 31542 11716
rect 32493 11713 32505 11716
rect 32539 11713 32551 11747
rect 32493 11707 32551 11713
rect 32674 11704 32680 11756
rect 32732 11744 32738 11756
rect 34517 11747 34575 11753
rect 34517 11744 34529 11747
rect 32732 11716 34529 11744
rect 32732 11704 32738 11716
rect 34517 11713 34529 11716
rect 34563 11713 34575 11747
rect 34517 11707 34575 11713
rect 34784 11747 34842 11753
rect 34784 11713 34796 11747
rect 34830 11744 34842 11747
rect 36170 11744 36176 11756
rect 34830 11716 36176 11744
rect 34830 11713 34842 11716
rect 34784 11707 34842 11713
rect 36170 11704 36176 11716
rect 36228 11704 36234 11756
rect 36354 11744 36360 11756
rect 36315 11716 36360 11744
rect 36354 11704 36360 11716
rect 36412 11704 36418 11756
rect 36449 11747 36507 11753
rect 36449 11713 36461 11747
rect 36495 11744 36507 11747
rect 36538 11744 36544 11756
rect 36495 11716 36544 11744
rect 36495 11713 36507 11716
rect 36449 11707 36507 11713
rect 36538 11704 36544 11716
rect 36596 11704 36602 11756
rect 42610 11704 42616 11756
rect 42668 11744 42674 11756
rect 42705 11747 42763 11753
rect 42705 11744 42717 11747
rect 42668 11716 42717 11744
rect 42668 11704 42674 11716
rect 42705 11713 42717 11716
rect 42751 11713 42763 11747
rect 42705 11707 42763 11713
rect 29270 11636 29276 11688
rect 29328 11676 29334 11688
rect 29454 11676 29460 11688
rect 29328 11648 29373 11676
rect 29415 11648 29460 11676
rect 29328 11636 29334 11648
rect 29454 11636 29460 11648
rect 29512 11636 29518 11688
rect 29549 11679 29607 11685
rect 29549 11645 29561 11679
rect 29595 11676 29607 11679
rect 29822 11676 29828 11688
rect 29595 11648 29828 11676
rect 29595 11645 29607 11648
rect 29549 11639 29607 11645
rect 29822 11636 29828 11648
rect 29880 11636 29886 11688
rect 36633 11679 36691 11685
rect 36633 11676 36645 11679
rect 35912 11648 36645 11676
rect 35912 11620 35940 11648
rect 36633 11645 36645 11648
rect 36679 11645 36691 11679
rect 36633 11639 36691 11645
rect 30098 11608 30104 11620
rect 29196 11580 30104 11608
rect 29089 11571 29147 11577
rect 30098 11568 30104 11580
rect 30156 11568 30162 11620
rect 32677 11611 32735 11617
rect 32677 11577 32689 11611
rect 32723 11608 32735 11611
rect 33594 11608 33600 11620
rect 32723 11580 33600 11608
rect 32723 11577 32735 11580
rect 32677 11571 32735 11577
rect 33594 11568 33600 11580
rect 33652 11568 33658 11620
rect 35894 11608 35900 11620
rect 35855 11580 35900 11608
rect 35894 11568 35900 11580
rect 35952 11568 35958 11620
rect 35986 11568 35992 11620
rect 36044 11608 36050 11620
rect 42518 11608 42524 11620
rect 36044 11580 42524 11608
rect 36044 11568 36050 11580
rect 42518 11568 42524 11580
rect 42576 11568 42582 11620
rect 28445 11543 28503 11549
rect 28445 11509 28457 11543
rect 28491 11509 28503 11543
rect 28626 11540 28632 11552
rect 28587 11512 28632 11540
rect 28445 11503 28503 11509
rect 28626 11500 28632 11512
rect 28684 11500 28690 11552
rect 29546 11500 29552 11552
rect 29604 11540 29610 11552
rect 30834 11540 30840 11552
rect 29604 11512 30840 11540
rect 29604 11500 29610 11512
rect 30834 11500 30840 11512
rect 30892 11500 30898 11552
rect 36538 11500 36544 11552
rect 36596 11540 36602 11552
rect 36596 11512 36641 11540
rect 36596 11500 36602 11512
rect 40310 11500 40316 11552
rect 40368 11540 40374 11552
rect 41046 11540 41052 11552
rect 40368 11512 41052 11540
rect 40368 11500 40374 11512
rect 41046 11500 41052 11512
rect 41104 11500 41110 11552
rect 42720 11540 42748 11707
rect 43180 11676 43208 11784
rect 43254 11704 43260 11756
rect 43312 11744 43318 11756
rect 43605 11747 43663 11753
rect 43605 11744 43617 11747
rect 43312 11716 43617 11744
rect 43312 11704 43318 11716
rect 43605 11713 43617 11716
rect 43651 11713 43663 11747
rect 43732 11744 43760 11784
rect 43990 11772 43996 11824
rect 44048 11812 44054 11824
rect 45434 11815 45492 11821
rect 45434 11812 45446 11815
rect 44048 11784 45446 11812
rect 44048 11772 44054 11784
rect 45434 11781 45446 11784
rect 45480 11781 45492 11815
rect 45572 11812 45600 11852
rect 46566 11840 46572 11852
rect 46624 11840 46630 11892
rect 48041 11883 48099 11889
rect 48041 11849 48053 11883
rect 48087 11880 48099 11883
rect 48406 11880 48412 11892
rect 48087 11852 48412 11880
rect 48087 11849 48099 11852
rect 48041 11843 48099 11849
rect 48406 11840 48412 11852
rect 48464 11880 48470 11892
rect 48682 11880 48688 11892
rect 48464 11852 48688 11880
rect 48464 11840 48470 11852
rect 48682 11840 48688 11852
rect 48740 11840 48746 11892
rect 55398 11880 55404 11892
rect 54036 11852 55404 11880
rect 53926 11812 53932 11824
rect 45572 11784 51672 11812
rect 53887 11784 53932 11812
rect 45434 11775 45492 11781
rect 45189 11747 45247 11753
rect 45189 11744 45201 11747
rect 43732 11716 45201 11744
rect 43605 11707 43663 11713
rect 45189 11713 45201 11716
rect 45235 11744 45247 11747
rect 46014 11744 46020 11756
rect 45235 11716 46020 11744
rect 45235 11713 45247 11716
rect 45189 11707 45247 11713
rect 46014 11704 46020 11716
rect 46072 11704 46078 11756
rect 46566 11704 46572 11756
rect 46624 11744 46630 11756
rect 47949 11747 48007 11753
rect 47949 11744 47961 11747
rect 46624 11716 47961 11744
rect 46624 11704 46630 11716
rect 47949 11713 47961 11716
rect 47995 11744 48007 11747
rect 48774 11744 48780 11756
rect 47995 11716 48780 11744
rect 47995 11713 48007 11716
rect 47949 11707 48007 11713
rect 48774 11704 48780 11716
rect 48832 11704 48838 11756
rect 49053 11747 49111 11753
rect 49053 11713 49065 11747
rect 49099 11713 49111 11747
rect 51442 11744 51448 11756
rect 51403 11716 51448 11744
rect 49053 11707 49111 11713
rect 43349 11679 43407 11685
rect 43349 11676 43361 11679
rect 43180 11648 43361 11676
rect 43349 11645 43361 11648
rect 43395 11645 43407 11679
rect 43349 11639 43407 11645
rect 48590 11636 48596 11688
rect 48648 11676 48654 11688
rect 49068 11676 49096 11707
rect 51442 11704 51448 11716
rect 51500 11704 51506 11756
rect 51534 11676 51540 11688
rect 48648 11648 51540 11676
rect 48648 11636 48654 11648
rect 51534 11636 51540 11648
rect 51592 11636 51598 11688
rect 51644 11676 51672 11784
rect 53926 11772 53932 11784
rect 53984 11772 53990 11824
rect 51994 11704 52000 11756
rect 52052 11744 52058 11756
rect 54036 11744 54064 11852
rect 55398 11840 55404 11852
rect 55456 11840 55462 11892
rect 56045 11883 56103 11889
rect 56045 11849 56057 11883
rect 56091 11849 56103 11883
rect 56045 11843 56103 11849
rect 54113 11815 54171 11821
rect 54113 11781 54125 11815
rect 54159 11812 54171 11815
rect 55122 11812 55128 11824
rect 54159 11784 55128 11812
rect 54159 11781 54171 11784
rect 54113 11775 54171 11781
rect 55122 11772 55128 11784
rect 55180 11812 55186 11824
rect 56060 11812 56088 11843
rect 55180 11784 56088 11812
rect 55180 11772 55186 11784
rect 54205 11747 54263 11753
rect 54205 11744 54217 11747
rect 52052 11716 54217 11744
rect 52052 11704 52058 11716
rect 54205 11713 54217 11716
rect 54251 11713 54263 11747
rect 54921 11747 54979 11753
rect 54921 11744 54933 11747
rect 54205 11707 54263 11713
rect 54404 11716 54933 11744
rect 51721 11679 51779 11685
rect 51721 11676 51733 11679
rect 51644 11648 51733 11676
rect 51721 11645 51733 11648
rect 51767 11645 51779 11679
rect 51721 11639 51779 11645
rect 51350 11568 51356 11620
rect 51408 11608 51414 11620
rect 51629 11611 51687 11617
rect 51629 11608 51641 11611
rect 51408 11580 51641 11608
rect 51408 11568 51414 11580
rect 51629 11577 51641 11580
rect 51675 11577 51687 11611
rect 51629 11571 51687 11577
rect 44729 11543 44787 11549
rect 44729 11540 44741 11543
rect 42720 11512 44741 11540
rect 44729 11509 44741 11512
rect 44775 11509 44787 11543
rect 48682 11540 48688 11552
rect 48643 11512 48688 11540
rect 44729 11503 44787 11509
rect 48682 11500 48688 11512
rect 48740 11540 48746 11552
rect 48866 11540 48872 11552
rect 48740 11512 48872 11540
rect 48740 11500 48746 11512
rect 48866 11500 48872 11512
rect 48924 11500 48930 11552
rect 51736 11540 51764 11639
rect 53929 11611 53987 11617
rect 53929 11577 53941 11611
rect 53975 11608 53987 11611
rect 54404 11608 54432 11716
rect 54921 11713 54933 11716
rect 54967 11713 54979 11747
rect 54921 11707 54979 11713
rect 54662 11676 54668 11688
rect 54623 11648 54668 11676
rect 54662 11636 54668 11648
rect 54720 11636 54726 11688
rect 53975 11580 54432 11608
rect 53975 11577 53987 11580
rect 53929 11571 53987 11577
rect 55582 11540 55588 11552
rect 51736 11512 55588 11540
rect 55582 11500 55588 11512
rect 55640 11500 55646 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 5442 11336 5448 11348
rect 5403 11308 5448 11336
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 8018 11296 8024 11348
rect 8076 11336 8082 11348
rect 9493 11339 9551 11345
rect 9493 11336 9505 11339
rect 8076 11308 9505 11336
rect 8076 11296 8082 11308
rect 9493 11305 9505 11308
rect 9539 11305 9551 11339
rect 9493 11299 9551 11305
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 12897 11339 12955 11345
rect 12897 11336 12909 11339
rect 12492 11308 12909 11336
rect 12492 11296 12498 11308
rect 12897 11305 12909 11308
rect 12943 11305 12955 11339
rect 12897 11299 12955 11305
rect 14093 11339 14151 11345
rect 14093 11305 14105 11339
rect 14139 11336 14151 11339
rect 14366 11336 14372 11348
rect 14139 11308 14372 11336
rect 14139 11305 14151 11308
rect 14093 11299 14151 11305
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 16850 11296 16856 11348
rect 16908 11336 16914 11348
rect 17589 11339 17647 11345
rect 17589 11336 17601 11339
rect 16908 11308 17601 11336
rect 16908 11296 16914 11308
rect 17589 11305 17601 11308
rect 17635 11305 17647 11339
rect 21542 11336 21548 11348
rect 21503 11308 21548 11336
rect 17589 11299 17647 11305
rect 21542 11296 21548 11308
rect 21600 11296 21606 11348
rect 23385 11339 23443 11345
rect 23385 11305 23397 11339
rect 23431 11305 23443 11339
rect 23566 11336 23572 11348
rect 23527 11308 23572 11336
rect 23385 11299 23443 11305
rect 12345 11271 12403 11277
rect 12345 11237 12357 11271
rect 12391 11268 12403 11271
rect 12618 11268 12624 11280
rect 12391 11240 12624 11268
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 13170 11268 13176 11280
rect 12820 11240 13176 11268
rect 2038 11160 2044 11212
rect 2096 11200 2102 11212
rect 2590 11200 2596 11212
rect 2096 11172 2596 11200
rect 2096 11160 2102 11172
rect 2590 11160 2596 11172
rect 2648 11200 2654 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 2648 11172 4077 11200
rect 2648 11160 2654 11172
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 10870 11160 10876 11212
rect 10928 11200 10934 11212
rect 12820 11200 12848 11240
rect 13170 11228 13176 11240
rect 13228 11228 13234 11280
rect 13357 11271 13415 11277
rect 13357 11237 13369 11271
rect 13403 11268 13415 11271
rect 15654 11268 15660 11280
rect 13403 11240 15660 11268
rect 13403 11237 13415 11240
rect 13357 11231 13415 11237
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 15930 11228 15936 11280
rect 15988 11268 15994 11280
rect 22922 11268 22928 11280
rect 15988 11240 22928 11268
rect 15988 11228 15994 11240
rect 22922 11228 22928 11240
rect 22980 11228 22986 11280
rect 23017 11271 23075 11277
rect 23017 11237 23029 11271
rect 23063 11268 23075 11271
rect 23106 11268 23112 11280
rect 23063 11240 23112 11268
rect 23063 11237 23075 11240
rect 23017 11231 23075 11237
rect 23106 11228 23112 11240
rect 23164 11228 23170 11280
rect 23400 11268 23428 11299
rect 23566 11296 23572 11308
rect 23624 11296 23630 11348
rect 34790 11336 34796 11348
rect 34751 11308 34796 11336
rect 34790 11296 34796 11308
rect 34848 11296 34854 11348
rect 35176 11308 35388 11336
rect 24486 11268 24492 11280
rect 23400 11240 24492 11268
rect 24486 11228 24492 11240
rect 24544 11228 24550 11280
rect 26878 11228 26884 11280
rect 26936 11268 26942 11280
rect 35066 11268 35072 11280
rect 26936 11240 35072 11268
rect 26936 11228 26942 11240
rect 35066 11228 35072 11240
rect 35124 11228 35130 11280
rect 10928 11172 12848 11200
rect 13081 11203 13139 11209
rect 10928 11160 10934 11172
rect 13081 11169 13093 11203
rect 13127 11200 13139 11203
rect 13446 11200 13452 11212
rect 13127 11172 13452 11200
rect 13127 11169 13139 11172
rect 13081 11163 13139 11169
rect 2130 11092 2136 11144
rect 2188 11132 2194 11144
rect 2685 11135 2743 11141
rect 2685 11132 2697 11135
rect 2188 11104 2697 11132
rect 2188 11092 2194 11104
rect 2685 11101 2697 11104
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 9950 11092 9956 11144
rect 10008 11132 10014 11144
rect 10045 11135 10103 11141
rect 10045 11132 10057 11135
rect 10008 11104 10057 11132
rect 10008 11092 10014 11104
rect 10045 11101 10057 11104
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 11514 11132 11520 11144
rect 10284 11104 11520 11132
rect 10284 11092 10290 11104
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12250 11132 12256 11144
rect 12207 11104 12256 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 13096 11132 13124 11163
rect 13446 11160 13452 11172
rect 13504 11200 13510 11212
rect 16301 11203 16359 11209
rect 13504 11172 14320 11200
rect 13504 11160 13510 11172
rect 12676 11104 13124 11132
rect 13173 11135 13231 11141
rect 12676 11092 12682 11104
rect 13173 11101 13185 11135
rect 13219 11132 13231 11135
rect 13722 11132 13728 11144
rect 13219 11104 13728 11132
rect 13219 11101 13231 11104
rect 13173 11095 13231 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 14090 11132 14096 11144
rect 14051 11104 14096 11132
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 14292 11141 14320 11172
rect 16301 11169 16313 11203
rect 16347 11200 16359 11203
rect 16390 11200 16396 11212
rect 16347 11172 16396 11200
rect 16347 11169 16359 11172
rect 16301 11163 16359 11169
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 16577 11203 16635 11209
rect 16577 11169 16589 11203
rect 16623 11200 16635 11203
rect 17126 11200 17132 11212
rect 16623 11172 17132 11200
rect 16623 11169 16635 11172
rect 16577 11163 16635 11169
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 18046 11200 18052 11212
rect 18007 11172 18052 11200
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 22554 11200 22560 11212
rect 22204 11172 22560 11200
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 16908 11104 17785 11132
rect 16908 11092 16914 11104
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 17865 11135 17923 11141
rect 17865 11101 17877 11135
rect 17911 11101 17923 11135
rect 17865 11095 17923 11101
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11132 18015 11135
rect 19426 11132 19432 11144
rect 18003 11104 19432 11132
rect 18003 11101 18015 11104
rect 17957 11095 18015 11101
rect 1854 11064 1860 11076
rect 1815 11036 1860 11064
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 2041 11067 2099 11073
rect 2041 11033 2053 11067
rect 2087 11064 2099 11067
rect 2590 11064 2596 11076
rect 2087 11036 2596 11064
rect 2087 11033 2099 11036
rect 2041 11027 2099 11033
rect 2590 11024 2596 11036
rect 2648 11024 2654 11076
rect 4332 11067 4390 11073
rect 4332 11033 4344 11067
rect 4378 11064 4390 11067
rect 4890 11064 4896 11076
rect 4378 11036 4896 11064
rect 4378 11033 4390 11036
rect 4332 11027 4390 11033
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 7926 11064 7932 11076
rect 6972 11036 7932 11064
rect 6972 11024 6978 11036
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 9398 11064 9404 11076
rect 9359 11036 9404 11064
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 9968 11036 10272 11064
rect 2498 10996 2504 11008
rect 2459 10968 2504 10996
rect 2498 10956 2504 10968
rect 2556 10956 2562 11008
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 9968 10996 9996 11036
rect 10134 10996 10140 11008
rect 7064 10968 9996 10996
rect 10095 10968 10140 10996
rect 7064 10956 7070 10968
rect 10134 10956 10140 10968
rect 10192 10956 10198 11008
rect 10244 10996 10272 11036
rect 11790 11024 11796 11076
rect 11848 11064 11854 11076
rect 12894 11064 12900 11076
rect 11848 11036 12900 11064
rect 11848 11024 11854 11036
rect 12894 11024 12900 11036
rect 12952 11024 12958 11076
rect 16482 11024 16488 11076
rect 16540 11064 16546 11076
rect 17880 11064 17908 11095
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 22204 11141 22232 11172
rect 22554 11160 22560 11172
rect 22612 11160 22618 11212
rect 26050 11160 26056 11212
rect 26108 11200 26114 11212
rect 29546 11200 29552 11212
rect 26108 11172 29552 11200
rect 26108 11160 26114 11172
rect 29546 11160 29552 11172
rect 29604 11160 29610 11212
rect 29914 11200 29920 11212
rect 29702 11172 29920 11200
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11101 22247 11135
rect 22189 11095 22247 11101
rect 22278 11092 22284 11144
rect 22336 11132 22342 11144
rect 22465 11135 22523 11141
rect 22465 11132 22477 11135
rect 22336 11104 22477 11132
rect 22336 11092 22342 11104
rect 22465 11101 22477 11104
rect 22511 11101 22523 11135
rect 22572 11132 22600 11160
rect 24765 11135 24823 11141
rect 22572 11104 23520 11132
rect 22465 11095 22523 11101
rect 21174 11064 21180 11076
rect 16540 11036 17908 11064
rect 21135 11036 21180 11064
rect 16540 11024 16546 11036
rect 21174 11024 21180 11036
rect 21232 11024 21238 11076
rect 21361 11067 21419 11073
rect 21361 11033 21373 11067
rect 21407 11064 21419 11067
rect 22005 11067 22063 11073
rect 21407 11036 21772 11064
rect 21407 11033 21419 11036
rect 21361 11027 21419 11033
rect 21744 11008 21772 11036
rect 22005 11033 22017 11067
rect 22051 11064 22063 11067
rect 23385 11067 23443 11073
rect 23385 11064 23397 11067
rect 22051 11036 23397 11064
rect 22051 11033 22063 11036
rect 22005 11027 22063 11033
rect 23385 11033 23397 11036
rect 23431 11033 23443 11067
rect 23492 11064 23520 11104
rect 24765 11101 24777 11135
rect 24811 11132 24823 11135
rect 27430 11132 27436 11144
rect 24811 11104 27436 11132
rect 24811 11101 24823 11104
rect 24765 11095 24823 11101
rect 27430 11092 27436 11104
rect 27488 11092 27494 11144
rect 28169 11135 28227 11141
rect 28169 11101 28181 11135
rect 28215 11132 28227 11135
rect 28626 11132 28632 11144
rect 28215 11104 28632 11132
rect 28215 11101 28227 11104
rect 28169 11095 28227 11101
rect 28626 11092 28632 11104
rect 28684 11092 28690 11144
rect 29702 11122 29730 11172
rect 29914 11160 29920 11172
rect 29972 11200 29978 11212
rect 35176 11200 35204 11308
rect 35253 11271 35311 11277
rect 35253 11237 35265 11271
rect 35299 11237 35311 11271
rect 35360 11268 35388 11308
rect 35434 11296 35440 11348
rect 35492 11336 35498 11348
rect 36081 11339 36139 11345
rect 36081 11336 36093 11339
rect 35492 11308 36093 11336
rect 35492 11296 35498 11308
rect 36081 11305 36093 11308
rect 36127 11305 36139 11339
rect 36081 11299 36139 11305
rect 36170 11296 36176 11348
rect 36228 11336 36234 11348
rect 36228 11308 36273 11336
rect 36228 11296 36234 11308
rect 36814 11296 36820 11348
rect 36872 11336 36878 11348
rect 43070 11336 43076 11348
rect 36872 11308 43076 11336
rect 36872 11296 36878 11308
rect 43070 11296 43076 11308
rect 43128 11296 43134 11348
rect 43254 11336 43260 11348
rect 43215 11308 43260 11336
rect 43254 11296 43260 11308
rect 43312 11296 43318 11348
rect 44450 11296 44456 11348
rect 44508 11336 44514 11348
rect 47765 11339 47823 11345
rect 47765 11336 47777 11339
rect 44508 11308 47777 11336
rect 44508 11296 44514 11308
rect 47765 11305 47777 11308
rect 47811 11305 47823 11339
rect 47765 11299 47823 11305
rect 39942 11268 39948 11280
rect 35360 11240 39948 11268
rect 35253 11231 35311 11237
rect 29972 11172 35204 11200
rect 29972 11160 29978 11172
rect 29702 11094 29776 11122
rect 23492 11036 24808 11064
rect 23385 11027 23443 11033
rect 15562 10996 15568 11008
rect 10244 10968 15568 10996
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 21726 10956 21732 11008
rect 21784 10996 21790 11008
rect 22373 10999 22431 11005
rect 22373 10996 22385 10999
rect 21784 10968 22385 10996
rect 21784 10956 21790 10968
rect 22373 10965 22385 10968
rect 22419 10965 22431 10999
rect 24780 10996 24808 11036
rect 24854 11024 24860 11076
rect 24912 11064 24918 11076
rect 25010 11067 25068 11073
rect 25010 11064 25022 11067
rect 24912 11036 25022 11064
rect 24912 11024 24918 11036
rect 25010 11033 25022 11036
rect 25056 11033 25068 11067
rect 25010 11027 25068 11033
rect 25222 11024 25228 11076
rect 25280 11064 25286 11076
rect 28353 11067 28411 11073
rect 28353 11064 28365 11067
rect 25280 11036 28365 11064
rect 25280 11024 25286 11036
rect 28353 11033 28365 11036
rect 28399 11033 28411 11067
rect 28534 11064 28540 11076
rect 28495 11036 28540 11064
rect 28353 11027 28411 11033
rect 28534 11024 28540 11036
rect 28592 11024 28598 11076
rect 29454 11024 29460 11076
rect 29512 11064 29518 11076
rect 29549 11067 29607 11073
rect 29549 11064 29561 11067
rect 29512 11036 29561 11064
rect 29512 11024 29518 11036
rect 29549 11033 29561 11036
rect 29595 11033 29607 11067
rect 29549 11027 29607 11033
rect 29748 11005 29776 11094
rect 29822 11092 29828 11144
rect 29880 11132 29886 11144
rect 30098 11132 30104 11144
rect 29880 11104 29925 11132
rect 30059 11104 30104 11132
rect 29880 11092 29886 11104
rect 30098 11092 30104 11104
rect 30156 11092 30162 11144
rect 33778 11092 33784 11144
rect 33836 11132 33842 11144
rect 34701 11135 34759 11141
rect 34701 11132 34713 11135
rect 33836 11104 34713 11132
rect 33836 11092 33842 11104
rect 34701 11101 34713 11104
rect 34747 11101 34759 11135
rect 34701 11095 34759 11101
rect 35069 11135 35127 11141
rect 35069 11101 35081 11135
rect 35115 11101 35127 11135
rect 35268 11132 35296 11231
rect 39942 11228 39948 11240
rect 40000 11228 40006 11280
rect 40586 11228 40592 11280
rect 40644 11268 40650 11280
rect 40773 11271 40831 11277
rect 40773 11268 40785 11271
rect 40644 11240 40785 11268
rect 40644 11228 40650 11240
rect 40773 11237 40785 11240
rect 40819 11237 40831 11271
rect 40773 11231 40831 11237
rect 36538 11200 36544 11212
rect 36004 11172 36544 11200
rect 35268 11124 35664 11132
rect 35702 11127 35760 11133
rect 35702 11124 35714 11127
rect 35268 11104 35714 11124
rect 35069 11095 35127 11101
rect 35636 11096 35714 11104
rect 29914 11064 29920 11076
rect 29875 11036 29920 11064
rect 29914 11024 29920 11036
rect 29972 11024 29978 11076
rect 35084 11064 35112 11095
rect 35702 11093 35714 11096
rect 35748 11093 35760 11127
rect 35702 11087 35760 11093
rect 35805 11067 35863 11073
rect 35084 11036 35664 11064
rect 26145 10999 26203 11005
rect 26145 10996 26157 10999
rect 24780 10968 26157 10996
rect 22373 10959 22431 10965
rect 26145 10965 26157 10968
rect 26191 10965 26203 10999
rect 26145 10959 26203 10965
rect 29733 10999 29791 11005
rect 29733 10965 29745 10999
rect 29779 10965 29791 10999
rect 29733 10959 29791 10965
rect 34146 10956 34152 11008
rect 34204 10996 34210 11008
rect 35434 10996 35440 11008
rect 34204 10968 35440 10996
rect 34204 10956 34210 10968
rect 35434 10956 35440 10968
rect 35492 10956 35498 11008
rect 35636 10996 35664 11036
rect 35805 11033 35817 11067
rect 35851 11064 35863 11067
rect 36004 11064 36032 11172
rect 36538 11160 36544 11172
rect 36596 11160 36602 11212
rect 36648 11172 37044 11200
rect 36170 11132 36176 11144
rect 36131 11104 36176 11132
rect 36170 11092 36176 11104
rect 36228 11132 36234 11144
rect 36648 11132 36676 11172
rect 36228 11104 36676 11132
rect 36725 11135 36783 11141
rect 36228 11092 36234 11104
rect 36725 11101 36737 11135
rect 36771 11132 36783 11135
rect 36814 11132 36820 11144
rect 36771 11104 36820 11132
rect 36771 11101 36783 11104
rect 36725 11095 36783 11101
rect 36814 11092 36820 11104
rect 36872 11092 36878 11144
rect 36909 11135 36967 11141
rect 36909 11101 36921 11135
rect 36955 11101 36967 11135
rect 37016 11132 37044 11172
rect 38378 11160 38384 11212
rect 38436 11200 38442 11212
rect 42889 11203 42947 11209
rect 42889 11200 42901 11203
rect 38436 11172 42901 11200
rect 38436 11160 38442 11172
rect 42889 11169 42901 11172
rect 42935 11169 42947 11203
rect 43622 11200 43628 11212
rect 42889 11163 42947 11169
rect 42996 11172 43628 11200
rect 38930 11132 38936 11144
rect 37016 11104 38936 11132
rect 36909 11095 36967 11101
rect 35851 11036 36032 11064
rect 35851 11033 35863 11036
rect 35805 11027 35863 11033
rect 36078 11024 36084 11076
rect 36136 11064 36142 11076
rect 36354 11064 36360 11076
rect 36136 11036 36360 11064
rect 36136 11024 36142 11036
rect 36354 11024 36360 11036
rect 36412 11064 36418 11076
rect 36924 11064 36952 11095
rect 38930 11092 38936 11104
rect 38988 11092 38994 11144
rect 40862 11092 40868 11144
rect 40920 11132 40926 11144
rect 40957 11135 41015 11141
rect 40957 11132 40969 11135
rect 40920 11104 40969 11132
rect 40920 11092 40926 11104
rect 40957 11101 40969 11104
rect 41003 11101 41015 11135
rect 40957 11095 41015 11101
rect 41046 11092 41052 11144
rect 41104 11132 41110 11144
rect 42521 11135 42579 11141
rect 41104 11104 41149 11132
rect 41104 11092 41110 11104
rect 42521 11101 42533 11135
rect 42567 11101 42579 11135
rect 42702 11132 42708 11144
rect 42663 11104 42708 11132
rect 42521 11095 42579 11101
rect 36412 11036 36952 11064
rect 36412 11024 36418 11036
rect 37090 11024 37096 11076
rect 37148 11064 37154 11076
rect 40770 11064 40776 11076
rect 37148 11036 38654 11064
rect 40731 11036 40776 11064
rect 37148 11024 37154 11036
rect 35710 10996 35716 11008
rect 35636 10968 35716 10996
rect 35710 10956 35716 10968
rect 35768 10956 35774 11008
rect 35923 10999 35981 11005
rect 35923 10965 35935 10999
rect 35969 10996 35981 10999
rect 36170 10996 36176 11008
rect 35969 10968 36176 10996
rect 35969 10965 35981 10968
rect 35923 10959 35981 10965
rect 36170 10956 36176 10968
rect 36228 10956 36234 11008
rect 36538 10956 36544 11008
rect 36596 10996 36602 11008
rect 36817 10999 36875 11005
rect 36817 10996 36829 10999
rect 36596 10968 36829 10996
rect 36596 10956 36602 10968
rect 36817 10965 36829 10968
rect 36863 10965 36875 10999
rect 38626 10996 38654 11036
rect 40770 11024 40776 11036
rect 40828 11024 40834 11076
rect 42536 11064 42564 11095
rect 42702 11092 42708 11104
rect 42760 11092 42766 11144
rect 42797 11135 42855 11141
rect 42797 11101 42809 11135
rect 42843 11132 42855 11135
rect 42996 11132 43024 11172
rect 43622 11160 43628 11172
rect 43680 11160 43686 11212
rect 42843 11104 43024 11132
rect 42843 11101 42855 11104
rect 42797 11095 42855 11101
rect 43070 11092 43076 11144
rect 43128 11132 43134 11144
rect 43714 11132 43720 11144
rect 43128 11104 43720 11132
rect 43128 11092 43134 11104
rect 43714 11092 43720 11104
rect 43772 11092 43778 11144
rect 47670 11132 47676 11144
rect 47631 11104 47676 11132
rect 47670 11092 47676 11104
rect 47728 11092 47734 11144
rect 43162 11064 43168 11076
rect 42536 11036 43168 11064
rect 42536 10996 42564 11036
rect 43162 11024 43168 11036
rect 43220 11024 43226 11076
rect 47780 11064 47808 11299
rect 48590 11268 48596 11280
rect 48551 11240 48596 11268
rect 48590 11228 48596 11240
rect 48648 11228 48654 11280
rect 51353 11271 51411 11277
rect 51353 11237 51365 11271
rect 51399 11268 51411 11271
rect 51626 11268 51632 11280
rect 51399 11240 51632 11268
rect 51399 11237 51411 11240
rect 51353 11231 51411 11237
rect 51626 11228 51632 11240
rect 51684 11228 51690 11280
rect 48406 11132 48412 11144
rect 48367 11104 48412 11132
rect 48406 11092 48412 11104
rect 48464 11092 48470 11144
rect 48501 11135 48559 11141
rect 48501 11101 48513 11135
rect 48547 11101 48559 11135
rect 51350 11132 51356 11144
rect 51311 11104 51356 11132
rect 48501 11095 48559 11101
rect 48516 11064 48544 11095
rect 51350 11092 51356 11104
rect 51408 11092 51414 11144
rect 51534 11092 51540 11144
rect 51592 11132 51598 11144
rect 51629 11135 51687 11141
rect 51629 11132 51641 11135
rect 51592 11104 51641 11132
rect 51592 11092 51598 11104
rect 51629 11101 51641 11104
rect 51675 11101 51687 11135
rect 51629 11095 51687 11101
rect 47780 11036 48544 11064
rect 38626 10968 42564 10996
rect 36817 10959 36875 10965
rect 51442 10956 51448 11008
rect 51500 10996 51506 11008
rect 51537 10999 51595 11005
rect 51537 10996 51549 10999
rect 51500 10968 51549 10996
rect 51500 10956 51506 10968
rect 51537 10965 51549 10968
rect 51583 10965 51595 10999
rect 51537 10959 51595 10965
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 4890 10792 4896 10804
rect 4851 10764 4896 10792
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5442 10792 5448 10804
rect 5307 10764 5448 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 12802 10792 12808 10804
rect 7576 10764 12808 10792
rect 2308 10727 2366 10733
rect 2308 10693 2320 10727
rect 2354 10724 2366 10727
rect 2498 10724 2504 10736
rect 2354 10696 2504 10724
rect 2354 10693 2366 10696
rect 2308 10687 2366 10693
rect 2498 10684 2504 10696
rect 2556 10684 2562 10736
rect 2590 10684 2596 10736
rect 2648 10724 2654 10736
rect 7576 10724 7604 10764
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 12989 10795 13047 10801
rect 12989 10761 13001 10795
rect 13035 10792 13047 10795
rect 13262 10792 13268 10804
rect 13035 10764 13268 10792
rect 13035 10761 13047 10764
rect 12989 10755 13047 10761
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 15562 10792 15568 10804
rect 15523 10764 15568 10792
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 19521 10795 19579 10801
rect 19521 10761 19533 10795
rect 19567 10761 19579 10795
rect 19521 10755 19579 10761
rect 21269 10795 21327 10801
rect 21269 10761 21281 10795
rect 21315 10792 21327 10795
rect 22094 10792 22100 10804
rect 21315 10764 22100 10792
rect 21315 10761 21327 10764
rect 21269 10755 21327 10761
rect 2648 10696 7604 10724
rect 9484 10727 9542 10733
rect 2648 10684 2654 10696
rect 9484 10693 9496 10727
rect 9530 10724 9542 10727
rect 10134 10724 10140 10736
rect 9530 10696 10140 10724
rect 9530 10693 9542 10696
rect 9484 10687 9542 10693
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 14734 10724 14740 10736
rect 12820 10696 14740 10724
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 5074 10656 5080 10668
rect 5035 10628 5080 10656
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 5718 10656 5724 10668
rect 5399 10628 5724 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 7190 10656 7196 10668
rect 7151 10628 7196 10656
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 7340 10628 7389 10656
rect 7340 10616 7346 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 8018 10656 8024 10668
rect 7515 10628 8024 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 11790 10656 11796 10668
rect 9140 10628 11796 10656
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10588 7067 10591
rect 9140 10588 9168 10628
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 12158 10616 12164 10668
rect 12216 10656 12222 10668
rect 12345 10659 12403 10665
rect 12345 10656 12357 10659
rect 12216 10628 12357 10656
rect 12216 10616 12222 10628
rect 12345 10625 12357 10628
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 7055 10560 9168 10588
rect 9217 10591 9275 10597
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 9217 10557 9229 10591
rect 9263 10557 9275 10591
rect 11514 10588 11520 10600
rect 11475 10560 11520 10588
rect 9217 10551 9275 10557
rect 7285 10523 7343 10529
rect 7285 10489 7297 10523
rect 7331 10520 7343 10523
rect 7466 10520 7472 10532
rect 7331 10492 7472 10520
rect 7331 10489 7343 10492
rect 7285 10483 7343 10489
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 1394 10452 1400 10464
rect 1355 10424 1400 10452
rect 1394 10412 1400 10424
rect 1452 10412 1458 10464
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 9232 10452 9260 10551
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 12069 10591 12127 10597
rect 12069 10557 12081 10591
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 10594 10520 10600 10532
rect 10507 10492 10600 10520
rect 10594 10480 10600 10492
rect 10652 10520 10658 10532
rect 12084 10520 12112 10551
rect 12250 10548 12256 10600
rect 12308 10588 12314 10600
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12308 10560 12541 10588
rect 12308 10548 12314 10560
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 10652 10492 12112 10520
rect 10652 10480 10658 10492
rect 12342 10480 12348 10532
rect 12400 10520 12406 10532
rect 12820 10520 12848 10696
rect 12894 10616 12900 10668
rect 12952 10656 12958 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12952 10628 13001 10656
rect 12952 10616 12958 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 13446 10656 13452 10668
rect 12989 10619 13047 10625
rect 13188 10628 13452 10656
rect 13081 10591 13139 10597
rect 13081 10557 13093 10591
rect 13127 10588 13139 10591
rect 13188 10588 13216 10628
rect 13446 10616 13452 10628
rect 13504 10616 13510 10668
rect 13740 10665 13768 10696
rect 14734 10684 14740 10696
rect 14792 10684 14798 10736
rect 17862 10724 17868 10736
rect 15856 10696 17868 10724
rect 15856 10665 15884 10696
rect 17862 10684 17868 10696
rect 17920 10684 17926 10736
rect 18408 10727 18466 10733
rect 18408 10693 18420 10727
rect 18454 10724 18466 10727
rect 18782 10724 18788 10736
rect 18454 10696 18788 10724
rect 18454 10693 18466 10696
rect 18408 10687 18466 10693
rect 18782 10684 18788 10696
rect 18840 10684 18846 10736
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10625 13783 10659
rect 13725 10619 13783 10625
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 16758 10656 16764 10668
rect 16071 10628 16764 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 16850 10616 16856 10668
rect 16908 10656 16914 10668
rect 17037 10659 17095 10665
rect 16908 10628 16953 10656
rect 16908 10616 16914 10628
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 19150 10656 19156 10668
rect 17083 10628 19156 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 19150 10616 19156 10628
rect 19208 10656 19214 10668
rect 19536 10656 19564 10755
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 22481 10795 22539 10801
rect 22481 10792 22493 10795
rect 22204 10764 22493 10792
rect 22204 10736 22232 10764
rect 22481 10761 22493 10764
rect 22527 10761 22539 10795
rect 22481 10755 22539 10761
rect 22649 10795 22707 10801
rect 22649 10761 22661 10795
rect 22695 10792 22707 10795
rect 23106 10792 23112 10804
rect 22695 10764 23112 10792
rect 22695 10761 22707 10764
rect 22649 10755 22707 10761
rect 23106 10752 23112 10764
rect 23164 10752 23170 10804
rect 24673 10795 24731 10801
rect 24673 10761 24685 10795
rect 24719 10792 24731 10795
rect 24854 10792 24860 10804
rect 24719 10764 24860 10792
rect 24719 10761 24731 10764
rect 24673 10755 24731 10761
rect 24854 10752 24860 10764
rect 24912 10752 24918 10804
rect 40310 10792 40316 10804
rect 40271 10764 40316 10792
rect 40310 10752 40316 10764
rect 40368 10752 40374 10804
rect 40405 10795 40463 10801
rect 40405 10761 40417 10795
rect 40451 10792 40463 10795
rect 40862 10792 40868 10804
rect 40451 10764 40868 10792
rect 40451 10761 40463 10764
rect 40405 10755 40463 10761
rect 40862 10752 40868 10764
rect 40920 10752 40926 10804
rect 48314 10752 48320 10804
rect 48372 10792 48378 10804
rect 49329 10795 49387 10801
rect 49329 10792 49341 10795
rect 48372 10764 49341 10792
rect 48372 10752 48378 10764
rect 49329 10761 49341 10764
rect 49375 10761 49387 10795
rect 49329 10755 49387 10761
rect 21174 10724 21180 10736
rect 21087 10696 21180 10724
rect 21100 10665 21128 10696
rect 21174 10684 21180 10696
rect 21232 10724 21238 10736
rect 22186 10724 22192 10736
rect 21232 10696 22192 10724
rect 21232 10684 21238 10696
rect 22186 10684 22192 10696
rect 22244 10684 22250 10736
rect 22278 10684 22284 10736
rect 22336 10724 22342 10736
rect 38654 10724 38660 10736
rect 22336 10696 22600 10724
rect 38615 10696 38660 10724
rect 22336 10684 22342 10696
rect 22572 10668 22600 10696
rect 38654 10684 38660 10696
rect 38712 10684 38718 10736
rect 38948 10696 40356 10724
rect 19208 10628 19564 10656
rect 21085 10659 21143 10665
rect 19208 10616 19214 10628
rect 21085 10625 21097 10659
rect 21131 10625 21143 10659
rect 21085 10619 21143 10625
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10656 21327 10659
rect 21726 10656 21732 10668
rect 21315 10628 21732 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 21726 10616 21732 10628
rect 21784 10616 21790 10668
rect 22554 10616 22560 10668
rect 22612 10616 22618 10668
rect 24857 10659 24915 10665
rect 24857 10625 24869 10659
rect 24903 10656 24915 10659
rect 24946 10656 24952 10668
rect 24903 10628 24952 10656
rect 24903 10625 24915 10628
rect 24857 10619 24915 10625
rect 24946 10616 24952 10628
rect 25004 10616 25010 10668
rect 27890 10656 27896 10668
rect 27851 10628 27896 10656
rect 27890 10616 27896 10628
rect 27948 10616 27954 10668
rect 28077 10659 28135 10665
rect 28077 10625 28089 10659
rect 28123 10625 28135 10659
rect 28077 10619 28135 10625
rect 13127 10560 13216 10588
rect 13127 10557 13139 10560
rect 13081 10551 13139 10557
rect 13262 10548 13268 10600
rect 13320 10588 13326 10600
rect 15746 10588 15752 10600
rect 13320 10560 13365 10588
rect 15707 10560 15752 10588
rect 13320 10548 13326 10560
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 15930 10588 15936 10600
rect 15891 10560 15936 10588
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 16482 10548 16488 10600
rect 16540 10588 16546 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16540 10560 16957 10588
rect 16540 10548 16546 10560
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 16945 10551 17003 10557
rect 17126 10548 17132 10600
rect 17184 10588 17190 10600
rect 17402 10588 17408 10600
rect 17184 10560 17408 10588
rect 17184 10548 17190 10560
rect 17402 10548 17408 10560
rect 17460 10548 17466 10600
rect 18138 10588 18144 10600
rect 18099 10560 18144 10588
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 27614 10588 27620 10600
rect 19168 10560 27620 10588
rect 12400 10492 12848 10520
rect 13188 10492 16804 10520
rect 12400 10480 12406 10492
rect 9490 10452 9496 10464
rect 9232 10424 9496 10452
rect 9490 10412 9496 10424
rect 9548 10452 9554 10464
rect 10962 10452 10968 10464
rect 9548 10424 10968 10452
rect 9548 10412 9554 10424
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 12802 10412 12808 10464
rect 12860 10452 12866 10464
rect 13188 10452 13216 10492
rect 12860 10424 13216 10452
rect 12860 10412 12866 10424
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13780 10424 13829 10452
rect 13780 10412 13786 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 16666 10452 16672 10464
rect 16627 10424 16672 10452
rect 13817 10415 13875 10421
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 16776 10452 16804 10492
rect 19168 10452 19196 10560
rect 27614 10548 27620 10560
rect 27672 10588 27678 10600
rect 28092 10588 28120 10619
rect 29914 10616 29920 10668
rect 29972 10656 29978 10668
rect 30742 10656 30748 10668
rect 29972 10628 30748 10656
rect 29972 10616 29978 10628
rect 30742 10616 30748 10628
rect 30800 10656 30806 10668
rect 31205 10659 31263 10665
rect 31205 10656 31217 10659
rect 30800 10628 31217 10656
rect 30800 10616 30806 10628
rect 31205 10625 31217 10628
rect 31251 10625 31263 10659
rect 38470 10656 38476 10668
rect 38431 10628 38476 10656
rect 31205 10619 31263 10625
rect 38470 10616 38476 10628
rect 38528 10656 38534 10668
rect 38948 10656 38976 10696
rect 39114 10656 39120 10668
rect 38528 10628 38976 10656
rect 39075 10628 39120 10656
rect 38528 10616 38534 10628
rect 39114 10616 39120 10628
rect 39172 10616 39178 10668
rect 39574 10616 39580 10668
rect 39632 10656 39638 10668
rect 40221 10659 40279 10665
rect 40221 10656 40233 10659
rect 39632 10628 40233 10656
rect 39632 10616 39638 10628
rect 40221 10625 40233 10628
rect 40267 10625 40279 10659
rect 40328 10656 40356 10696
rect 40681 10659 40739 10665
rect 40681 10656 40693 10659
rect 40328 10628 40693 10656
rect 40221 10619 40279 10625
rect 40681 10625 40693 10628
rect 40727 10625 40739 10659
rect 40681 10619 40739 10625
rect 47578 10616 47584 10668
rect 47636 10656 47642 10668
rect 48205 10659 48263 10665
rect 48205 10656 48217 10659
rect 47636 10628 48217 10656
rect 47636 10616 47642 10628
rect 48205 10625 48217 10628
rect 48251 10625 48263 10659
rect 48205 10619 48263 10625
rect 27672 10560 28120 10588
rect 31113 10591 31171 10597
rect 27672 10548 27678 10560
rect 31113 10557 31125 10591
rect 31159 10557 31171 10591
rect 31113 10551 31171 10557
rect 24946 10480 24952 10532
rect 25004 10520 25010 10532
rect 25590 10520 25596 10532
rect 25004 10492 25596 10520
rect 25004 10480 25010 10492
rect 25590 10480 25596 10492
rect 25648 10480 25654 10532
rect 31128 10520 31156 10551
rect 47118 10548 47124 10600
rect 47176 10588 47182 10600
rect 47949 10591 48007 10597
rect 47949 10588 47961 10591
rect 47176 10560 47961 10588
rect 47176 10548 47182 10560
rect 47949 10557 47961 10560
rect 47995 10557 48007 10591
rect 47949 10551 48007 10557
rect 31202 10520 31208 10532
rect 31128 10492 31208 10520
rect 31202 10480 31208 10492
rect 31260 10480 31266 10532
rect 40770 10520 40776 10532
rect 39408 10492 40776 10520
rect 16776 10424 19196 10452
rect 21726 10412 21732 10464
rect 21784 10452 21790 10464
rect 22465 10455 22523 10461
rect 22465 10452 22477 10455
rect 21784 10424 22477 10452
rect 21784 10412 21790 10424
rect 22465 10421 22477 10424
rect 22511 10421 22523 10455
rect 27982 10452 27988 10464
rect 27943 10424 27988 10452
rect 22465 10415 22523 10421
rect 27982 10412 27988 10424
rect 28040 10412 28046 10464
rect 31478 10452 31484 10464
rect 31439 10424 31484 10452
rect 31478 10412 31484 10424
rect 31536 10412 31542 10464
rect 38562 10412 38568 10464
rect 38620 10452 38626 10464
rect 38838 10452 38844 10464
rect 38620 10424 38844 10452
rect 38620 10412 38626 10424
rect 38838 10412 38844 10424
rect 38896 10452 38902 10464
rect 39408 10461 39436 10492
rect 40770 10480 40776 10492
rect 40828 10480 40834 10532
rect 39393 10455 39451 10461
rect 39393 10452 39405 10455
rect 38896 10424 39405 10452
rect 38896 10412 38902 10424
rect 39393 10421 39405 10424
rect 39439 10421 39451 10455
rect 39574 10452 39580 10464
rect 39535 10424 39580 10452
rect 39393 10415 39451 10421
rect 39574 10412 39580 10424
rect 39632 10412 39638 10464
rect 40586 10452 40592 10464
rect 40547 10424 40592 10452
rect 40586 10412 40592 10424
rect 40644 10412 40650 10464
rect 40681 10455 40739 10461
rect 40681 10421 40693 10455
rect 40727 10452 40739 10455
rect 41322 10452 41328 10464
rect 40727 10424 41328 10452
rect 40727 10421 40739 10424
rect 40681 10415 40739 10421
rect 41322 10412 41328 10424
rect 41380 10412 41386 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 2130 10248 2136 10260
rect 2091 10220 2136 10248
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 3418 10248 3424 10260
rect 2516 10220 3424 10248
rect 2516 10053 2544 10220
rect 3418 10208 3424 10220
rect 3476 10248 3482 10260
rect 6273 10251 6331 10257
rect 6273 10248 6285 10251
rect 3476 10220 6285 10248
rect 3476 10208 3482 10220
rect 6273 10217 6285 10220
rect 6319 10217 6331 10251
rect 6273 10211 6331 10217
rect 6457 10251 6515 10257
rect 6457 10217 6469 10251
rect 6503 10248 6515 10251
rect 7282 10248 7288 10260
rect 6503 10220 7288 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 6288 10180 6316 10211
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 7745 10251 7803 10257
rect 7745 10217 7757 10251
rect 7791 10248 7803 10251
rect 10042 10248 10048 10260
rect 7791 10220 10048 10248
rect 7791 10217 7803 10220
rect 7745 10211 7803 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10226 10248 10232 10260
rect 10183 10220 10232 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 13262 10248 13268 10260
rect 11572 10220 13268 10248
rect 11572 10208 11578 10220
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 16853 10251 16911 10257
rect 16853 10248 16865 10251
rect 15804 10220 16865 10248
rect 15804 10208 15810 10220
rect 16853 10217 16865 10220
rect 16899 10217 16911 10251
rect 38010 10248 38016 10260
rect 16853 10211 16911 10217
rect 22066 10220 38016 10248
rect 7377 10183 7435 10189
rect 6288 10152 7052 10180
rect 2682 10112 2688 10124
rect 2643 10084 2688 10112
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 6362 10112 6368 10124
rect 6227 10084 6368 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 6362 10072 6368 10084
rect 6420 10112 6426 10124
rect 6822 10112 6828 10124
rect 6420 10084 6828 10112
rect 6420 10072 6426 10084
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10013 2559 10047
rect 2501 10007 2559 10013
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 3326 10044 3332 10056
rect 2639 10016 3332 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 5994 10044 6000 10056
rect 5955 10016 6000 10044
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10044 6331 10047
rect 6730 10044 6736 10056
rect 6319 10016 6736 10044
rect 6319 10013 6331 10016
rect 6273 10007 6331 10013
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10013 6975 10047
rect 7024 10044 7052 10152
rect 7377 10149 7389 10183
rect 7423 10180 7435 10183
rect 8478 10180 8484 10192
rect 7423 10152 8484 10180
rect 7423 10149 7435 10152
rect 7377 10143 7435 10149
rect 8478 10140 8484 10152
rect 8536 10140 8542 10192
rect 22066 10180 22094 10220
rect 38010 10208 38016 10220
rect 38068 10248 38074 10260
rect 38470 10248 38476 10260
rect 38068 10220 38476 10248
rect 38068 10208 38074 10220
rect 38470 10208 38476 10220
rect 38528 10208 38534 10260
rect 39114 10248 39120 10260
rect 39075 10220 39120 10248
rect 39114 10208 39120 10220
rect 39172 10208 39178 10260
rect 40770 10208 40776 10260
rect 40828 10248 40834 10260
rect 42613 10251 42671 10257
rect 42613 10248 42625 10251
rect 40828 10220 42625 10248
rect 40828 10208 40834 10220
rect 42613 10217 42625 10220
rect 42659 10217 42671 10251
rect 47578 10248 47584 10260
rect 47539 10220 47584 10248
rect 42613 10211 42671 10217
rect 47578 10208 47584 10220
rect 47636 10208 47642 10260
rect 47854 10208 47860 10260
rect 47912 10248 47918 10260
rect 47949 10251 48007 10257
rect 47949 10248 47961 10251
rect 47912 10220 47961 10248
rect 47912 10208 47918 10220
rect 47949 10217 47961 10220
rect 47995 10217 48007 10251
rect 47949 10211 48007 10217
rect 51442 10208 51448 10260
rect 51500 10248 51506 10260
rect 52917 10251 52975 10257
rect 52917 10248 52929 10251
rect 51500 10220 52929 10248
rect 51500 10208 51506 10220
rect 52917 10217 52929 10220
rect 52963 10217 52975 10251
rect 52917 10211 52975 10217
rect 9876 10152 22094 10180
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7469 10115 7527 10121
rect 7469 10112 7481 10115
rect 7248 10084 7481 10112
rect 7248 10072 7254 10084
rect 7469 10081 7481 10084
rect 7515 10081 7527 10115
rect 7469 10075 7527 10081
rect 7650 10044 7656 10056
rect 7024 10016 7656 10044
rect 6917 10007 6975 10013
rect 6932 9976 6960 10007
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 9876 10053 9904 10152
rect 22462 10140 22468 10192
rect 22520 10180 22526 10192
rect 22649 10183 22707 10189
rect 22649 10180 22661 10183
rect 22520 10152 22661 10180
rect 22520 10140 22526 10152
rect 22649 10149 22661 10152
rect 22695 10149 22707 10183
rect 22649 10143 22707 10149
rect 42242 10140 42248 10192
rect 42300 10180 42306 10192
rect 48682 10180 48688 10192
rect 42300 10152 48688 10180
rect 42300 10140 42306 10152
rect 48682 10140 48688 10152
rect 48740 10140 48746 10192
rect 13722 10112 13728 10124
rect 12268 10084 13728 10112
rect 12268 10053 12296 10084
rect 13722 10072 13728 10084
rect 13780 10072 13786 10124
rect 16850 10072 16856 10124
rect 16908 10112 16914 10124
rect 17037 10115 17095 10121
rect 17037 10112 17049 10115
rect 16908 10084 17049 10112
rect 16908 10072 16914 10084
rect 17037 10081 17049 10084
rect 17083 10081 17095 10115
rect 17037 10075 17095 10081
rect 17313 10115 17371 10121
rect 17313 10081 17325 10115
rect 17359 10112 17371 10115
rect 18046 10112 18052 10124
rect 17359 10084 18052 10112
rect 17359 10081 17371 10084
rect 17313 10075 17371 10081
rect 18046 10072 18052 10084
rect 18104 10072 18110 10124
rect 26326 10112 26332 10124
rect 25056 10084 26332 10112
rect 25056 10056 25084 10084
rect 26326 10072 26332 10084
rect 26384 10072 26390 10124
rect 27430 10112 27436 10124
rect 27391 10084 27436 10112
rect 27430 10072 27436 10084
rect 27488 10072 27494 10124
rect 30653 10115 30711 10121
rect 30653 10081 30665 10115
rect 30699 10112 30711 10115
rect 31662 10112 31668 10124
rect 30699 10084 31668 10112
rect 30699 10081 30711 10084
rect 30653 10075 30711 10081
rect 31662 10072 31668 10084
rect 31720 10072 31726 10124
rect 42426 10072 42432 10124
rect 42484 10112 42490 10124
rect 46293 10115 46351 10121
rect 46293 10112 46305 10115
rect 42484 10084 46305 10112
rect 42484 10072 42490 10084
rect 46293 10081 46305 10084
rect 46339 10081 46351 10115
rect 48038 10112 48044 10124
rect 47999 10084 48044 10112
rect 46293 10075 46351 10081
rect 48038 10072 48044 10084
rect 48096 10072 48102 10124
rect 51074 10072 51080 10124
rect 51132 10112 51138 10124
rect 51534 10112 51540 10124
rect 51132 10084 51540 10112
rect 51132 10072 51138 10084
rect 51534 10072 51540 10084
rect 51592 10072 51598 10124
rect 9861 10047 9919 10053
rect 9861 10044 9873 10047
rect 9824 10016 9873 10044
rect 9824 10004 9830 10016
rect 9861 10013 9873 10016
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12529 10047 12587 10053
rect 12529 10044 12541 10047
rect 12253 10007 12311 10013
rect 12406 10016 12541 10044
rect 7466 9976 7472 9988
rect 6932 9948 7472 9976
rect 7466 9936 7472 9948
rect 7524 9936 7530 9988
rect 8478 9936 8484 9988
rect 8536 9976 8542 9988
rect 12406 9976 12434 10016
rect 12529 10013 12541 10016
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10044 13139 10047
rect 13354 10044 13360 10056
rect 13127 10016 13360 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10044 13507 10047
rect 14090 10044 14096 10056
rect 13495 10016 14096 10044
rect 13495 10013 13507 10016
rect 13449 10007 13507 10013
rect 13464 9976 13492 10007
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 15657 10047 15715 10053
rect 15657 10013 15669 10047
rect 15703 10044 15715 10047
rect 15838 10044 15844 10056
rect 15703 10016 15844 10044
rect 15703 10013 15715 10016
rect 15657 10007 15715 10013
rect 15838 10004 15844 10016
rect 15896 10044 15902 10056
rect 16482 10044 16488 10056
rect 15896 10016 16488 10044
rect 15896 10004 15902 10016
rect 16482 10004 16488 10016
rect 16540 10044 16546 10056
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16540 10016 17141 10044
rect 16540 10004 16546 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 17221 10047 17279 10053
rect 17221 10013 17233 10047
rect 17267 10044 17279 10047
rect 20070 10044 20076 10056
rect 17267 10016 20076 10044
rect 17267 10013 17279 10016
rect 17221 10007 17279 10013
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 21910 10004 21916 10056
rect 21968 10044 21974 10056
rect 22005 10047 22063 10053
rect 22005 10044 22017 10047
rect 21968 10016 22017 10044
rect 21968 10004 21974 10016
rect 22005 10013 22017 10016
rect 22051 10013 22063 10047
rect 22005 10007 22063 10013
rect 22098 10047 22156 10053
rect 22098 10013 22110 10047
rect 22144 10013 22156 10047
rect 22098 10007 22156 10013
rect 8536 9948 12434 9976
rect 13188 9948 13492 9976
rect 13541 9979 13599 9985
rect 8536 9936 8542 9948
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 12158 9908 12164 9920
rect 11112 9880 12164 9908
rect 11112 9868 11118 9880
rect 12158 9868 12164 9880
rect 12216 9908 12222 9920
rect 13188 9908 13216 9948
rect 13541 9945 13553 9979
rect 13587 9976 13599 9979
rect 13587 9948 16436 9976
rect 13587 9945 13599 9948
rect 13541 9939 13599 9945
rect 12216 9880 13216 9908
rect 12216 9868 12222 9880
rect 13446 9868 13452 9920
rect 13504 9908 13510 9920
rect 13556 9908 13584 9939
rect 13504 9880 13584 9908
rect 15749 9911 15807 9917
rect 13504 9868 13510 9880
rect 15749 9877 15761 9911
rect 15795 9908 15807 9911
rect 16298 9908 16304 9920
rect 15795 9880 16304 9908
rect 15795 9877 15807 9880
rect 15749 9871 15807 9877
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 16408 9908 16436 9948
rect 21726 9936 21732 9988
rect 21784 9976 21790 9988
rect 22112 9976 22140 10007
rect 22462 10004 22468 10056
rect 22520 10053 22526 10056
rect 22520 10044 22528 10053
rect 22520 10016 22565 10044
rect 22520 10007 22528 10016
rect 22520 10004 22526 10007
rect 24578 10004 24584 10056
rect 24636 10044 24642 10056
rect 24946 10053 24952 10056
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 24636 10016 24777 10044
rect 24636 10004 24642 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 24913 10047 24952 10053
rect 24913 10013 24925 10047
rect 24913 10007 24952 10013
rect 24946 10004 24952 10007
rect 25004 10004 25010 10056
rect 25038 10004 25044 10056
rect 25096 10044 25102 10056
rect 25096 10016 25189 10044
rect 25096 10004 25102 10016
rect 25222 10004 25228 10056
rect 25280 10053 25286 10056
rect 25280 10044 25288 10053
rect 30926 10044 30932 10056
rect 25280 10016 25325 10044
rect 30887 10016 30932 10044
rect 25280 10007 25288 10016
rect 25280 10004 25286 10007
rect 30926 10004 30932 10016
rect 30984 10004 30990 10056
rect 36173 10047 36231 10053
rect 36173 10013 36185 10047
rect 36219 10013 36231 10047
rect 36173 10007 36231 10013
rect 36357 10047 36415 10053
rect 36357 10013 36369 10047
rect 36403 10044 36415 10047
rect 36446 10044 36452 10056
rect 36403 10016 36452 10044
rect 36403 10013 36415 10016
rect 36357 10007 36415 10013
rect 21784 9948 22140 9976
rect 22281 9979 22339 9985
rect 21784 9936 21790 9948
rect 22281 9945 22293 9979
rect 22327 9945 22339 9979
rect 22281 9939 22339 9945
rect 22373 9979 22431 9985
rect 22373 9945 22385 9979
rect 22419 9976 22431 9979
rect 23658 9976 23664 9988
rect 22419 9948 23664 9976
rect 22419 9945 22431 9948
rect 22373 9939 22431 9945
rect 22296 9908 22324 9939
rect 23658 9936 23664 9948
rect 23716 9936 23722 9988
rect 25133 9979 25191 9985
rect 25133 9945 25145 9979
rect 25179 9976 25191 9979
rect 27700 9979 27758 9985
rect 25179 9948 27660 9976
rect 25179 9945 25191 9948
rect 25133 9939 25191 9945
rect 22738 9908 22744 9920
rect 16408 9880 22744 9908
rect 22738 9868 22744 9880
rect 22796 9868 22802 9920
rect 23382 9868 23388 9920
rect 23440 9908 23446 9920
rect 25409 9911 25467 9917
rect 25409 9908 25421 9911
rect 23440 9880 25421 9908
rect 23440 9868 23446 9880
rect 25409 9877 25421 9880
rect 25455 9877 25467 9911
rect 27632 9908 27660 9948
rect 27700 9945 27712 9979
rect 27746 9976 27758 9979
rect 28074 9976 28080 9988
rect 27746 9948 28080 9976
rect 27746 9945 27758 9948
rect 27700 9939 27758 9945
rect 28074 9936 28080 9948
rect 28132 9936 28138 9988
rect 36188 9976 36216 10007
rect 36446 10004 36452 10016
rect 36504 10044 36510 10056
rect 37001 10047 37059 10053
rect 37001 10044 37013 10047
rect 36504 10016 37013 10044
rect 36504 10004 36510 10016
rect 37001 10013 37013 10016
rect 37047 10013 37059 10047
rect 37642 10044 37648 10056
rect 37603 10016 37648 10044
rect 37001 10007 37059 10013
rect 37642 10004 37648 10016
rect 37700 10004 37706 10056
rect 37829 10047 37887 10053
rect 37829 10013 37841 10047
rect 37875 10013 37887 10047
rect 38838 10044 38844 10056
rect 38799 10016 38844 10044
rect 37829 10007 37887 10013
rect 36538 9976 36544 9988
rect 36188 9948 36544 9976
rect 36538 9936 36544 9948
rect 36596 9976 36602 9988
rect 36817 9979 36875 9985
rect 36817 9976 36829 9979
rect 36596 9948 36829 9976
rect 36596 9936 36602 9948
rect 36817 9945 36829 9948
rect 36863 9945 36875 9979
rect 37182 9976 37188 9988
rect 37143 9948 37188 9976
rect 36817 9939 36875 9945
rect 37182 9936 37188 9948
rect 37240 9936 37246 9988
rect 37274 9936 37280 9988
rect 37332 9976 37338 9988
rect 37844 9976 37872 10007
rect 38838 10004 38844 10016
rect 38896 10004 38902 10056
rect 41230 10044 41236 10056
rect 41191 10016 41236 10044
rect 41230 10004 41236 10016
rect 41288 10004 41294 10056
rect 41322 10004 41328 10056
rect 41380 10044 41386 10056
rect 41489 10047 41547 10053
rect 41489 10044 41501 10047
rect 41380 10016 41501 10044
rect 41380 10004 41386 10016
rect 41489 10013 41501 10016
rect 41535 10013 41547 10047
rect 41489 10007 41547 10013
rect 46109 10047 46167 10053
rect 46109 10013 46121 10047
rect 46155 10013 46167 10047
rect 46109 10007 46167 10013
rect 46385 10047 46443 10053
rect 46385 10013 46397 10047
rect 46431 10044 46443 10047
rect 46566 10044 46572 10056
rect 46431 10016 46572 10044
rect 46431 10013 46443 10016
rect 46385 10007 46443 10013
rect 37332 9948 37872 9976
rect 37332 9936 37338 9948
rect 37918 9936 37924 9988
rect 37976 9976 37982 9988
rect 44634 9976 44640 9988
rect 37976 9948 44640 9976
rect 37976 9936 37982 9948
rect 44634 9936 44640 9948
rect 44692 9936 44698 9988
rect 46124 9976 46152 10007
rect 46566 10004 46572 10016
rect 46624 10004 46630 10056
rect 47765 10047 47823 10053
rect 47765 10013 47777 10047
rect 47811 10013 47823 10047
rect 47765 10007 47823 10013
rect 46474 9976 46480 9988
rect 46124 9948 46480 9976
rect 46474 9936 46480 9948
rect 46532 9976 46538 9988
rect 47780 9976 47808 10007
rect 51626 10004 51632 10056
rect 51684 10044 51690 10056
rect 51793 10047 51851 10053
rect 51793 10044 51805 10047
rect 51684 10016 51805 10044
rect 51684 10004 51690 10016
rect 51793 10013 51805 10016
rect 51839 10013 51851 10047
rect 51793 10007 51851 10013
rect 48774 9976 48780 9988
rect 46532 9948 48780 9976
rect 46532 9936 46538 9948
rect 48774 9936 48780 9948
rect 48832 9936 48838 9988
rect 28166 9908 28172 9920
rect 27632 9880 28172 9908
rect 25409 9871 25467 9877
rect 28166 9868 28172 9880
rect 28224 9868 28230 9920
rect 28810 9908 28816 9920
rect 28771 9880 28816 9908
rect 28810 9868 28816 9880
rect 28868 9868 28874 9920
rect 30742 9868 30748 9920
rect 30800 9908 30806 9920
rect 32033 9911 32091 9917
rect 32033 9908 32045 9911
rect 30800 9880 32045 9908
rect 30800 9868 30806 9880
rect 32033 9877 32045 9880
rect 32079 9877 32091 9911
rect 32033 9871 32091 9877
rect 36265 9911 36323 9917
rect 36265 9877 36277 9911
rect 36311 9908 36323 9911
rect 36446 9908 36452 9920
rect 36311 9880 36452 9908
rect 36311 9877 36323 9880
rect 36265 9871 36323 9877
rect 36446 9868 36452 9880
rect 36504 9868 36510 9920
rect 37458 9868 37464 9920
rect 37516 9908 37522 9920
rect 37737 9911 37795 9917
rect 37737 9908 37749 9911
rect 37516 9880 37749 9908
rect 37516 9868 37522 9880
rect 37737 9877 37749 9880
rect 37783 9877 37795 9911
rect 37737 9871 37795 9877
rect 38930 9868 38936 9920
rect 38988 9908 38994 9920
rect 39301 9911 39359 9917
rect 39301 9908 39313 9911
rect 38988 9880 39313 9908
rect 38988 9868 38994 9880
rect 39301 9877 39313 9880
rect 39347 9877 39359 9911
rect 45922 9908 45928 9920
rect 45883 9880 45928 9908
rect 39301 9871 39359 9877
rect 45922 9868 45928 9880
rect 45980 9868 45986 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 2593 9707 2651 9713
rect 2593 9704 2605 9707
rect 1452 9676 2605 9704
rect 1452 9664 1458 9676
rect 2593 9673 2605 9676
rect 2639 9673 2651 9707
rect 2593 9667 2651 9673
rect 5074 9664 5080 9716
rect 5132 9704 5138 9716
rect 15473 9707 15531 9713
rect 15473 9704 15485 9707
rect 5132 9676 15485 9704
rect 5132 9664 5138 9676
rect 15473 9673 15485 9676
rect 15519 9673 15531 9707
rect 16666 9704 16672 9716
rect 15473 9667 15531 9673
rect 15672 9676 16672 9704
rect 2501 9639 2559 9645
rect 2501 9605 2513 9639
rect 2547 9636 2559 9639
rect 3326 9636 3332 9648
rect 2547 9608 3332 9636
rect 2547 9605 2559 9608
rect 2501 9599 2559 9605
rect 3326 9596 3332 9608
rect 3384 9596 3390 9648
rect 10045 9639 10103 9645
rect 10045 9605 10057 9639
rect 10091 9636 10103 9639
rect 10594 9636 10600 9648
rect 10091 9608 10600 9636
rect 10091 9605 10103 9608
rect 10045 9599 10103 9605
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 12526 9596 12532 9648
rect 12584 9636 12590 9648
rect 12584 9608 14872 9636
rect 12584 9596 12590 9608
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 1412 9432 1440 9531
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 8297 9571 8355 9577
rect 8297 9568 8309 9571
rect 8260 9540 8309 9568
rect 8260 9528 8266 9540
rect 8297 9537 8309 9540
rect 8343 9537 8355 9571
rect 8297 9531 8355 9537
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 9950 9568 9956 9580
rect 9907 9540 9956 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 13265 9571 13323 9577
rect 12492 9540 12537 9568
rect 12492 9528 12498 9540
rect 13265 9537 13277 9571
rect 13311 9568 13323 9571
rect 13354 9568 13360 9580
rect 13311 9540 13360 9568
rect 13311 9537 13323 9540
rect 13265 9531 13323 9537
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 14844 9577 14872 9608
rect 14918 9596 14924 9648
rect 14976 9636 14982 9648
rect 15013 9639 15071 9645
rect 15013 9636 15025 9639
rect 14976 9608 15025 9636
rect 14976 9596 14982 9608
rect 15013 9605 15025 9608
rect 15059 9605 15071 9639
rect 15013 9599 15071 9605
rect 15672 9577 15700 9676
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 21744 9676 22232 9704
rect 17218 9636 17224 9648
rect 15764 9608 17224 9636
rect 15764 9577 15792 9608
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 21744 9636 21772 9676
rect 17328 9608 21772 9636
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9568 14887 9571
rect 15657 9571 15715 9577
rect 14875 9540 15516 9568
rect 14875 9537 14887 9540
rect 14829 9531 14887 9537
rect 2682 9500 2688 9512
rect 2643 9472 2688 9500
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 4890 9460 4896 9512
rect 4948 9500 4954 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 4948 9472 6929 9500
rect 4948 9460 4954 9472
rect 6917 9469 6929 9472
rect 6963 9500 6975 9503
rect 7190 9500 7196 9512
rect 6963 9472 7196 9500
rect 6963 9469 6975 9472
rect 6917 9463 6975 9469
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7466 9500 7472 9512
rect 7427 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9500 7895 9503
rect 11054 9500 11060 9512
rect 7883 9472 11060 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 13170 9500 13176 9512
rect 13131 9472 13176 9500
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 5994 9432 6000 9444
rect 1412 9404 6000 9432
rect 5994 9392 6000 9404
rect 6052 9392 6058 9444
rect 7282 9432 7288 9444
rect 7243 9404 7288 9432
rect 7282 9392 7288 9404
rect 7340 9392 7346 9444
rect 7377 9435 7435 9441
rect 7377 9401 7389 9435
rect 7423 9432 7435 9435
rect 8294 9432 8300 9444
rect 7423 9404 8300 9432
rect 7423 9401 7435 9404
rect 7377 9395 7435 9401
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 8478 9432 8484 9444
rect 8439 9404 8484 9432
rect 8478 9392 8484 9404
rect 8536 9392 8542 9444
rect 14090 9392 14096 9444
rect 14148 9432 14154 9444
rect 14918 9432 14924 9444
rect 14148 9404 14924 9432
rect 14148 9392 14154 9404
rect 14918 9392 14924 9404
rect 14976 9392 14982 9444
rect 15488 9432 15516 9540
rect 15657 9537 15669 9571
rect 15703 9537 15715 9571
rect 15657 9531 15715 9537
rect 15749 9571 15807 9577
rect 15749 9537 15761 9571
rect 15795 9537 15807 9571
rect 15749 9531 15807 9537
rect 15838 9500 15844 9512
rect 15799 9472 15844 9500
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 15930 9460 15936 9512
rect 15988 9500 15994 9512
rect 15988 9472 16033 9500
rect 15988 9460 15994 9472
rect 15488 9404 15700 9432
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 2133 9367 2191 9373
rect 2133 9333 2145 9367
rect 2179 9364 2191 9367
rect 2406 9364 2412 9376
rect 2179 9336 2412 9364
rect 2179 9333 2191 9336
rect 2133 9327 2191 9333
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 9858 9324 9864 9376
rect 9916 9364 9922 9376
rect 10229 9367 10287 9373
rect 10229 9364 10241 9367
rect 9916 9336 10241 9364
rect 9916 9324 9922 9336
rect 10229 9333 10241 9336
rect 10275 9333 10287 9367
rect 10229 9327 10287 9333
rect 13541 9367 13599 9373
rect 13541 9333 13553 9367
rect 13587 9364 13599 9367
rect 15562 9364 15568 9376
rect 13587 9336 15568 9364
rect 13587 9333 13599 9336
rect 13541 9327 13599 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 15672 9364 15700 9404
rect 17328 9364 17356 9608
rect 21818 9596 21824 9648
rect 21876 9636 21882 9648
rect 22066 9639 22124 9645
rect 22066 9636 22078 9639
rect 21876 9608 22078 9636
rect 21876 9596 21882 9608
rect 22066 9605 22078 9608
rect 22112 9605 22124 9639
rect 22204 9636 22232 9676
rect 22278 9664 22284 9716
rect 22336 9704 22342 9716
rect 23106 9704 23112 9716
rect 22336 9676 23112 9704
rect 22336 9664 22342 9676
rect 23106 9664 23112 9676
rect 23164 9664 23170 9716
rect 28074 9704 28080 9716
rect 28035 9676 28080 9704
rect 28074 9664 28080 9676
rect 28132 9664 28138 9716
rect 30926 9704 30932 9716
rect 23198 9636 23204 9648
rect 22204 9608 23204 9636
rect 22066 9599 22124 9605
rect 23198 9596 23204 9608
rect 23256 9636 23262 9648
rect 23382 9636 23388 9648
rect 23256 9608 23388 9636
rect 23256 9596 23262 9608
rect 23382 9596 23388 9608
rect 23440 9596 23446 9648
rect 28629 9639 28687 9645
rect 28629 9636 28641 9639
rect 25608 9608 28641 9636
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 18325 9571 18383 9577
rect 18325 9568 18337 9571
rect 18196 9540 18337 9568
rect 18196 9528 18202 9540
rect 18325 9537 18337 9540
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 18592 9571 18650 9577
rect 18592 9537 18604 9571
rect 18638 9568 18650 9571
rect 19150 9568 19156 9580
rect 18638 9540 19156 9568
rect 18638 9537 18650 9540
rect 18592 9531 18650 9537
rect 19150 9528 19156 9540
rect 19208 9528 19214 9580
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 25608 9568 25636 9608
rect 28629 9605 28641 9608
rect 28675 9636 28687 9639
rect 28810 9636 28816 9686
rect 28675 9634 28816 9636
rect 28868 9634 28874 9686
rect 28902 9634 28908 9686
rect 28960 9636 28966 9686
rect 30887 9676 30932 9704
rect 30926 9664 30932 9676
rect 30984 9664 30990 9716
rect 31202 9664 31208 9716
rect 31260 9704 31266 9716
rect 42242 9704 42248 9716
rect 31260 9676 42248 9704
rect 31260 9664 31266 9676
rect 42242 9664 42248 9676
rect 42300 9664 42306 9716
rect 42426 9704 42432 9716
rect 42387 9676 42432 9704
rect 42426 9664 42432 9676
rect 42484 9664 42490 9716
rect 31478 9636 31484 9648
rect 28960 9634 31340 9636
rect 28675 9608 28856 9634
rect 28920 9608 31340 9634
rect 31439 9608 31484 9636
rect 28675 9605 28687 9608
rect 28629 9599 28687 9605
rect 19392 9540 25636 9568
rect 25961 9571 26019 9577
rect 19392 9528 19398 9540
rect 25961 9537 25973 9571
rect 26007 9537 26019 9571
rect 25961 9531 26019 9537
rect 21821 9503 21879 9509
rect 21821 9469 21833 9503
rect 21867 9469 21879 9503
rect 24670 9500 24676 9512
rect 24631 9472 24676 9500
rect 21821 9463 21879 9469
rect 19426 9392 19432 9444
rect 19484 9432 19490 9444
rect 19705 9435 19763 9441
rect 19705 9432 19717 9435
rect 19484 9404 19717 9432
rect 19484 9392 19490 9404
rect 19705 9401 19717 9404
rect 19751 9401 19763 9435
rect 19705 9395 19763 9401
rect 15672 9336 17356 9364
rect 18138 9324 18144 9376
rect 18196 9364 18202 9376
rect 21836 9364 21864 9463
rect 24670 9460 24676 9472
rect 24728 9460 24734 9512
rect 24949 9503 25007 9509
rect 24949 9469 24961 9503
rect 24995 9500 25007 9503
rect 25222 9500 25228 9512
rect 24995 9472 25228 9500
rect 24995 9469 25007 9472
rect 24949 9463 25007 9469
rect 24964 9432 24992 9463
rect 25222 9460 25228 9472
rect 25280 9460 25286 9512
rect 25682 9460 25688 9512
rect 25740 9500 25746 9512
rect 25976 9500 26004 9531
rect 27982 9528 27988 9580
rect 28040 9568 28046 9580
rect 28353 9571 28411 9577
rect 28353 9568 28365 9571
rect 28040 9540 28365 9568
rect 28040 9528 28046 9540
rect 28353 9537 28365 9540
rect 28399 9568 28411 9571
rect 31205 9571 31263 9577
rect 28920 9568 29040 9569
rect 31205 9568 31217 9571
rect 28399 9541 31217 9568
rect 28399 9540 28948 9541
rect 29012 9540 31217 9541
rect 28399 9537 28411 9540
rect 28353 9531 28411 9537
rect 31205 9537 31217 9540
rect 31251 9537 31263 9571
rect 31205 9531 31263 9537
rect 25740 9472 26004 9500
rect 28261 9503 28319 9509
rect 25740 9460 25746 9472
rect 28261 9469 28273 9503
rect 28307 9469 28319 9503
rect 28261 9463 28319 9469
rect 28276 9432 28304 9463
rect 28626 9460 28632 9512
rect 28684 9500 28690 9512
rect 28721 9503 28779 9509
rect 28721 9500 28733 9503
rect 28684 9472 28733 9500
rect 28684 9460 28690 9472
rect 28721 9469 28733 9472
rect 28767 9500 28779 9503
rect 28902 9500 28908 9512
rect 28767 9472 28908 9500
rect 28767 9469 28779 9472
rect 28721 9463 28779 9469
rect 28902 9460 28908 9472
rect 28960 9460 28966 9512
rect 31114 9503 31172 9509
rect 31114 9469 31126 9503
rect 31160 9469 31172 9503
rect 31312 9500 31340 9608
rect 31478 9596 31484 9608
rect 31536 9596 31542 9648
rect 31588 9608 32904 9636
rect 31588 9509 31616 9608
rect 32876 9568 32904 9608
rect 33134 9596 33140 9648
rect 33192 9636 33198 9648
rect 33318 9636 33324 9648
rect 33192 9608 33324 9636
rect 33192 9596 33198 9608
rect 33318 9596 33324 9608
rect 33376 9596 33382 9648
rect 34054 9636 34060 9648
rect 33428 9608 34060 9636
rect 33428 9568 33456 9608
rect 34054 9596 34060 9608
rect 34112 9596 34118 9648
rect 35713 9639 35771 9645
rect 35713 9605 35725 9639
rect 35759 9636 35771 9639
rect 36814 9636 36820 9648
rect 35759 9608 36820 9636
rect 35759 9605 35771 9608
rect 35713 9599 35771 9605
rect 36814 9596 36820 9608
rect 36872 9596 36878 9648
rect 37642 9596 37648 9648
rect 37700 9636 37706 9648
rect 39025 9639 39083 9645
rect 39025 9636 39037 9639
rect 37700 9608 39037 9636
rect 37700 9596 37706 9608
rect 39025 9605 39037 9608
rect 39071 9605 39083 9639
rect 39025 9599 39083 9605
rect 42794 9596 42800 9648
rect 42852 9636 42858 9648
rect 45922 9645 45928 9648
rect 45916 9636 45928 9645
rect 42852 9608 42897 9636
rect 45883 9608 45928 9636
rect 42852 9596 42858 9608
rect 45916 9599 45928 9608
rect 45922 9596 45928 9599
rect 45980 9596 45986 9648
rect 49237 9639 49295 9645
rect 49237 9605 49249 9639
rect 49283 9605 49295 9639
rect 49237 9599 49295 9605
rect 49453 9639 49511 9645
rect 49453 9605 49465 9639
rect 49499 9636 49511 9639
rect 49694 9636 49700 9648
rect 49499 9608 49700 9636
rect 49499 9605 49511 9608
rect 49453 9599 49511 9605
rect 33594 9577 33600 9580
rect 32876 9540 33456 9568
rect 33577 9571 33600 9577
rect 33577 9537 33589 9571
rect 33577 9531 33600 9537
rect 33594 9528 33600 9531
rect 33652 9528 33658 9580
rect 36538 9528 36544 9580
rect 36596 9568 36602 9580
rect 37274 9568 37280 9580
rect 36596 9540 36641 9568
rect 37235 9540 37280 9568
rect 36596 9528 36602 9540
rect 37274 9528 37280 9540
rect 37332 9528 37338 9580
rect 38930 9568 38936 9580
rect 38891 9540 38936 9568
rect 38930 9528 38936 9540
rect 38988 9528 38994 9580
rect 39117 9571 39175 9577
rect 39117 9537 39129 9571
rect 39163 9568 39175 9571
rect 39574 9568 39580 9580
rect 39163 9540 39580 9568
rect 39163 9537 39175 9540
rect 39117 9531 39175 9537
rect 39574 9528 39580 9540
rect 39632 9528 39638 9580
rect 39758 9568 39764 9580
rect 39719 9540 39764 9568
rect 39758 9528 39764 9540
rect 39816 9528 39822 9580
rect 42610 9568 42616 9580
rect 42571 9540 42616 9568
rect 42610 9528 42616 9540
rect 42668 9528 42674 9580
rect 42702 9528 42708 9580
rect 42760 9568 42766 9580
rect 42760 9540 42805 9568
rect 42760 9528 42766 9540
rect 42886 9528 42892 9580
rect 42944 9577 42950 9580
rect 42944 9571 42973 9577
rect 42961 9537 42973 9571
rect 47118 9568 47124 9580
rect 42944 9531 42973 9537
rect 45664 9540 47124 9568
rect 42944 9528 42950 9531
rect 31573 9503 31631 9509
rect 31573 9500 31585 9503
rect 31312 9472 31585 9500
rect 31114 9463 31172 9469
rect 31573 9469 31585 9472
rect 31619 9469 31631 9503
rect 31573 9463 31631 9469
rect 31128 9432 31156 9463
rect 31846 9460 31852 9512
rect 31904 9500 31910 9512
rect 32674 9500 32680 9512
rect 31904 9472 32680 9500
rect 31904 9460 31910 9472
rect 32674 9460 32680 9472
rect 32732 9500 32738 9512
rect 33321 9503 33379 9509
rect 33321 9500 33333 9503
rect 32732 9472 33333 9500
rect 32732 9460 32738 9472
rect 33321 9469 33333 9472
rect 33367 9469 33379 9503
rect 33321 9463 33379 9469
rect 36357 9503 36415 9509
rect 36357 9469 36369 9503
rect 36403 9500 36415 9503
rect 37292 9500 37320 9528
rect 42794 9500 42800 9512
rect 36403 9472 37320 9500
rect 37660 9472 42800 9500
rect 36403 9469 36415 9472
rect 36357 9463 36415 9469
rect 33134 9432 33140 9444
rect 23124 9404 24992 9432
rect 25332 9404 26280 9432
rect 28276 9404 33140 9432
rect 18196 9336 21864 9364
rect 18196 9324 18202 9336
rect 22462 9324 22468 9376
rect 22520 9364 22526 9376
rect 23124 9364 23152 9404
rect 22520 9336 23152 9364
rect 22520 9324 22526 9336
rect 23198 9324 23204 9376
rect 23256 9364 23262 9376
rect 23256 9336 23301 9364
rect 23256 9324 23262 9336
rect 23382 9324 23388 9376
rect 23440 9364 23446 9376
rect 25332 9364 25360 9404
rect 26142 9364 26148 9376
rect 23440 9336 25360 9364
rect 26103 9336 26148 9364
rect 23440 9324 23446 9336
rect 26142 9324 26148 9336
rect 26200 9324 26206 9376
rect 26252 9364 26280 9404
rect 33134 9392 33140 9404
rect 33192 9392 33198 9444
rect 37660 9432 37688 9472
rect 42794 9460 42800 9472
rect 42852 9460 42858 9512
rect 45664 9509 45692 9540
rect 47118 9528 47124 9540
rect 47176 9528 47182 9580
rect 43073 9503 43131 9509
rect 43073 9469 43085 9503
rect 43119 9469 43131 9503
rect 43073 9463 43131 9469
rect 45649 9503 45707 9509
rect 45649 9469 45661 9503
rect 45695 9469 45707 9503
rect 49252 9500 49280 9599
rect 49694 9596 49700 9608
rect 49752 9596 49758 9648
rect 49510 9500 49516 9512
rect 49252 9472 49516 9500
rect 45649 9463 45707 9469
rect 39758 9432 39764 9444
rect 34624 9404 37688 9432
rect 37752 9404 39764 9432
rect 30190 9364 30196 9376
rect 26252 9336 30196 9364
rect 30190 9324 30196 9336
rect 30248 9324 30254 9376
rect 30834 9324 30840 9376
rect 30892 9364 30898 9376
rect 34624 9364 34652 9404
rect 30892 9336 34652 9364
rect 34701 9367 34759 9373
rect 30892 9324 30898 9336
rect 34701 9333 34713 9367
rect 34747 9364 34759 9367
rect 35342 9364 35348 9376
rect 34747 9336 35348 9364
rect 34747 9333 34759 9336
rect 34701 9327 34759 9333
rect 35342 9324 35348 9336
rect 35400 9324 35406 9376
rect 35802 9364 35808 9376
rect 35763 9336 35808 9364
rect 35802 9324 35808 9336
rect 35860 9364 35866 9376
rect 36170 9364 36176 9376
rect 35860 9336 36176 9364
rect 35860 9324 35866 9336
rect 36170 9324 36176 9336
rect 36228 9324 36234 9376
rect 36722 9364 36728 9376
rect 36683 9336 36728 9364
rect 36722 9324 36728 9336
rect 36780 9324 36786 9376
rect 36814 9324 36820 9376
rect 36872 9364 36878 9376
rect 37507 9367 37565 9373
rect 37507 9364 37519 9367
rect 36872 9336 37519 9364
rect 36872 9324 36878 9336
rect 37507 9333 37519 9336
rect 37553 9364 37565 9367
rect 37752 9364 37780 9404
rect 39758 9392 39764 9404
rect 39816 9392 39822 9444
rect 39850 9392 39856 9444
rect 39908 9432 39914 9444
rect 43088 9432 43116 9463
rect 49510 9460 49516 9472
rect 49568 9460 49574 9512
rect 39908 9404 43116 9432
rect 39908 9392 39914 9404
rect 43162 9392 43168 9444
rect 43220 9432 43226 9444
rect 45370 9432 45376 9444
rect 43220 9404 45376 9432
rect 43220 9392 43226 9404
rect 45370 9392 45376 9404
rect 45428 9392 45434 9444
rect 46952 9404 49464 9432
rect 37553 9336 37780 9364
rect 37553 9333 37565 9336
rect 37507 9327 37565 9333
rect 38470 9324 38476 9376
rect 38528 9364 38534 9376
rect 39577 9367 39635 9373
rect 39577 9364 39589 9367
rect 38528 9336 39589 9364
rect 38528 9324 38534 9336
rect 39577 9333 39589 9336
rect 39623 9333 39635 9367
rect 39577 9327 39635 9333
rect 41690 9324 41696 9376
rect 41748 9364 41754 9376
rect 46290 9364 46296 9376
rect 41748 9336 46296 9364
rect 41748 9324 41754 9336
rect 46290 9324 46296 9336
rect 46348 9364 46354 9376
rect 46952 9364 46980 9404
rect 49436 9376 49464 9404
rect 46348 9336 46980 9364
rect 46348 9324 46354 9336
rect 47026 9324 47032 9376
rect 47084 9364 47090 9376
rect 48498 9364 48504 9376
rect 47084 9336 48504 9364
rect 47084 9324 47090 9336
rect 48498 9324 48504 9336
rect 48556 9324 48562 9376
rect 49418 9364 49424 9376
rect 49331 9336 49424 9364
rect 49418 9324 49424 9336
rect 49476 9324 49482 9376
rect 49602 9364 49608 9376
rect 49563 9336 49608 9364
rect 49602 9324 49608 9336
rect 49660 9324 49666 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 5902 9160 5908 9172
rect 5863 9132 5908 9160
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 8202 9160 8208 9172
rect 8163 9132 8208 9160
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 9309 9163 9367 9169
rect 9309 9129 9321 9163
rect 9355 9160 9367 9163
rect 9398 9160 9404 9172
rect 9355 9132 9404 9160
rect 9355 9129 9367 9132
rect 9309 9123 9367 9129
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 10042 9160 10048 9172
rect 10003 9132 10048 9160
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 10318 9160 10324 9172
rect 10279 9132 10324 9160
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 13538 9160 13544 9172
rect 13499 9132 13544 9160
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 14304 9163 14362 9169
rect 14304 9160 14316 9163
rect 13780 9132 14316 9160
rect 13780 9120 13786 9132
rect 14304 9129 14316 9132
rect 14350 9129 14362 9163
rect 14304 9123 14362 9129
rect 19150 9120 19156 9172
rect 19208 9160 19214 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 19208 9132 19257 9160
rect 19208 9120 19214 9132
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 19245 9123 19303 9129
rect 19352 9132 22094 9160
rect 13078 9092 13084 9104
rect 12912 9064 13084 9092
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 4525 9027 4583 9033
rect 4525 9024 4537 9027
rect 1912 8996 4537 9024
rect 1912 8984 1918 8996
rect 4525 8993 4537 8996
rect 4571 8993 4583 9027
rect 4525 8987 4583 8993
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 2406 8956 2412 8968
rect 2367 8928 2412 8956
rect 2406 8916 2412 8928
rect 2464 8916 2470 8968
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 4540 8956 4568 8987
rect 4614 8956 4620 8968
rect 4540 8928 4620 8956
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 8846 8956 8852 8968
rect 8435 8928 8852 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 4792 8891 4850 8897
rect 4792 8857 4804 8891
rect 4838 8888 4850 8891
rect 5166 8888 5172 8900
rect 4838 8860 5172 8888
rect 4838 8857 4850 8860
rect 4792 8851 4850 8857
rect 5166 8848 5172 8860
rect 5224 8848 5230 8900
rect 8220 8888 8248 8919
rect 8846 8916 8852 8928
rect 8904 8956 8910 8968
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 8904 8928 9137 8956
rect 8904 8916 8910 8928
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9858 8956 9864 8968
rect 9819 8928 9864 8956
rect 9125 8919 9183 8925
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 12912 8965 12940 9064
rect 13078 9052 13084 9064
rect 13136 9052 13142 9104
rect 13446 9092 13452 9104
rect 13188 9064 13452 9092
rect 13078 8965 13084 8968
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8925 12955 8959
rect 12897 8919 12955 8925
rect 13045 8959 13084 8965
rect 13045 8925 13057 8959
rect 13045 8919 13084 8925
rect 13078 8916 13084 8919
rect 13136 8916 13142 8968
rect 13188 8965 13216 9064
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 19352 9092 19380 9132
rect 20162 9092 20168 9104
rect 14384 9064 19380 9092
rect 19444 9064 20168 9092
rect 13262 8984 13268 9036
rect 13320 8984 13326 9036
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8925 13231 8959
rect 13280 8956 13308 8984
rect 13403 8959 13461 8965
rect 13403 8956 13415 8959
rect 13280 8928 13415 8956
rect 13173 8919 13231 8925
rect 13403 8925 13415 8928
rect 13449 8956 13461 8959
rect 13538 8956 13544 8968
rect 13449 8928 13544 8956
rect 13449 8925 13461 8928
rect 13403 8919 13461 8925
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 8941 8891 8999 8897
rect 8941 8888 8953 8891
rect 8220 8860 8953 8888
rect 8941 8857 8953 8860
rect 8987 8888 8999 8891
rect 10042 8888 10048 8900
rect 8987 8860 10048 8888
rect 8987 8857 8999 8860
rect 8941 8851 8999 8857
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 14090 8888 14096 8900
rect 13320 8860 13365 8888
rect 14051 8860 14096 8888
rect 13320 8848 13326 8860
rect 14090 8848 14096 8860
rect 14148 8848 14154 8900
rect 1397 8823 1455 8829
rect 1397 8789 1409 8823
rect 1443 8820 1455 8823
rect 2038 8820 2044 8832
rect 1443 8792 2044 8820
rect 1443 8789 1455 8792
rect 1397 8783 1455 8789
rect 2038 8780 2044 8792
rect 2096 8780 2102 8832
rect 2222 8820 2228 8832
rect 2183 8792 2228 8820
rect 2222 8780 2228 8792
rect 2280 8780 2286 8832
rect 2869 8823 2927 8829
rect 2869 8789 2881 8823
rect 2915 8820 2927 8823
rect 5810 8820 5816 8832
rect 2915 8792 5816 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 5810 8780 5816 8792
rect 5868 8780 5874 8832
rect 14277 8823 14335 8829
rect 14277 8789 14289 8823
rect 14323 8820 14335 8823
rect 14384 8820 14412 9064
rect 15189 9027 15247 9033
rect 15189 8993 15201 9027
rect 15235 9024 15247 9027
rect 16025 9027 16083 9033
rect 16025 9024 16037 9027
rect 15235 8996 16037 9024
rect 15235 8993 15247 8996
rect 15189 8987 15247 8993
rect 16025 8993 16037 8996
rect 16071 8993 16083 9027
rect 16025 8987 16083 8993
rect 16393 9027 16451 9033
rect 16393 8993 16405 9027
rect 16439 9024 16451 9027
rect 19334 9024 19340 9036
rect 16439 8996 19340 9024
rect 16439 8993 16451 8996
rect 16393 8987 16451 8993
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 15382 8959 15440 8965
rect 15382 8925 15394 8959
rect 15428 8925 15440 8959
rect 15382 8919 15440 8925
rect 15473 8959 15531 8965
rect 15473 8925 15485 8959
rect 15519 8956 15531 8959
rect 15746 8956 15752 8968
rect 15519 8928 15752 8956
rect 15519 8925 15531 8928
rect 15473 8919 15531 8925
rect 14323 8792 14412 8820
rect 14461 8823 14519 8829
rect 14323 8789 14335 8792
rect 14277 8783 14335 8789
rect 14461 8789 14473 8823
rect 14507 8820 14519 8823
rect 14826 8820 14832 8832
rect 14507 8792 14832 8820
rect 14507 8789 14519 8792
rect 14461 8783 14519 8789
rect 14826 8780 14832 8792
rect 14884 8780 14890 8832
rect 15010 8820 15016 8832
rect 14971 8792 15016 8820
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 15304 8820 15332 8919
rect 15397 8888 15425 8919
rect 15746 8916 15752 8928
rect 15804 8956 15810 8968
rect 15930 8956 15936 8968
rect 15804 8928 15936 8956
rect 15804 8916 15810 8928
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 16209 8959 16267 8965
rect 16209 8925 16221 8959
rect 16255 8925 16267 8959
rect 16209 8919 16267 8925
rect 15838 8888 15844 8900
rect 15397 8860 15844 8888
rect 15838 8848 15844 8860
rect 15896 8848 15902 8900
rect 16224 8888 16252 8919
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 16485 8959 16543 8965
rect 16356 8928 16401 8956
rect 16356 8916 16362 8928
rect 16485 8925 16497 8959
rect 16531 8956 16543 8959
rect 17402 8956 17408 8968
rect 16531 8928 17408 8956
rect 16531 8925 16543 8928
rect 16485 8919 16543 8925
rect 17402 8916 17408 8928
rect 17460 8916 17466 8968
rect 19444 8965 19472 9064
rect 20162 9052 20168 9064
rect 20220 9052 20226 9104
rect 21726 9052 21732 9104
rect 21784 9092 21790 9104
rect 21913 9095 21971 9101
rect 21913 9092 21925 9095
rect 21784 9064 21925 9092
rect 21784 9052 21790 9064
rect 21913 9061 21925 9064
rect 21959 9061 21971 9095
rect 22066 9092 22094 9132
rect 22554 9120 22560 9172
rect 22612 9160 22618 9172
rect 23198 9160 23204 9172
rect 22612 9132 23204 9160
rect 22612 9120 22618 9132
rect 23198 9120 23204 9132
rect 23256 9120 23262 9172
rect 25130 9120 25136 9172
rect 25188 9160 25194 9172
rect 25409 9163 25467 9169
rect 25409 9160 25421 9163
rect 25188 9132 25421 9160
rect 25188 9120 25194 9132
rect 25409 9129 25421 9132
rect 25455 9129 25467 9163
rect 25409 9123 25467 9129
rect 33321 9163 33379 9169
rect 33321 9129 33333 9163
rect 33367 9160 33379 9163
rect 33594 9160 33600 9172
rect 33367 9132 33600 9160
rect 33367 9129 33379 9132
rect 33321 9123 33379 9129
rect 33594 9120 33600 9132
rect 33652 9120 33658 9172
rect 33870 9120 33876 9172
rect 33928 9160 33934 9172
rect 37366 9160 37372 9172
rect 33928 9132 37372 9160
rect 33928 9120 33934 9132
rect 37366 9120 37372 9132
rect 37424 9120 37430 9172
rect 37550 9120 37556 9172
rect 37608 9160 37614 9172
rect 39850 9160 39856 9172
rect 37608 9132 39856 9160
rect 37608 9120 37614 9132
rect 39850 9120 39856 9132
rect 39908 9120 39914 9172
rect 41782 9120 41788 9172
rect 41840 9160 41846 9172
rect 42153 9163 42211 9169
rect 42153 9160 42165 9163
rect 41840 9132 42165 9160
rect 41840 9120 41846 9132
rect 42153 9129 42165 9132
rect 42199 9129 42211 9163
rect 42153 9123 42211 9129
rect 42242 9120 42248 9172
rect 42300 9160 42306 9172
rect 46198 9160 46204 9172
rect 42300 9132 46204 9160
rect 42300 9120 42306 9132
rect 46198 9120 46204 9132
rect 46256 9120 46262 9172
rect 46290 9120 46296 9172
rect 46348 9160 46354 9172
rect 50985 9163 51043 9169
rect 50985 9160 50997 9163
rect 46348 9132 46393 9160
rect 46492 9132 50997 9160
rect 46348 9120 46354 9132
rect 23014 9092 23020 9104
rect 22066 9064 23020 9092
rect 21913 9055 21971 9061
rect 23014 9052 23020 9064
rect 23072 9052 23078 9104
rect 24762 9052 24768 9104
rect 24820 9092 24826 9104
rect 24820 9064 28764 9092
rect 24820 9052 24826 9064
rect 24670 9024 24676 9036
rect 21836 8996 24676 9024
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8956 19763 8959
rect 19978 8956 19984 8968
rect 19751 8928 19984 8956
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 19978 8916 19984 8928
rect 20036 8916 20042 8968
rect 16850 8888 16856 8900
rect 16224 8860 16856 8888
rect 16850 8848 16856 8860
rect 16908 8848 16914 8900
rect 17034 8848 17040 8900
rect 17092 8888 17098 8900
rect 21836 8888 21864 8996
rect 24670 8984 24676 8996
rect 24728 8984 24734 9036
rect 28736 9024 28764 9064
rect 28902 9052 28908 9104
rect 28960 9092 28966 9104
rect 44542 9092 44548 9104
rect 28960 9064 44548 9092
rect 28960 9052 28966 9064
rect 44542 9052 44548 9064
rect 44600 9052 44606 9104
rect 44726 9052 44732 9104
rect 44784 9092 44790 9104
rect 46492 9092 46520 9132
rect 50985 9129 50997 9132
rect 51031 9129 51043 9163
rect 50985 9123 51043 9129
rect 44784 9064 46520 9092
rect 44784 9052 44790 9064
rect 33594 9024 33600 9036
rect 28736 8996 33600 9024
rect 33594 8984 33600 8996
rect 33652 8984 33658 9036
rect 36725 9027 36783 9033
rect 36725 9024 36737 9027
rect 36464 8996 36737 9024
rect 22097 8959 22155 8965
rect 22097 8925 22109 8959
rect 22143 8956 22155 8959
rect 22554 8956 22560 8968
rect 22143 8928 22560 8956
rect 22143 8925 22155 8928
rect 22097 8919 22155 8925
rect 22554 8916 22560 8928
rect 22612 8916 22618 8968
rect 22646 8916 22652 8968
rect 22704 8956 22710 8968
rect 22833 8959 22891 8965
rect 22833 8956 22845 8959
rect 22704 8928 22845 8956
rect 22704 8916 22710 8928
rect 22833 8925 22845 8928
rect 22879 8925 22891 8959
rect 22833 8919 22891 8925
rect 23109 8959 23167 8965
rect 23109 8925 23121 8959
rect 23155 8956 23167 8959
rect 24578 8956 24584 8968
rect 23155 8928 24584 8956
rect 23155 8925 23167 8928
rect 23109 8919 23167 8925
rect 17092 8860 21864 8888
rect 17092 8848 17098 8860
rect 21910 8848 21916 8900
rect 21968 8888 21974 8900
rect 23124 8888 23152 8919
rect 24578 8916 24584 8928
rect 24636 8956 24642 8968
rect 24765 8959 24823 8965
rect 24765 8956 24777 8959
rect 24636 8928 24777 8956
rect 24636 8916 24642 8928
rect 24765 8925 24777 8928
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 24858 8959 24916 8965
rect 24858 8925 24870 8959
rect 24904 8925 24916 8959
rect 25038 8956 25044 8968
rect 24999 8928 25044 8956
rect 24858 8919 24916 8925
rect 21968 8860 23152 8888
rect 21968 8848 21974 8860
rect 23198 8848 23204 8900
rect 23256 8888 23262 8900
rect 24873 8888 24901 8919
rect 25038 8916 25044 8928
rect 25096 8916 25102 8968
rect 25222 8916 25228 8968
rect 25280 8965 25286 8968
rect 25280 8956 25288 8965
rect 25280 8928 25325 8956
rect 25280 8919 25288 8928
rect 25280 8916 25286 8919
rect 27798 8916 27804 8968
rect 27856 8956 27862 8968
rect 27985 8959 28043 8965
rect 27985 8956 27997 8959
rect 27856 8928 27997 8956
rect 27856 8916 27862 8928
rect 27985 8925 27997 8928
rect 28031 8925 28043 8959
rect 27985 8919 28043 8925
rect 28629 8959 28687 8965
rect 28629 8925 28641 8959
rect 28675 8956 28687 8959
rect 28810 8956 28816 8968
rect 28675 8928 28816 8956
rect 28675 8925 28687 8928
rect 28629 8919 28687 8925
rect 28810 8916 28816 8928
rect 28868 8916 28874 8968
rect 28902 8916 28908 8968
rect 28960 8916 28966 8968
rect 33502 8956 33508 8968
rect 33463 8928 33508 8956
rect 33502 8916 33508 8928
rect 33560 8916 33566 8968
rect 33870 8965 33876 8968
rect 33827 8959 33876 8965
rect 33827 8925 33839 8959
rect 33873 8925 33876 8959
rect 33827 8919 33876 8925
rect 33870 8916 33876 8919
rect 33928 8916 33934 8968
rect 33965 8959 34023 8965
rect 33965 8925 33977 8959
rect 34011 8956 34023 8959
rect 34054 8956 34060 8968
rect 34011 8928 34060 8956
rect 34011 8925 34023 8928
rect 33965 8919 34023 8925
rect 34054 8916 34060 8928
rect 34112 8916 34118 8968
rect 34238 8916 34244 8968
rect 34296 8956 34302 8968
rect 36262 8956 36268 8968
rect 34296 8928 36268 8956
rect 34296 8916 34302 8928
rect 36262 8916 36268 8928
rect 36320 8916 36326 8968
rect 36464 8956 36492 8996
rect 36725 8993 36737 8996
rect 36771 8993 36783 9027
rect 36725 8987 36783 8993
rect 36817 9027 36875 9033
rect 36817 8993 36829 9027
rect 36863 9024 36875 9027
rect 37458 9024 37464 9036
rect 36863 8996 37320 9024
rect 37419 8996 37464 9024
rect 36863 8993 36875 8996
rect 36817 8987 36875 8993
rect 36630 8956 36636 8968
rect 36372 8928 36492 8956
rect 36591 8928 36636 8956
rect 23256 8860 24901 8888
rect 25133 8891 25191 8897
rect 23256 8848 23262 8860
rect 25133 8857 25145 8891
rect 25179 8888 25191 8891
rect 26050 8888 26056 8900
rect 25179 8860 26056 8888
rect 25179 8857 25191 8860
rect 25133 8851 25191 8857
rect 26050 8848 26056 8860
rect 26108 8848 26114 8900
rect 27706 8848 27712 8900
rect 27764 8888 27770 8900
rect 27764 8860 28488 8888
rect 27764 8848 27770 8860
rect 16574 8820 16580 8832
rect 15304 8792 16580 8820
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 19484 8792 19625 8820
rect 19484 8780 19490 8792
rect 19613 8789 19625 8792
rect 19659 8789 19671 8823
rect 19613 8783 19671 8789
rect 22094 8780 22100 8832
rect 22152 8820 22158 8832
rect 22738 8820 22744 8832
rect 22152 8792 22744 8820
rect 22152 8780 22158 8792
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 27801 8823 27859 8829
rect 27801 8789 27813 8823
rect 27847 8820 27859 8823
rect 27890 8820 27896 8832
rect 27847 8792 27896 8820
rect 27847 8789 27859 8792
rect 27801 8783 27859 8789
rect 27890 8780 27896 8792
rect 27948 8780 27954 8832
rect 28460 8829 28488 8860
rect 28534 8848 28540 8900
rect 28592 8888 28598 8900
rect 28920 8888 28948 8916
rect 28592 8860 28948 8888
rect 33597 8891 33655 8897
rect 28592 8848 28598 8860
rect 33597 8857 33609 8891
rect 33643 8857 33655 8891
rect 33597 8851 33655 8857
rect 28445 8823 28503 8829
rect 28445 8789 28457 8823
rect 28491 8820 28503 8823
rect 28902 8820 28908 8832
rect 28491 8792 28908 8820
rect 28491 8789 28503 8792
rect 28445 8783 28503 8789
rect 28902 8780 28908 8792
rect 28960 8780 28966 8832
rect 33612 8820 33640 8851
rect 33686 8848 33692 8900
rect 33744 8888 33750 8900
rect 35526 8888 35532 8900
rect 33744 8860 35532 8888
rect 33744 8848 33750 8860
rect 35526 8848 35532 8860
rect 35584 8848 35590 8900
rect 36372 8832 36400 8928
rect 36630 8916 36636 8928
rect 36688 8916 36694 8968
rect 36909 8959 36967 8965
rect 36909 8925 36921 8959
rect 36955 8956 36967 8959
rect 37182 8956 37188 8968
rect 36955 8928 37188 8956
rect 36955 8925 36967 8928
rect 36909 8919 36967 8925
rect 37182 8916 37188 8928
rect 37240 8916 37246 8968
rect 37292 8956 37320 8996
rect 37458 8984 37464 8996
rect 37516 9024 37522 9036
rect 37516 8996 38884 9024
rect 37516 8984 37522 8996
rect 37642 8956 37648 8968
rect 37292 8928 37648 8956
rect 37642 8916 37648 8928
rect 37700 8916 37706 8968
rect 37734 8916 37740 8968
rect 37792 8956 37798 8968
rect 38856 8965 38884 8996
rect 41506 8984 41512 9036
rect 41564 9024 41570 9036
rect 41564 8996 42564 9024
rect 41564 8984 41570 8996
rect 38841 8959 38899 8965
rect 37792 8928 37837 8956
rect 37792 8916 37798 8928
rect 38841 8925 38853 8959
rect 38887 8925 38899 8959
rect 38841 8919 38899 8925
rect 39025 8959 39083 8965
rect 39025 8925 39037 8959
rect 39071 8956 39083 8959
rect 39114 8956 39120 8968
rect 39071 8928 39120 8956
rect 39071 8925 39083 8928
rect 39025 8919 39083 8925
rect 39114 8916 39120 8928
rect 39172 8916 39178 8968
rect 42426 8956 42432 8968
rect 41984 8928 42432 8956
rect 36998 8848 37004 8900
rect 37056 8888 37062 8900
rect 41874 8888 41880 8900
rect 37056 8860 41880 8888
rect 37056 8848 37062 8860
rect 41874 8848 41880 8860
rect 41932 8848 41938 8900
rect 41984 8897 42012 8928
rect 42426 8916 42432 8928
rect 42484 8916 42490 8968
rect 42536 8956 42564 8996
rect 45002 8984 45008 9036
rect 45060 9024 45066 9036
rect 45060 8996 45324 9024
rect 45060 8984 45066 8996
rect 43162 8956 43168 8968
rect 42536 8928 43168 8956
rect 43162 8916 43168 8928
rect 43220 8916 43226 8968
rect 44910 8916 44916 8968
rect 44968 8956 44974 8968
rect 45296 8965 45324 8996
rect 45370 8984 45376 9036
rect 45428 9024 45434 9036
rect 46658 9024 46664 9036
rect 45428 8996 46664 9024
rect 45428 8984 45434 8996
rect 46658 8984 46664 8996
rect 46716 8984 46722 9036
rect 51534 9024 51540 9036
rect 51495 8996 51540 9024
rect 51534 8984 51540 8996
rect 51592 8984 51598 9036
rect 45189 8959 45247 8965
rect 45189 8956 45201 8959
rect 44968 8928 45201 8956
rect 44968 8916 44974 8928
rect 45189 8925 45201 8928
rect 45235 8925 45247 8959
rect 45189 8919 45247 8925
rect 45281 8959 45339 8965
rect 45281 8925 45293 8959
rect 45327 8925 45339 8959
rect 45281 8919 45339 8925
rect 45649 8959 45707 8965
rect 45649 8925 45661 8959
rect 45695 8956 45707 8959
rect 47026 8956 47032 8968
rect 45695 8928 47032 8956
rect 45695 8925 45707 8928
rect 45649 8919 45707 8925
rect 42242 8897 42248 8900
rect 41969 8891 42027 8897
rect 41969 8857 41981 8891
rect 42015 8857 42027 8891
rect 42185 8891 42248 8897
rect 42185 8888 42197 8891
rect 41969 8851 42027 8857
rect 42076 8860 42197 8888
rect 34790 8820 34796 8832
rect 33612 8792 34796 8820
rect 34790 8780 34796 8792
rect 34848 8780 34854 8832
rect 36354 8780 36360 8832
rect 36412 8780 36418 8832
rect 36449 8823 36507 8829
rect 36449 8789 36461 8823
rect 36495 8820 36507 8823
rect 36906 8820 36912 8832
rect 36495 8792 36912 8820
rect 36495 8789 36507 8792
rect 36449 8783 36507 8789
rect 36906 8780 36912 8792
rect 36964 8780 36970 8832
rect 38746 8780 38752 8832
rect 38804 8820 38810 8832
rect 42076 8820 42104 8860
rect 42185 8857 42197 8860
rect 42231 8857 42248 8891
rect 42185 8851 42248 8857
rect 42242 8848 42248 8851
rect 42300 8848 42306 8900
rect 44174 8848 44180 8900
rect 44232 8888 44238 8900
rect 45373 8891 45431 8897
rect 45373 8888 45385 8891
rect 44232 8860 45385 8888
rect 44232 8848 44238 8860
rect 45373 8857 45385 8860
rect 45419 8857 45431 8891
rect 45373 8851 45431 8857
rect 45462 8848 45468 8900
rect 45520 8897 45526 8900
rect 46124 8897 46152 8928
rect 47026 8916 47032 8928
rect 47084 8916 47090 8968
rect 47118 8916 47124 8968
rect 47176 8956 47182 8968
rect 48225 8959 48283 8965
rect 48225 8956 48237 8959
rect 47176 8928 48237 8956
rect 47176 8916 47182 8928
rect 48225 8925 48237 8928
rect 48271 8925 48283 8959
rect 49694 8956 49700 8968
rect 48225 8919 48283 8925
rect 48332 8928 49700 8956
rect 45520 8891 45549 8897
rect 45537 8857 45549 8891
rect 45520 8851 45549 8857
rect 46109 8891 46167 8897
rect 46109 8857 46121 8891
rect 46155 8857 46167 8891
rect 46290 8888 46296 8900
rect 46348 8897 46354 8900
rect 46348 8891 46383 8897
rect 46235 8860 46296 8888
rect 46109 8851 46167 8857
rect 45520 8848 45526 8851
rect 46290 8848 46296 8860
rect 46371 8888 46383 8891
rect 48332 8888 48360 8928
rect 49694 8916 49700 8928
rect 49752 8916 49758 8968
rect 50801 8959 50859 8965
rect 50801 8956 50813 8959
rect 50540 8928 50813 8956
rect 46371 8860 48360 8888
rect 48492 8891 48550 8897
rect 46371 8857 46383 8860
rect 46348 8851 46383 8857
rect 48492 8857 48504 8891
rect 48538 8888 48550 8891
rect 48590 8888 48596 8900
rect 48538 8860 48596 8888
rect 48538 8857 48550 8860
rect 48492 8851 48550 8857
rect 46348 8848 46354 8851
rect 48590 8848 48596 8860
rect 48648 8848 48654 8900
rect 50540 8888 50568 8928
rect 50801 8925 50813 8928
rect 50847 8925 50859 8959
rect 50801 8919 50859 8925
rect 51074 8916 51080 8968
rect 51132 8956 51138 8968
rect 51132 8928 51177 8956
rect 51132 8916 51138 8928
rect 48700 8860 50568 8888
rect 42334 8820 42340 8832
rect 38804 8792 42104 8820
rect 42295 8792 42340 8820
rect 38804 8780 38810 8792
rect 42334 8780 42340 8792
rect 42392 8780 42398 8832
rect 45005 8823 45063 8829
rect 45005 8789 45017 8823
rect 45051 8820 45063 8823
rect 46198 8820 46204 8832
rect 45051 8792 46204 8820
rect 45051 8789 45063 8792
rect 45005 8783 45063 8789
rect 46198 8780 46204 8792
rect 46256 8780 46262 8832
rect 46477 8823 46535 8829
rect 46477 8789 46489 8823
rect 46523 8820 46535 8823
rect 46566 8820 46572 8832
rect 46523 8792 46572 8820
rect 46523 8789 46535 8792
rect 46477 8783 46535 8789
rect 46566 8780 46572 8792
rect 46624 8780 46630 8832
rect 46658 8780 46664 8832
rect 46716 8820 46722 8832
rect 48700 8820 48728 8860
rect 46716 8792 48728 8820
rect 46716 8780 46722 8792
rect 49510 8780 49516 8832
rect 49568 8820 49574 8832
rect 49605 8823 49663 8829
rect 49605 8820 49617 8823
rect 49568 8792 49617 8820
rect 49568 8780 49574 8792
rect 49605 8789 49617 8792
rect 49651 8789 49663 8823
rect 50540 8820 50568 8860
rect 50617 8891 50675 8897
rect 50617 8857 50629 8891
rect 50663 8888 50675 8891
rect 51782 8891 51840 8897
rect 51782 8888 51794 8891
rect 50663 8860 51794 8888
rect 50663 8857 50675 8860
rect 50617 8851 50675 8857
rect 51782 8857 51794 8860
rect 51828 8857 51840 8891
rect 51782 8851 51840 8857
rect 52730 8820 52736 8832
rect 50540 8792 52736 8820
rect 49605 8783 49663 8789
rect 52730 8780 52736 8792
rect 52788 8780 52794 8832
rect 52914 8820 52920 8832
rect 52875 8792 52920 8820
rect 52914 8780 52920 8792
rect 52972 8780 52978 8832
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 5166 8616 5172 8628
rect 5127 8588 5172 8616
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 13722 8616 13728 8628
rect 5868 8588 13728 8616
rect 5868 8576 5874 8588
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 17034 8616 17040 8628
rect 13832 8588 17040 8616
rect 2222 8557 2228 8560
rect 2216 8548 2228 8557
rect 2183 8520 2228 8548
rect 2216 8511 2228 8520
rect 2222 8508 2228 8511
rect 2280 8508 2286 8560
rect 5537 8551 5595 8557
rect 5537 8517 5549 8551
rect 5583 8548 5595 8551
rect 5902 8548 5908 8560
rect 5583 8520 5908 8548
rect 5583 8517 5595 8520
rect 5537 8511 5595 8517
rect 5902 8508 5908 8520
rect 5960 8508 5966 8560
rect 13538 8508 13544 8560
rect 13596 8548 13602 8560
rect 13832 8548 13860 8588
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 17862 8576 17868 8628
rect 17920 8616 17926 8628
rect 19889 8619 19947 8625
rect 17920 8588 19840 8616
rect 17920 8576 17926 8588
rect 13596 8520 13860 8548
rect 13596 8508 13602 8520
rect 15562 8508 15568 8560
rect 15620 8548 15626 8560
rect 19812 8548 19840 8588
rect 19889 8585 19901 8619
rect 19935 8616 19947 8619
rect 20070 8616 20076 8628
rect 19935 8588 20076 8616
rect 19935 8585 19947 8588
rect 19889 8579 19947 8585
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 22465 8619 22523 8625
rect 22465 8616 22477 8619
rect 20180 8588 22477 8616
rect 20180 8548 20208 8588
rect 22465 8585 22477 8588
rect 22511 8585 22523 8619
rect 25038 8616 25044 8628
rect 22465 8579 22523 8585
rect 24964 8588 25044 8616
rect 15620 8520 19748 8548
rect 19812 8520 20208 8548
rect 15620 8508 15626 8520
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 1949 8483 2007 8489
rect 1949 8480 1961 8483
rect 1912 8452 1961 8480
rect 1912 8440 1918 8452
rect 1949 8449 1961 8452
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8480 5687 8483
rect 5718 8480 5724 8492
rect 5675 8452 5724 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 5368 8412 5396 8443
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 16850 8440 16856 8492
rect 16908 8480 16914 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16908 8452 16957 8480
rect 16908 8440 16914 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 18138 8440 18144 8492
rect 18196 8480 18202 8492
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18196 8452 18521 8480
rect 18196 8440 18202 8452
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18776 8483 18834 8489
rect 18776 8449 18788 8483
rect 18822 8480 18834 8483
rect 19242 8480 19248 8492
rect 18822 8452 19248 8480
rect 18822 8449 18834 8452
rect 18776 8443 18834 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 19720 8480 19748 8520
rect 21174 8508 21180 8560
rect 21232 8548 21238 8560
rect 22189 8551 22247 8557
rect 22189 8548 22201 8551
rect 21232 8520 22201 8548
rect 21232 8508 21238 8520
rect 22189 8517 22201 8520
rect 22235 8517 22247 8551
rect 22189 8511 22247 8517
rect 24394 8508 24400 8560
rect 24452 8548 24458 8560
rect 24964 8557 24992 8588
rect 25038 8576 25044 8588
rect 25096 8576 25102 8628
rect 25317 8619 25375 8625
rect 25317 8585 25329 8619
rect 25363 8616 25375 8619
rect 25958 8616 25964 8628
rect 25363 8588 25964 8616
rect 25363 8585 25375 8588
rect 25317 8579 25375 8585
rect 25958 8576 25964 8588
rect 26016 8576 26022 8628
rect 28626 8616 28632 8628
rect 27540 8588 28632 8616
rect 24949 8551 25007 8557
rect 24452 8520 24808 8548
rect 24452 8508 24458 8520
rect 24780 8492 24808 8520
rect 24949 8517 24961 8551
rect 24995 8517 25007 8551
rect 27540 8548 27568 8588
rect 28626 8576 28632 8588
rect 28684 8576 28690 8628
rect 30466 8576 30472 8628
rect 30524 8616 30530 8628
rect 30524 8588 33456 8616
rect 30524 8576 30530 8588
rect 24949 8511 25007 8517
rect 25056 8520 27568 8548
rect 27617 8551 27675 8557
rect 21266 8480 21272 8492
rect 19720 8452 21272 8480
rect 21266 8440 21272 8452
rect 21324 8440 21330 8492
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21784 8452 21833 8480
rect 21784 8440 21790 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21941 8483 21999 8489
rect 21941 8480 21953 8483
rect 21821 8443 21879 8449
rect 21929 8449 21953 8480
rect 21987 8449 21999 8483
rect 21929 8443 21999 8449
rect 15010 8412 15016 8424
rect 5368 8384 15016 8412
rect 15010 8372 15016 8384
rect 15068 8372 15074 8424
rect 15286 8412 15292 8424
rect 15247 8384 15292 8412
rect 15286 8372 15292 8384
rect 15344 8372 15350 8424
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8412 15623 8415
rect 15746 8412 15752 8424
rect 15611 8384 15752 8412
rect 15611 8381 15623 8384
rect 15565 8375 15623 8381
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 16666 8412 16672 8424
rect 16627 8384 16672 8412
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 3326 8344 3332 8356
rect 3239 8316 3332 8344
rect 3326 8304 3332 8316
rect 3384 8344 3390 8356
rect 6730 8344 6736 8356
rect 3384 8316 6736 8344
rect 3384 8304 3390 8316
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 15304 8344 15332 8372
rect 16942 8344 16948 8356
rect 15304 8316 16948 8344
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 21818 8304 21824 8356
rect 21876 8344 21882 8356
rect 21929 8344 21957 8443
rect 22094 8440 22100 8492
rect 22152 8480 22158 8492
rect 22327 8483 22385 8489
rect 22152 8452 22197 8480
rect 22152 8440 22158 8452
rect 22327 8449 22339 8483
rect 22373 8480 22385 8483
rect 22462 8480 22468 8492
rect 22373 8452 22468 8480
rect 22373 8449 22385 8452
rect 22327 8443 22385 8449
rect 22462 8440 22468 8452
rect 22520 8440 22526 8492
rect 24578 8440 24584 8492
rect 24636 8480 24642 8492
rect 24673 8483 24731 8489
rect 24673 8480 24685 8483
rect 24636 8452 24685 8480
rect 24636 8440 24642 8452
rect 24673 8449 24685 8452
rect 24719 8449 24731 8483
rect 24673 8443 24731 8449
rect 24762 8440 24768 8492
rect 24820 8480 24826 8492
rect 25056 8489 25084 8520
rect 27617 8517 27629 8551
rect 27663 8517 27675 8551
rect 27617 8511 27675 8517
rect 25222 8489 25228 8492
rect 25041 8483 25099 8489
rect 24820 8452 24865 8480
rect 24820 8440 24826 8452
rect 25041 8449 25053 8483
rect 25087 8449 25099 8483
rect 25041 8443 25099 8449
rect 25179 8483 25228 8489
rect 25179 8449 25191 8483
rect 25225 8449 25228 8483
rect 25179 8443 25228 8449
rect 25222 8440 25228 8443
rect 25280 8440 25286 8492
rect 27632 8412 27660 8511
rect 27706 8508 27712 8560
rect 27764 8548 27770 8560
rect 27801 8551 27859 8557
rect 27801 8548 27813 8551
rect 27764 8520 27813 8548
rect 27764 8508 27770 8520
rect 27801 8517 27813 8520
rect 27847 8517 27859 8551
rect 27801 8511 27859 8517
rect 28445 8551 28503 8557
rect 28445 8517 28457 8551
rect 28491 8548 28503 8551
rect 28718 8548 28724 8560
rect 28491 8520 28724 8548
rect 28491 8517 28503 8520
rect 28445 8511 28503 8517
rect 28718 8508 28724 8520
rect 28776 8508 28782 8560
rect 28810 8508 28816 8560
rect 28868 8548 28874 8560
rect 28921 8551 28979 8557
rect 28921 8548 28933 8551
rect 28868 8520 28933 8548
rect 28868 8508 28874 8520
rect 28921 8517 28933 8520
rect 28967 8517 28979 8551
rect 33318 8548 33324 8560
rect 28921 8511 28979 8517
rect 30024 8520 32260 8548
rect 33279 8520 33324 8548
rect 30024 8480 30052 8520
rect 30190 8480 30196 8492
rect 22480 8384 27660 8412
rect 27724 8452 30052 8480
rect 30151 8452 30196 8480
rect 22480 8356 22508 8384
rect 21876 8316 21957 8344
rect 21876 8304 21882 8316
rect 22462 8304 22468 8356
rect 22520 8304 22526 8356
rect 26142 8304 26148 8356
rect 26200 8344 26206 8356
rect 27724 8344 27752 8452
rect 30190 8440 30196 8452
rect 30248 8440 30254 8492
rect 30469 8483 30527 8489
rect 30469 8449 30481 8483
rect 30515 8480 30527 8483
rect 30926 8480 30932 8492
rect 30515 8452 30932 8480
rect 30515 8449 30527 8452
rect 30469 8443 30527 8449
rect 30926 8440 30932 8452
rect 30984 8480 30990 8492
rect 32125 8483 32183 8489
rect 32125 8480 32137 8483
rect 30984 8452 32137 8480
rect 30984 8440 30990 8452
rect 32125 8449 32137 8452
rect 32171 8449 32183 8483
rect 32125 8443 32183 8449
rect 32232 8412 32260 8520
rect 33318 8508 33324 8520
rect 33376 8508 33382 8560
rect 33428 8548 33456 8588
rect 33502 8576 33508 8628
rect 33560 8616 33566 8628
rect 33689 8619 33747 8625
rect 33689 8616 33701 8619
rect 33560 8588 33701 8616
rect 33560 8576 33566 8588
rect 33689 8585 33701 8588
rect 33735 8585 33747 8619
rect 33689 8579 33747 8585
rect 33870 8576 33876 8628
rect 33928 8616 33934 8628
rect 39574 8616 39580 8628
rect 33928 8588 39580 8616
rect 33928 8576 33934 8588
rect 39574 8576 39580 8588
rect 39632 8576 39638 8628
rect 39669 8619 39727 8625
rect 39669 8585 39681 8619
rect 39715 8616 39727 8619
rect 41598 8616 41604 8628
rect 39715 8588 41604 8616
rect 39715 8585 39727 8588
rect 39669 8579 39727 8585
rect 41598 8576 41604 8588
rect 41656 8616 41662 8628
rect 41782 8616 41788 8628
rect 41656 8588 41788 8616
rect 41656 8576 41662 8588
rect 41782 8576 41788 8588
rect 41840 8576 41846 8628
rect 41874 8576 41880 8628
rect 41932 8616 41938 8628
rect 45462 8616 45468 8628
rect 41932 8588 45140 8616
rect 41932 8576 41938 8588
rect 42797 8551 42855 8557
rect 42797 8548 42809 8551
rect 33428 8520 42809 8548
rect 42797 8517 42809 8520
rect 42843 8517 42855 8551
rect 42797 8511 42855 8517
rect 42886 8508 42892 8560
rect 42944 8557 42950 8560
rect 42944 8551 42973 8557
rect 42961 8517 42973 8551
rect 44726 8548 44732 8560
rect 44687 8520 44732 8548
rect 42944 8511 42973 8517
rect 42944 8508 42950 8511
rect 44726 8508 44732 8520
rect 44784 8508 44790 8560
rect 45002 8548 45008 8560
rect 44963 8520 45008 8548
rect 45002 8508 45008 8520
rect 45060 8508 45066 8560
rect 45112 8557 45140 8588
rect 45204 8588 45468 8616
rect 45204 8557 45232 8588
rect 45462 8576 45468 8588
rect 45520 8576 45526 8628
rect 48590 8616 48596 8628
rect 48551 8588 48596 8616
rect 48590 8576 48596 8588
rect 48648 8576 48654 8628
rect 49694 8576 49700 8628
rect 49752 8616 49758 8628
rect 50449 8619 50507 8625
rect 50449 8616 50461 8619
rect 49752 8588 50461 8616
rect 49752 8576 49758 8588
rect 50449 8585 50461 8588
rect 50495 8585 50507 8619
rect 50449 8579 50507 8585
rect 50617 8619 50675 8625
rect 50617 8585 50629 8619
rect 50663 8616 50675 8619
rect 51074 8616 51080 8628
rect 50663 8588 51080 8616
rect 50663 8585 50675 8588
rect 50617 8579 50675 8585
rect 51074 8576 51080 8588
rect 51132 8576 51138 8628
rect 45097 8551 45155 8557
rect 45097 8517 45109 8551
rect 45143 8517 45155 8551
rect 45204 8551 45273 8557
rect 45204 8520 45227 8551
rect 45097 8511 45155 8517
rect 45215 8517 45227 8520
rect 45261 8517 45273 8551
rect 45215 8511 45273 8517
rect 46198 8508 46204 8560
rect 46256 8548 46262 8560
rect 50249 8551 50307 8557
rect 46256 8520 49004 8548
rect 46256 8508 46262 8520
rect 32950 8440 32956 8492
rect 33008 8480 33014 8492
rect 33505 8483 33563 8489
rect 33505 8480 33517 8483
rect 33008 8452 33517 8480
rect 33008 8440 33014 8452
rect 33505 8449 33517 8452
rect 33551 8449 33563 8483
rect 33505 8443 33563 8449
rect 35253 8483 35311 8489
rect 35253 8449 35265 8483
rect 35299 8480 35311 8483
rect 36173 8483 36231 8489
rect 36173 8480 36185 8483
rect 35299 8452 36185 8480
rect 35299 8449 35311 8452
rect 35253 8443 35311 8449
rect 36173 8449 36185 8452
rect 36219 8449 36231 8483
rect 36173 8443 36231 8449
rect 33870 8412 33876 8424
rect 32232 8384 33876 8412
rect 33870 8372 33876 8384
rect 33928 8372 33934 8424
rect 35069 8415 35127 8421
rect 35069 8381 35081 8415
rect 35115 8412 35127 8415
rect 35342 8412 35348 8424
rect 35115 8384 35348 8412
rect 35115 8381 35127 8384
rect 35069 8375 35127 8381
rect 35342 8372 35348 8384
rect 35400 8372 35406 8424
rect 36188 8412 36216 8443
rect 36538 8440 36544 8492
rect 36596 8480 36602 8492
rect 37737 8483 37795 8489
rect 37737 8480 37749 8483
rect 36596 8452 37749 8480
rect 36596 8440 36602 8452
rect 37737 8449 37749 8452
rect 37783 8449 37795 8483
rect 38746 8480 38752 8492
rect 38707 8452 38752 8480
rect 37737 8443 37795 8449
rect 38746 8440 38752 8452
rect 38804 8440 38810 8492
rect 38933 8483 38991 8489
rect 38933 8449 38945 8483
rect 38979 8449 38991 8483
rect 38933 8443 38991 8449
rect 39577 8483 39635 8489
rect 39577 8449 39589 8483
rect 39623 8480 39635 8483
rect 39758 8480 39764 8492
rect 39623 8452 39764 8480
rect 39623 8449 39635 8452
rect 39577 8443 39635 8449
rect 36814 8412 36820 8424
rect 36188 8384 36820 8412
rect 36814 8372 36820 8384
rect 36872 8372 36878 8424
rect 36998 8372 37004 8424
rect 37056 8412 37062 8424
rect 38948 8412 38976 8443
rect 39758 8440 39764 8452
rect 39816 8440 39822 8492
rect 41506 8440 41512 8492
rect 41564 8480 41570 8492
rect 41601 8483 41659 8489
rect 41601 8480 41613 8483
rect 41564 8452 41613 8480
rect 41564 8440 41570 8452
rect 41601 8449 41613 8452
rect 41647 8449 41659 8483
rect 41601 8443 41659 8449
rect 41877 8483 41935 8489
rect 41877 8449 41889 8483
rect 41923 8480 41935 8483
rect 42334 8480 42340 8492
rect 41923 8452 42340 8480
rect 41923 8449 41935 8452
rect 41877 8443 41935 8449
rect 42334 8440 42340 8452
rect 42392 8440 42398 8492
rect 42610 8480 42616 8492
rect 42523 8452 42616 8480
rect 42610 8440 42616 8452
rect 42668 8440 42674 8492
rect 42702 8440 42708 8492
rect 42760 8480 42766 8492
rect 44910 8480 44916 8492
rect 42760 8452 42805 8480
rect 42996 8452 44916 8480
rect 42760 8440 42766 8452
rect 37056 8384 38976 8412
rect 37056 8372 37062 8384
rect 26200 8316 27752 8344
rect 27985 8347 28043 8353
rect 26200 8304 26206 8316
rect 27985 8313 27997 8347
rect 28031 8344 28043 8347
rect 28534 8344 28540 8356
rect 28031 8316 28540 8344
rect 28031 8313 28043 8316
rect 27985 8307 28043 8313
rect 28534 8304 28540 8316
rect 28592 8304 28598 8356
rect 29089 8347 29147 8353
rect 29089 8313 29101 8347
rect 29135 8344 29147 8347
rect 30374 8344 30380 8356
rect 29135 8316 30380 8344
rect 29135 8313 29147 8316
rect 29089 8307 29147 8313
rect 30374 8304 30380 8316
rect 30432 8304 30438 8356
rect 32306 8344 32312 8356
rect 32219 8316 32312 8344
rect 32306 8304 32312 8316
rect 32364 8344 32370 8356
rect 36354 8344 36360 8356
rect 32364 8316 33272 8344
rect 36315 8316 36360 8344
rect 32364 8304 32370 8316
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 9398 8276 9404 8288
rect 8996 8248 9404 8276
rect 8996 8236 9002 8248
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 21358 8236 21364 8288
rect 21416 8276 21422 8288
rect 27614 8276 27620 8288
rect 21416 8248 27620 8276
rect 21416 8236 21422 8248
rect 27614 8236 27620 8248
rect 27672 8236 27678 8288
rect 27801 8279 27859 8285
rect 27801 8245 27813 8279
rect 27847 8276 27859 8279
rect 27890 8276 27896 8288
rect 27847 8248 27896 8276
rect 27847 8245 27859 8248
rect 27801 8239 27859 8245
rect 27890 8236 27896 8248
rect 27948 8236 27954 8288
rect 28718 8236 28724 8288
rect 28776 8276 28782 8288
rect 28905 8279 28963 8285
rect 28905 8276 28917 8279
rect 28776 8248 28917 8276
rect 28776 8236 28782 8248
rect 28905 8245 28917 8248
rect 28951 8245 28963 8279
rect 28905 8239 28963 8245
rect 28994 8236 29000 8288
rect 29052 8276 29058 8288
rect 33134 8276 33140 8288
rect 29052 8248 33140 8276
rect 29052 8236 29058 8248
rect 33134 8236 33140 8248
rect 33192 8236 33198 8288
rect 33244 8276 33272 8316
rect 36354 8304 36360 8316
rect 36412 8304 36418 8356
rect 37918 8344 37924 8356
rect 37831 8316 37924 8344
rect 37918 8304 37924 8316
rect 37976 8344 37982 8356
rect 38562 8344 38568 8356
rect 37976 8316 38568 8344
rect 37976 8304 37982 8316
rect 38562 8304 38568 8316
rect 38620 8304 38626 8356
rect 38948 8344 38976 8384
rect 39114 8372 39120 8424
rect 39172 8412 39178 8424
rect 42628 8412 42656 8440
rect 42996 8412 43024 8452
rect 44910 8440 44916 8452
rect 44968 8440 44974 8492
rect 48774 8480 48780 8492
rect 45296 8452 48360 8480
rect 48735 8452 48780 8480
rect 39172 8384 43024 8412
rect 43073 8415 43131 8421
rect 39172 8372 39178 8384
rect 43073 8381 43085 8415
rect 43119 8381 43131 8415
rect 43073 8375 43131 8381
rect 41690 8344 41696 8356
rect 38948 8316 41696 8344
rect 41690 8304 41696 8316
rect 41748 8304 41754 8356
rect 41785 8347 41843 8353
rect 41785 8313 41797 8347
rect 41831 8344 41843 8347
rect 42429 8347 42487 8353
rect 42429 8344 42441 8347
rect 41831 8316 42441 8344
rect 41831 8313 41843 8316
rect 41785 8307 41843 8313
rect 42429 8313 42441 8316
rect 42475 8313 42487 8347
rect 43088 8344 43116 8375
rect 44542 8372 44548 8424
rect 44600 8412 44606 8424
rect 45296 8412 45324 8452
rect 44600 8384 45324 8412
rect 45373 8415 45431 8421
rect 44600 8372 44606 8384
rect 45373 8381 45385 8415
rect 45419 8412 45431 8415
rect 48222 8412 48228 8424
rect 45419 8384 48228 8412
rect 45419 8381 45431 8384
rect 45373 8375 45431 8381
rect 48222 8372 48228 8384
rect 48280 8372 48286 8424
rect 48332 8412 48360 8452
rect 48774 8440 48780 8452
rect 48832 8440 48838 8492
rect 48976 8489 49004 8520
rect 50249 8517 50261 8551
rect 50295 8517 50307 8551
rect 50249 8511 50307 8517
rect 48961 8483 49019 8489
rect 48961 8449 48973 8483
rect 49007 8449 49019 8483
rect 48961 8443 49019 8449
rect 49053 8483 49111 8489
rect 49053 8449 49065 8483
rect 49099 8480 49111 8483
rect 49602 8480 49608 8492
rect 49099 8452 49608 8480
rect 49099 8449 49111 8452
rect 49053 8443 49111 8449
rect 49602 8440 49608 8452
rect 49660 8440 49666 8492
rect 50264 8480 50292 8511
rect 52454 8480 52460 8492
rect 50264 8452 52460 8480
rect 52454 8440 52460 8452
rect 52512 8480 52518 8492
rect 52914 8480 52920 8492
rect 52512 8452 52920 8480
rect 52512 8440 52518 8452
rect 52914 8440 52920 8452
rect 52972 8440 52978 8492
rect 49694 8412 49700 8424
rect 48332 8384 49700 8412
rect 49694 8372 49700 8384
rect 49752 8372 49758 8424
rect 54846 8412 54852 8424
rect 51046 8384 54852 8412
rect 51046 8344 51074 8384
rect 54846 8372 54852 8384
rect 54904 8372 54910 8424
rect 43088 8316 51074 8344
rect 42429 8307 42487 8313
rect 33686 8276 33692 8288
rect 33244 8248 33692 8276
rect 33686 8236 33692 8248
rect 33744 8236 33750 8288
rect 35434 8276 35440 8288
rect 35395 8248 35440 8276
rect 35434 8236 35440 8248
rect 35492 8236 35498 8288
rect 35802 8236 35808 8288
rect 35860 8276 35866 8288
rect 36998 8276 37004 8288
rect 35860 8248 37004 8276
rect 35860 8236 35866 8248
rect 36998 8236 37004 8248
rect 37056 8236 37062 8288
rect 37182 8236 37188 8288
rect 37240 8276 37246 8288
rect 38749 8279 38807 8285
rect 38749 8276 38761 8279
rect 37240 8248 38761 8276
rect 37240 8236 37246 8248
rect 38749 8245 38761 8248
rect 38795 8245 38807 8279
rect 38749 8239 38807 8245
rect 41417 8279 41475 8285
rect 41417 8245 41429 8279
rect 41463 8276 41475 8279
rect 41506 8276 41512 8288
rect 41463 8248 41512 8276
rect 41463 8245 41475 8248
rect 41417 8239 41475 8245
rect 41506 8236 41512 8248
rect 41564 8236 41570 8288
rect 49418 8236 49424 8288
rect 49476 8276 49482 8288
rect 50433 8279 50491 8285
rect 50433 8276 50445 8279
rect 49476 8248 50445 8276
rect 49476 8236 49482 8248
rect 50433 8245 50445 8248
rect 50479 8245 50491 8279
rect 50433 8239 50491 8245
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 5994 8072 6000 8084
rect 4448 8044 5580 8072
rect 5955 8044 6000 8072
rect 2682 7964 2688 8016
rect 2740 8004 2746 8016
rect 4157 8007 4215 8013
rect 4157 8004 4169 8007
rect 2740 7976 4169 8004
rect 2740 7964 2746 7976
rect 4157 7973 4169 7976
rect 4203 7973 4215 8007
rect 4157 7967 4215 7973
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 4448 7936 4476 8044
rect 5552 8004 5580 8044
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 9309 8075 9367 8081
rect 9309 8041 9321 8075
rect 9355 8072 9367 8075
rect 10042 8072 10048 8084
rect 9355 8044 10048 8072
rect 9355 8041 9367 8044
rect 9309 8035 9367 8041
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8041 10195 8075
rect 13078 8072 13084 8084
rect 13039 8044 13084 8072
rect 10137 8035 10195 8041
rect 10152 8004 10180 8035
rect 13078 8032 13084 8044
rect 13136 8032 13142 8084
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14277 8075 14335 8081
rect 14277 8072 14289 8075
rect 14240 8044 14289 8072
rect 14240 8032 14246 8044
rect 14277 8041 14289 8044
rect 14323 8072 14335 8075
rect 17494 8072 17500 8084
rect 14323 8044 17500 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 19242 8072 19248 8084
rect 19203 8044 19248 8072
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 23106 8032 23112 8084
rect 23164 8072 23170 8084
rect 24670 8072 24676 8084
rect 23164 8044 24676 8072
rect 23164 8032 23170 8044
rect 24670 8032 24676 8044
rect 24728 8072 24734 8084
rect 25133 8075 25191 8081
rect 25133 8072 25145 8075
rect 24728 8044 25145 8072
rect 24728 8032 24734 8044
rect 25133 8041 25145 8044
rect 25179 8041 25191 8075
rect 25492 8075 25550 8081
rect 25492 8072 25504 8075
rect 25133 8035 25191 8041
rect 25424 8044 25504 8072
rect 5552 7976 6408 8004
rect 4614 7936 4620 7948
rect 1719 7908 4476 7936
rect 4575 7908 4620 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 6270 7868 6276 7880
rect 2731 7840 6276 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 3973 7803 4031 7809
rect 3973 7769 3985 7803
rect 4019 7769 4031 7803
rect 3973 7763 4031 7769
rect 4884 7803 4942 7809
rect 4884 7769 4896 7803
rect 4930 7800 4942 7803
rect 5258 7800 5264 7812
rect 4930 7772 5264 7800
rect 4930 7769 4942 7772
rect 4884 7763 4942 7769
rect 2866 7732 2872 7744
rect 2827 7704 2872 7732
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 3988 7732 4016 7763
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 6380 7800 6408 7976
rect 9048 7976 10180 8004
rect 7742 7896 7748 7948
rect 7800 7936 7806 7948
rect 8478 7936 8484 7948
rect 7800 7908 8484 7936
rect 7800 7896 7806 7908
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 8110 7868 8116 7880
rect 8071 7840 8116 7868
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 9048 7877 9076 7976
rect 13906 7964 13912 8016
rect 13964 8004 13970 8016
rect 17586 8004 17592 8016
rect 13964 7976 17592 8004
rect 13964 7964 13970 7976
rect 17586 7964 17592 7976
rect 17644 7964 17650 8016
rect 24302 7964 24308 8016
rect 24360 8004 24366 8016
rect 24360 7976 25360 8004
rect 24360 7964 24366 7976
rect 10962 7896 10968 7948
rect 11020 7936 11026 7948
rect 11701 7939 11759 7945
rect 11701 7936 11713 7939
rect 11020 7908 11713 7936
rect 11020 7896 11026 7908
rect 11701 7905 11713 7908
rect 11747 7905 11759 7939
rect 11701 7899 11759 7905
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7936 15715 7939
rect 15930 7936 15936 7948
rect 15703 7908 15936 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 15930 7896 15936 7908
rect 15988 7896 15994 7948
rect 19242 7896 19248 7948
rect 19300 7936 19306 7948
rect 21082 7936 21088 7948
rect 19300 7908 21088 7936
rect 19300 7896 19306 7908
rect 21082 7896 21088 7908
rect 21140 7936 21146 7948
rect 25130 7936 25136 7948
rect 21140 7908 25136 7936
rect 21140 7896 21146 7908
rect 25130 7896 25136 7908
rect 25188 7896 25194 7948
rect 9033 7871 9091 7877
rect 9033 7868 9045 7871
rect 8904 7840 9045 7868
rect 8904 7828 8910 7840
rect 9033 7837 9045 7840
rect 9079 7837 9091 7871
rect 10042 7868 10048 7880
rect 10003 7840 10048 7868
rect 9033 7831 9091 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 12250 7828 12256 7880
rect 12308 7868 12314 7880
rect 15286 7868 15292 7880
rect 12308 7840 15292 7868
rect 12308 7828 12314 7840
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 15470 7868 15476 7880
rect 15431 7840 15476 7868
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 15562 7828 15568 7880
rect 15620 7868 15626 7880
rect 15620 7840 15665 7868
rect 15620 7828 15626 7840
rect 15746 7828 15752 7880
rect 15804 7868 15810 7880
rect 19426 7868 19432 7880
rect 15804 7840 15849 7868
rect 19387 7840 19432 7868
rect 15804 7828 15810 7840
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7868 19763 7871
rect 19978 7868 19984 7880
rect 19751 7840 19984 7868
rect 19751 7837 19763 7840
rect 19705 7831 19763 7837
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 25222 7828 25228 7880
rect 25280 7828 25286 7880
rect 25332 7868 25360 7976
rect 25424 7936 25452 8044
rect 25492 8041 25504 8044
rect 25538 8041 25550 8075
rect 25492 8035 25550 8041
rect 27525 8075 27583 8081
rect 27525 8041 27537 8075
rect 27571 8041 27583 8075
rect 27525 8035 27583 8041
rect 27540 8004 27568 8035
rect 27614 8032 27620 8084
rect 27672 8072 27678 8084
rect 27672 8044 27844 8072
rect 27672 8032 27678 8044
rect 27709 8007 27767 8013
rect 27540 7976 27660 8004
rect 25590 7936 25596 7948
rect 25424 7908 25596 7936
rect 25590 7896 25596 7908
rect 25648 7896 25654 7948
rect 27632 7868 27660 7976
rect 27709 7973 27721 8007
rect 27755 7973 27767 8007
rect 27816 8004 27844 8044
rect 27890 8032 27896 8084
rect 27948 8072 27954 8084
rect 29733 8075 29791 8081
rect 29733 8072 29745 8075
rect 27948 8044 29745 8072
rect 27948 8032 27954 8044
rect 29733 8041 29745 8044
rect 29779 8041 29791 8075
rect 32582 8072 32588 8084
rect 29733 8035 29791 8041
rect 31036 8044 32588 8072
rect 31036 8004 31064 8044
rect 32582 8032 32588 8044
rect 32640 8032 32646 8084
rect 46474 8072 46480 8084
rect 32692 8044 46336 8072
rect 46435 8044 46480 8072
rect 27816 7976 31064 8004
rect 27709 7967 27767 7973
rect 27724 7936 27752 7967
rect 32692 7936 32720 8044
rect 33045 8007 33103 8013
rect 33045 7973 33057 8007
rect 33091 8004 33103 8007
rect 33318 8004 33324 8016
rect 33091 7976 33324 8004
rect 33091 7973 33103 7976
rect 33045 7967 33103 7973
rect 33318 7964 33324 7976
rect 33376 7964 33382 8016
rect 34790 7964 34796 8016
rect 34848 8004 34854 8016
rect 35069 8007 35127 8013
rect 35069 8004 35081 8007
rect 34848 7976 35081 8004
rect 34848 7964 34854 7976
rect 35069 7973 35081 7976
rect 35115 7973 35127 8007
rect 35069 7967 35127 7973
rect 35526 7964 35532 8016
rect 35584 8004 35590 8016
rect 38378 8004 38384 8016
rect 35584 7976 38384 8004
rect 35584 7964 35590 7976
rect 38378 7964 38384 7976
rect 38436 7964 38442 8016
rect 38746 8004 38752 8016
rect 38707 7976 38752 8004
rect 38746 7964 38752 7976
rect 38804 7964 38810 8016
rect 42426 7964 42432 8016
rect 42484 8004 42490 8016
rect 42613 8007 42671 8013
rect 42613 8004 42625 8007
rect 42484 7976 42625 8004
rect 42484 7964 42490 7976
rect 42613 7973 42625 7976
rect 42659 7973 42671 8007
rect 46308 8004 46336 8044
rect 46474 8032 46480 8044
rect 46532 8032 46538 8084
rect 49694 8032 49700 8084
rect 49752 8072 49758 8084
rect 52917 8075 52975 8081
rect 52917 8072 52929 8075
rect 49752 8044 52929 8072
rect 49752 8032 49758 8044
rect 52917 8041 52929 8044
rect 52963 8041 52975 8075
rect 52917 8035 52975 8041
rect 49418 8004 49424 8016
rect 46308 7976 49424 8004
rect 42613 7967 42671 7973
rect 49418 7964 49424 7976
rect 49476 7964 49482 8016
rect 37734 7936 37740 7948
rect 27724 7908 31156 7936
rect 27890 7868 27896 7880
rect 25332 7840 25452 7868
rect 9674 7800 9680 7812
rect 6380 7772 9680 7800
rect 9674 7760 9680 7772
rect 9732 7760 9738 7812
rect 11968 7803 12026 7809
rect 11968 7769 11980 7803
rect 12014 7800 12026 7803
rect 12618 7800 12624 7812
rect 12014 7772 12624 7800
rect 12014 7769 12026 7772
rect 11968 7763 12026 7769
rect 12618 7760 12624 7772
rect 12676 7760 12682 7812
rect 14090 7800 14096 7812
rect 14051 7772 14096 7800
rect 14090 7760 14096 7772
rect 14148 7760 14154 7812
rect 14274 7760 14280 7812
rect 14332 7809 14338 7812
rect 14332 7803 14351 7809
rect 14339 7769 14351 7803
rect 14332 7763 14351 7769
rect 19613 7803 19671 7809
rect 19613 7769 19625 7803
rect 19659 7800 19671 7803
rect 20070 7800 20076 7812
rect 19659 7772 20076 7800
rect 19659 7769 19671 7772
rect 19613 7763 19671 7769
rect 14332 7760 14338 7763
rect 20070 7760 20076 7772
rect 20128 7760 20134 7812
rect 24486 7800 24492 7812
rect 24447 7772 24492 7800
rect 24486 7760 24492 7772
rect 24544 7760 24550 7812
rect 24705 7803 24763 7809
rect 24705 7769 24717 7803
rect 24751 7800 24763 7803
rect 25240 7800 25268 7828
rect 24751 7772 25268 7800
rect 25317 7803 25375 7809
rect 24751 7769 24763 7772
rect 24705 7763 24763 7769
rect 25317 7769 25329 7803
rect 25363 7800 25375 7803
rect 25424 7800 25452 7840
rect 25363 7772 25452 7800
rect 25532 7840 27594 7868
rect 27632 7840 27896 7868
rect 25363 7769 25375 7772
rect 25317 7763 25375 7769
rect 5534 7732 5540 7744
rect 3988 7704 5540 7732
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 8202 7732 8208 7744
rect 8163 7704 8208 7732
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 9490 7732 9496 7744
rect 8352 7704 9496 7732
rect 8352 7692 8358 7704
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 10226 7692 10232 7744
rect 10284 7732 10290 7744
rect 10505 7735 10563 7741
rect 10505 7732 10517 7735
rect 10284 7704 10517 7732
rect 10284 7692 10290 7704
rect 10505 7701 10517 7704
rect 10551 7732 10563 7735
rect 12434 7732 12440 7744
rect 10551 7704 12440 7732
rect 10551 7701 10563 7704
rect 10505 7695 10563 7701
rect 12434 7692 12440 7704
rect 12492 7692 12498 7744
rect 14458 7732 14464 7744
rect 14419 7704 14464 7732
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 15289 7735 15347 7741
rect 15289 7732 15301 7735
rect 14608 7704 15301 7732
rect 14608 7692 14614 7704
rect 15289 7701 15301 7704
rect 15335 7701 15347 7735
rect 15289 7695 15347 7701
rect 16206 7692 16212 7744
rect 16264 7732 16270 7744
rect 19334 7732 19340 7744
rect 16264 7704 19340 7732
rect 16264 7692 16270 7704
rect 19334 7692 19340 7704
rect 19392 7732 19398 7744
rect 20530 7732 20536 7744
rect 19392 7704 20536 7732
rect 19392 7692 19398 7704
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 21634 7692 21640 7744
rect 21692 7732 21698 7744
rect 24118 7732 24124 7744
rect 21692 7704 24124 7732
rect 21692 7692 21698 7704
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 24854 7732 24860 7744
rect 24815 7704 24860 7732
rect 24854 7692 24860 7704
rect 24912 7692 24918 7744
rect 25406 7692 25412 7744
rect 25464 7732 25470 7744
rect 25532 7741 25560 7840
rect 26234 7800 26240 7812
rect 26195 7772 26240 7800
rect 26234 7760 26240 7772
rect 26292 7760 26298 7812
rect 27341 7803 27399 7809
rect 27341 7769 27353 7803
rect 27387 7800 27399 7803
rect 27430 7800 27436 7812
rect 27387 7772 27436 7800
rect 27387 7769 27399 7772
rect 27341 7763 27399 7769
rect 27430 7760 27436 7772
rect 27488 7760 27494 7812
rect 27566 7800 27594 7840
rect 27890 7828 27896 7840
rect 27948 7828 27954 7880
rect 28166 7868 28172 7880
rect 28127 7840 28172 7868
rect 28166 7828 28172 7840
rect 28224 7828 28230 7880
rect 28445 7871 28503 7877
rect 28445 7837 28457 7871
rect 28491 7837 28503 7871
rect 28445 7831 28503 7837
rect 31021 7871 31079 7877
rect 31021 7837 31033 7871
rect 31067 7837 31079 7871
rect 31128 7868 31156 7908
rect 32508 7908 32720 7936
rect 32876 7908 37740 7936
rect 32508 7868 32536 7908
rect 31128 7840 32536 7868
rect 31021 7831 31079 7837
rect 27706 7800 27712 7812
rect 27566 7772 27712 7800
rect 27706 7760 27712 7772
rect 27764 7760 27770 7812
rect 28460 7800 28488 7831
rect 29549 7803 29607 7809
rect 29549 7800 29561 7803
rect 28000 7772 28488 7800
rect 28552 7772 29561 7800
rect 28000 7744 28028 7772
rect 25517 7735 25575 7741
rect 25517 7732 25529 7735
rect 25464 7704 25529 7732
rect 25464 7692 25470 7704
rect 25517 7701 25529 7704
rect 25563 7701 25575 7735
rect 25682 7732 25688 7744
rect 25643 7704 25688 7732
rect 25517 7695 25575 7701
rect 25682 7692 25688 7704
rect 25740 7692 25746 7744
rect 26326 7732 26332 7744
rect 26287 7704 26332 7732
rect 26326 7692 26332 7704
rect 26384 7692 26390 7744
rect 27551 7735 27609 7741
rect 27551 7701 27563 7735
rect 27597 7732 27609 7735
rect 27982 7732 27988 7744
rect 27597 7704 27988 7732
rect 27597 7701 27609 7704
rect 27551 7695 27609 7701
rect 27982 7692 27988 7704
rect 28040 7692 28046 7744
rect 28258 7692 28264 7744
rect 28316 7732 28322 7744
rect 28552 7732 28580 7772
rect 29549 7769 29561 7772
rect 29595 7769 29607 7803
rect 29549 7763 29607 7769
rect 28316 7704 28580 7732
rect 28316 7692 28322 7704
rect 28902 7692 28908 7744
rect 28960 7732 28966 7744
rect 29749 7735 29807 7741
rect 29749 7732 29761 7735
rect 28960 7704 29761 7732
rect 28960 7692 28966 7704
rect 29749 7701 29761 7704
rect 29795 7701 29807 7735
rect 29749 7695 29807 7701
rect 29917 7735 29975 7741
rect 29917 7701 29929 7735
rect 29963 7732 29975 7735
rect 30098 7732 30104 7744
rect 29963 7704 30104 7732
rect 29963 7701 29975 7704
rect 29917 7695 29975 7701
rect 30098 7692 30104 7704
rect 30156 7692 30162 7744
rect 31036 7732 31064 7831
rect 32674 7828 32680 7880
rect 32732 7868 32738 7880
rect 32876 7877 32904 7908
rect 37734 7896 37740 7908
rect 37792 7896 37798 7948
rect 39114 7936 39120 7948
rect 37844 7908 39120 7936
rect 32861 7871 32919 7877
rect 32861 7868 32873 7871
rect 32732 7840 32873 7868
rect 32732 7828 32738 7840
rect 32861 7837 32873 7840
rect 32907 7837 32919 7871
rect 32861 7831 32919 7837
rect 34701 7871 34759 7877
rect 34701 7837 34713 7871
rect 34747 7868 34759 7871
rect 35066 7868 35072 7880
rect 34747 7840 35072 7868
rect 34747 7837 34759 7840
rect 34701 7831 34759 7837
rect 35066 7828 35072 7840
rect 35124 7868 35130 7880
rect 35434 7868 35440 7880
rect 35124 7840 35440 7868
rect 35124 7828 35130 7840
rect 35434 7828 35440 7840
rect 35492 7828 35498 7880
rect 37844 7877 37872 7908
rect 39114 7896 39120 7908
rect 39172 7896 39178 7948
rect 40034 7896 40040 7948
rect 40092 7936 40098 7948
rect 41230 7936 41236 7948
rect 40092 7908 41236 7936
rect 40092 7896 40098 7908
rect 41230 7896 41236 7908
rect 41288 7896 41294 7948
rect 42886 7896 42892 7948
rect 42944 7936 42950 7948
rect 45281 7939 45339 7945
rect 45281 7936 45293 7939
rect 42944 7908 45293 7936
rect 42944 7896 42950 7908
rect 45281 7905 45293 7908
rect 45327 7936 45339 7939
rect 45462 7936 45468 7948
rect 45327 7908 45468 7936
rect 45327 7905 45339 7908
rect 45281 7899 45339 7905
rect 45462 7896 45468 7908
rect 45520 7896 45526 7948
rect 37829 7871 37887 7877
rect 37829 7837 37841 7871
rect 37875 7837 37887 7871
rect 38010 7868 38016 7880
rect 37971 7840 38016 7868
rect 37829 7831 37887 7837
rect 38010 7828 38016 7840
rect 38068 7828 38074 7880
rect 38562 7868 38568 7880
rect 38523 7840 38568 7868
rect 38562 7828 38568 7840
rect 38620 7828 38626 7880
rect 41506 7877 41512 7880
rect 41500 7868 41512 7877
rect 41467 7840 41512 7868
rect 41500 7831 41512 7840
rect 41506 7828 41512 7831
rect 41564 7828 41570 7880
rect 42334 7828 42340 7880
rect 42392 7868 42398 7880
rect 44174 7868 44180 7880
rect 42392 7840 44180 7868
rect 42392 7828 42398 7840
rect 44174 7828 44180 7840
rect 44232 7828 44238 7880
rect 44266 7828 44272 7880
rect 44324 7868 44330 7880
rect 45005 7871 45063 7877
rect 45005 7868 45017 7871
rect 44324 7840 45017 7868
rect 44324 7828 44330 7840
rect 45005 7837 45017 7840
rect 45051 7837 45063 7871
rect 52730 7868 52736 7880
rect 52691 7840 52736 7868
rect 45005 7831 45063 7837
rect 52730 7828 52736 7840
rect 52788 7828 52794 7880
rect 53006 7828 53012 7880
rect 53064 7868 53070 7880
rect 53064 7840 53109 7868
rect 53064 7828 53070 7840
rect 31288 7803 31346 7809
rect 31288 7769 31300 7803
rect 31334 7800 31346 7803
rect 32122 7800 32128 7812
rect 31334 7772 32128 7800
rect 31334 7769 31346 7772
rect 31288 7763 31346 7769
rect 32122 7760 32128 7772
rect 32180 7760 32186 7812
rect 32950 7800 32956 7812
rect 32416 7772 32956 7800
rect 31846 7732 31852 7744
rect 31036 7704 31852 7732
rect 31846 7692 31852 7704
rect 31904 7692 31910 7744
rect 32416 7741 32444 7772
rect 32950 7760 32956 7772
rect 33008 7760 33014 7812
rect 34790 7760 34796 7812
rect 34848 7800 34854 7812
rect 34885 7803 34943 7809
rect 34885 7800 34897 7803
rect 34848 7772 34897 7800
rect 34848 7760 34854 7772
rect 34885 7769 34897 7772
rect 34931 7769 34943 7803
rect 34885 7763 34943 7769
rect 34983 7772 38036 7800
rect 32401 7735 32459 7741
rect 32401 7701 32413 7735
rect 32447 7701 32459 7735
rect 32401 7695 32459 7701
rect 32582 7692 32588 7744
rect 32640 7732 32646 7744
rect 34983 7732 35011 7772
rect 32640 7704 35011 7732
rect 32640 7692 32646 7704
rect 35250 7692 35256 7744
rect 35308 7732 35314 7744
rect 35526 7732 35532 7744
rect 35308 7704 35532 7732
rect 35308 7692 35314 7704
rect 35526 7692 35532 7704
rect 35584 7732 35590 7744
rect 37182 7732 37188 7744
rect 35584 7704 37188 7732
rect 35584 7692 35590 7704
rect 37182 7692 37188 7704
rect 37240 7692 37246 7744
rect 37274 7692 37280 7744
rect 37332 7732 37338 7744
rect 37921 7735 37979 7741
rect 37921 7732 37933 7735
rect 37332 7704 37933 7732
rect 37332 7692 37338 7704
rect 37921 7701 37933 7704
rect 37967 7701 37979 7735
rect 38008 7732 38036 7772
rect 38102 7760 38108 7812
rect 38160 7800 38166 7812
rect 45922 7800 45928 7812
rect 38160 7772 45928 7800
rect 38160 7760 38166 7772
rect 45922 7760 45928 7772
rect 45980 7760 45986 7812
rect 46014 7760 46020 7812
rect 46072 7800 46078 7812
rect 46385 7803 46443 7809
rect 46385 7800 46397 7803
rect 46072 7772 46397 7800
rect 46072 7760 46078 7772
rect 46385 7769 46397 7772
rect 46431 7769 46443 7803
rect 46385 7763 46443 7769
rect 42518 7732 42524 7744
rect 38008 7704 42524 7732
rect 37921 7695 37979 7701
rect 42518 7692 42524 7704
rect 42576 7692 42582 7744
rect 52546 7732 52552 7744
rect 52507 7704 52552 7732
rect 52546 7692 52552 7704
rect 52604 7692 52610 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2593 7531 2651 7537
rect 2593 7528 2605 7531
rect 2096 7500 2605 7528
rect 2096 7488 2102 7500
rect 2593 7497 2605 7500
rect 2639 7497 2651 7531
rect 5258 7528 5264 7540
rect 5219 7500 5264 7528
rect 2593 7491 2651 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 12618 7528 12624 7540
rect 5460 7500 12434 7528
rect 12579 7500 12624 7528
rect 2501 7463 2559 7469
rect 2501 7429 2513 7463
rect 2547 7460 2559 7463
rect 4890 7460 4896 7472
rect 2547 7432 4896 7460
rect 2547 7429 2559 7432
rect 2501 7423 2559 7429
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 1486 7392 1492 7404
rect 1447 7364 1492 7392
rect 1486 7352 1492 7364
rect 1544 7352 1550 7404
rect 3510 7392 3516 7404
rect 3471 7364 3516 7392
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 5460 7401 5488 7500
rect 5629 7463 5687 7469
rect 5629 7429 5641 7463
rect 5675 7460 5687 7463
rect 5994 7460 6000 7472
rect 5675 7432 6000 7460
rect 5675 7429 5687 7432
rect 5629 7423 5687 7429
rect 5994 7420 6000 7432
rect 6052 7420 6058 7472
rect 7653 7463 7711 7469
rect 7653 7429 7665 7463
rect 7699 7460 7711 7463
rect 7699 7432 7972 7460
rect 7699 7429 7711 7432
rect 7653 7423 7711 7429
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 7742 7392 7748 7404
rect 5776 7364 5821 7392
rect 7703 7364 7748 7392
rect 5776 7352 5782 7364
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 7944 7392 7972 7432
rect 8202 7420 8208 7472
rect 8260 7420 8266 7472
rect 11885 7463 11943 7469
rect 11885 7429 11897 7463
rect 11931 7460 11943 7463
rect 12250 7460 12256 7472
rect 11931 7432 12256 7460
rect 11931 7429 11943 7432
rect 11885 7423 11943 7429
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 12406 7460 12434 7500
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 12989 7531 13047 7537
rect 12989 7497 13001 7531
rect 13035 7528 13047 7531
rect 13078 7528 13084 7540
rect 13035 7500 13084 7528
rect 13035 7497 13047 7500
rect 12989 7491 13047 7497
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 14090 7488 14096 7540
rect 14148 7528 14154 7540
rect 14148 7500 15424 7528
rect 14148 7488 14154 7500
rect 14550 7460 14556 7472
rect 12406 7432 14556 7460
rect 14550 7420 14556 7432
rect 14608 7420 14614 7472
rect 15396 7460 15424 7500
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 15528 7500 16681 7528
rect 15528 7488 15534 7500
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 16669 7491 16727 7497
rect 19455 7531 19513 7537
rect 19455 7497 19467 7531
rect 19501 7528 19513 7531
rect 20457 7531 20515 7537
rect 20457 7528 20469 7531
rect 19501 7500 20469 7528
rect 19501 7497 19513 7500
rect 19455 7491 19513 7497
rect 20457 7497 20469 7500
rect 20503 7528 20515 7531
rect 22830 7528 22836 7540
rect 20503 7500 22836 7528
rect 20503 7497 20515 7500
rect 20457 7491 20515 7497
rect 22830 7488 22836 7500
rect 22888 7488 22894 7540
rect 24854 7528 24860 7540
rect 22940 7500 24860 7528
rect 19242 7460 19248 7472
rect 15396 7432 19248 7460
rect 19242 7420 19248 7432
rect 19300 7460 19306 7472
rect 20257 7463 20315 7469
rect 20257 7460 20269 7463
rect 19300 7432 20269 7460
rect 19300 7420 19306 7432
rect 20257 7429 20269 7432
rect 20303 7429 20315 7463
rect 20257 7423 20315 7429
rect 8220 7392 8248 7420
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 7944 7364 8769 7392
rect 8757 7361 8769 7364
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9079 7364 10180 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 2682 7324 2688 7336
rect 2643 7296 2688 7324
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 6454 7324 6460 7336
rect 5592 7296 6460 7324
rect 5592 7284 5598 7296
rect 6454 7284 6460 7296
rect 6512 7324 6518 7336
rect 8113 7327 8171 7333
rect 8113 7324 8125 7327
rect 6512 7296 8125 7324
rect 6512 7284 6518 7296
rect 8113 7293 8125 7296
rect 8159 7293 8171 7327
rect 8113 7287 8171 7293
rect 8205 7327 8263 7333
rect 8205 7293 8217 7327
rect 8251 7324 8263 7327
rect 9214 7324 9220 7336
rect 8251 7296 9220 7324
rect 8251 7293 8263 7296
rect 8205 7287 8263 7293
rect 9214 7284 9220 7296
rect 9272 7284 9278 7336
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 10045 7327 10103 7333
rect 10045 7324 10057 7327
rect 9548 7296 10057 7324
rect 9548 7284 9554 7296
rect 10045 7293 10057 7296
rect 10091 7293 10103 7327
rect 10152 7324 10180 7364
rect 10226 7352 10232 7404
rect 10284 7392 10290 7404
rect 10284 7364 10329 7392
rect 10284 7352 10290 7364
rect 10410 7352 10416 7404
rect 10468 7392 10474 7404
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 10468 7364 11529 7392
rect 10468 7352 10474 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 12805 7395 12863 7401
rect 11747 7364 12572 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 12434 7324 12440 7336
rect 10152 7296 12440 7324
rect 10045 7287 10103 7293
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 9582 7216 9588 7268
rect 9640 7256 9646 7268
rect 9640 7228 12434 7256
rect 9640 7216 9646 7228
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 2866 7188 2872 7200
rect 2179 7160 2872 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 3326 7188 3332 7200
rect 3287 7160 3332 7188
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 10410 7188 10416 7200
rect 10371 7160 10416 7188
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 12406 7188 12434 7228
rect 12544 7188 12572 7364
rect 12805 7361 12817 7395
rect 12851 7361 12863 7395
rect 12805 7355 12863 7361
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13630 7392 13636 7404
rect 13127 7364 13636 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 12820 7324 12848 7355
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 15565 7395 15623 7401
rect 15565 7392 15577 7395
rect 15212 7364 15577 7392
rect 15212 7336 15240 7364
rect 15565 7361 15577 7364
rect 15611 7361 15623 7395
rect 16850 7392 16856 7404
rect 16811 7364 16856 7392
rect 15565 7355 15623 7361
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 19150 7392 19156 7404
rect 17083 7364 19156 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 22370 7392 22376 7404
rect 19260 7364 22376 7392
rect 14458 7324 14464 7336
rect 12820 7296 14464 7324
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 15194 7284 15200 7336
rect 15252 7284 15258 7336
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7324 15347 7327
rect 16666 7324 16672 7336
rect 15335 7296 16672 7324
rect 15335 7293 15347 7296
rect 15289 7287 15347 7293
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 16945 7327 17003 7333
rect 16945 7293 16957 7327
rect 16991 7293 17003 7327
rect 16945 7287 17003 7293
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7324 17187 7327
rect 17402 7324 17408 7336
rect 17175 7296 17408 7324
rect 17175 7293 17187 7296
rect 17129 7287 17187 7293
rect 16298 7216 16304 7268
rect 16356 7256 16362 7268
rect 16960 7256 16988 7287
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 17034 7256 17040 7268
rect 16356 7228 17040 7256
rect 16356 7216 16362 7228
rect 17034 7216 17040 7228
rect 17092 7216 17098 7268
rect 19260 7188 19288 7364
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 22940 7401 22968 7500
rect 24854 7488 24860 7500
rect 24912 7488 24918 7540
rect 25130 7528 25136 7540
rect 25091 7500 25136 7528
rect 25130 7488 25136 7500
rect 25188 7488 25194 7540
rect 25222 7488 25228 7540
rect 25280 7528 25286 7540
rect 26234 7528 26240 7540
rect 25280 7500 26240 7528
rect 25280 7488 25286 7500
rect 26234 7488 26240 7500
rect 26292 7488 26298 7540
rect 28166 7488 28172 7540
rect 28224 7528 28230 7540
rect 28810 7528 28816 7540
rect 28224 7500 28816 7528
rect 28224 7488 28230 7500
rect 28810 7488 28816 7500
rect 28868 7528 28874 7540
rect 30190 7528 30196 7540
rect 28868 7500 30196 7528
rect 28868 7488 28874 7500
rect 30190 7488 30196 7500
rect 30248 7488 30254 7540
rect 32122 7528 32128 7540
rect 32083 7500 32128 7528
rect 32122 7488 32128 7500
rect 32180 7488 32186 7540
rect 33870 7488 33876 7540
rect 33928 7528 33934 7540
rect 34330 7528 34336 7540
rect 33928 7500 34336 7528
rect 33928 7488 33934 7500
rect 34330 7488 34336 7500
rect 34388 7488 34394 7540
rect 34440 7500 37044 7528
rect 23109 7463 23167 7469
rect 23109 7429 23121 7463
rect 23155 7460 23167 7463
rect 23382 7460 23388 7472
rect 23155 7432 23388 7460
rect 23155 7429 23167 7432
rect 23109 7423 23167 7429
rect 23382 7420 23388 7432
rect 23440 7420 23446 7472
rect 24118 7460 24124 7472
rect 24079 7432 24124 7460
rect 24118 7420 24124 7432
rect 24176 7420 24182 7472
rect 24337 7463 24395 7469
rect 24337 7429 24349 7463
rect 24383 7460 24395 7463
rect 25406 7460 25412 7472
rect 24383 7432 25412 7460
rect 24383 7429 24395 7432
rect 24337 7423 24395 7429
rect 25406 7420 25412 7432
rect 25464 7420 25470 7472
rect 25498 7420 25504 7472
rect 25556 7460 25562 7472
rect 26510 7460 26516 7472
rect 25556 7432 26516 7460
rect 25556 7420 25562 7432
rect 26510 7420 26516 7432
rect 26568 7420 26574 7472
rect 27801 7463 27859 7469
rect 27801 7429 27813 7463
rect 27847 7429 27859 7463
rect 27982 7460 27988 7472
rect 27943 7432 27988 7460
rect 27801 7423 27859 7429
rect 22925 7395 22983 7401
rect 22925 7361 22937 7395
rect 22971 7361 22983 7395
rect 23198 7392 23204 7404
rect 23159 7364 23204 7392
rect 22925 7355 22983 7361
rect 23198 7352 23204 7364
rect 23256 7352 23262 7404
rect 25041 7395 25099 7401
rect 25041 7361 25053 7395
rect 25087 7392 25099 7395
rect 25222 7392 25228 7404
rect 25087 7364 25228 7392
rect 25087 7361 25099 7364
rect 25041 7355 25099 7361
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 25590 7352 25596 7404
rect 25648 7392 25654 7404
rect 25685 7395 25743 7401
rect 25685 7392 25697 7395
rect 25648 7364 25697 7392
rect 25648 7352 25654 7364
rect 25685 7361 25697 7364
rect 25731 7361 25743 7395
rect 27816 7392 27844 7423
rect 27982 7420 27988 7432
rect 28040 7420 28046 7472
rect 28442 7420 28448 7472
rect 28500 7460 28506 7472
rect 28721 7463 28779 7469
rect 28721 7460 28733 7463
rect 28500 7432 28733 7460
rect 28500 7420 28506 7432
rect 28721 7429 28733 7432
rect 28767 7429 28779 7463
rect 28721 7423 28779 7429
rect 28902 7420 28908 7472
rect 28960 7469 28966 7472
rect 28960 7463 28979 7469
rect 28967 7429 28979 7463
rect 30926 7460 30932 7472
rect 28960 7423 28979 7429
rect 30208 7432 30932 7460
rect 28960 7420 28966 7423
rect 25685 7355 25743 7361
rect 25792 7364 27844 7392
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 19484 7296 19656 7324
rect 19484 7284 19490 7296
rect 19628 7265 19656 7296
rect 20530 7284 20536 7336
rect 20588 7324 20594 7336
rect 25792 7324 25820 7364
rect 29914 7352 29920 7404
rect 29972 7392 29978 7404
rect 30208 7401 30236 7432
rect 30926 7420 30932 7432
rect 30984 7420 30990 7472
rect 34440 7460 34468 7500
rect 36906 7460 36912 7472
rect 32232 7432 34468 7460
rect 35176 7432 36912 7460
rect 30193 7395 30251 7401
rect 30193 7392 30205 7395
rect 29972 7364 30205 7392
rect 29972 7352 29978 7364
rect 30193 7361 30205 7364
rect 30239 7361 30251 7395
rect 30193 7355 30251 7361
rect 30377 7395 30435 7401
rect 30377 7361 30389 7395
rect 30423 7392 30435 7395
rect 30466 7392 30472 7404
rect 30423 7364 30472 7392
rect 30423 7361 30435 7364
rect 30377 7355 30435 7361
rect 30466 7352 30472 7364
rect 30524 7352 30530 7404
rect 31110 7392 31116 7404
rect 31071 7364 31116 7392
rect 31110 7352 31116 7364
rect 31168 7352 31174 7404
rect 27706 7324 27712 7336
rect 20588 7296 25820 7324
rect 26160 7296 27712 7324
rect 20588 7284 20594 7296
rect 19613 7259 19671 7265
rect 19613 7225 19625 7259
rect 19659 7256 19671 7259
rect 19978 7256 19984 7268
rect 19659 7228 19984 7256
rect 19659 7225 19671 7228
rect 19613 7219 19671 7225
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 20162 7216 20168 7268
rect 20220 7256 20226 7268
rect 20625 7259 20683 7265
rect 20625 7256 20637 7259
rect 20220 7228 20637 7256
rect 20220 7216 20226 7228
rect 20625 7225 20637 7228
rect 20671 7225 20683 7259
rect 20625 7219 20683 7225
rect 21266 7216 21272 7268
rect 21324 7256 21330 7268
rect 24394 7256 24400 7268
rect 21324 7228 24400 7256
rect 21324 7216 21330 7228
rect 12406 7160 19288 7188
rect 19334 7148 19340 7200
rect 19392 7188 19398 7200
rect 19429 7191 19487 7197
rect 19429 7188 19441 7191
rect 19392 7160 19441 7188
rect 19392 7148 19398 7160
rect 19429 7157 19441 7160
rect 19475 7157 19487 7191
rect 19429 7151 19487 7157
rect 19889 7191 19947 7197
rect 19889 7157 19901 7191
rect 19935 7188 19947 7191
rect 20254 7188 20260 7200
rect 19935 7160 20260 7188
rect 19935 7157 19947 7160
rect 19889 7151 19947 7157
rect 20254 7148 20260 7160
rect 20312 7188 20318 7200
rect 20441 7191 20499 7197
rect 20441 7188 20453 7191
rect 20312 7160 20453 7188
rect 20312 7148 20318 7160
rect 20441 7157 20453 7160
rect 20487 7188 20499 7191
rect 22462 7188 22468 7200
rect 20487 7160 22468 7188
rect 20487 7157 20499 7160
rect 20441 7151 20499 7157
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 22738 7188 22744 7200
rect 22699 7160 22744 7188
rect 22738 7148 22744 7160
rect 22796 7148 22802 7200
rect 24320 7197 24348 7228
rect 24394 7216 24400 7228
rect 24452 7216 24458 7268
rect 26160 7256 26188 7296
rect 27706 7284 27712 7296
rect 27764 7284 27770 7336
rect 27798 7284 27804 7336
rect 27856 7324 27862 7336
rect 32232 7324 32260 7432
rect 32309 7395 32367 7401
rect 32309 7361 32321 7395
rect 32355 7392 32367 7395
rect 34882 7392 34888 7404
rect 32355 7364 34888 7392
rect 32355 7361 32367 7364
rect 32309 7355 32367 7361
rect 34882 7352 34888 7364
rect 34940 7352 34946 7404
rect 35066 7392 35072 7404
rect 35027 7364 35072 7392
rect 35066 7352 35072 7364
rect 35124 7352 35130 7404
rect 35176 7401 35204 7432
rect 36906 7420 36912 7432
rect 36964 7420 36970 7472
rect 37016 7460 37044 7500
rect 37090 7488 37096 7540
rect 37148 7528 37154 7540
rect 42334 7528 42340 7540
rect 37148 7500 42340 7528
rect 37148 7488 37154 7500
rect 42334 7488 42340 7500
rect 42392 7488 42398 7540
rect 42444 7500 43576 7528
rect 41966 7460 41972 7472
rect 37016 7432 41972 7460
rect 41966 7420 41972 7432
rect 42024 7420 42030 7472
rect 35161 7395 35219 7401
rect 35161 7361 35173 7395
rect 35207 7361 35219 7395
rect 35161 7355 35219 7361
rect 35250 7352 35256 7404
rect 35308 7392 35314 7404
rect 35437 7395 35495 7401
rect 35308 7364 35353 7392
rect 35308 7352 35314 7364
rect 35437 7361 35449 7395
rect 35483 7392 35495 7395
rect 36170 7392 36176 7404
rect 35483 7364 36176 7392
rect 35483 7361 35495 7364
rect 35437 7355 35495 7361
rect 36170 7352 36176 7364
rect 36228 7352 36234 7404
rect 37458 7352 37464 7404
rect 37516 7392 37522 7404
rect 37993 7395 38051 7401
rect 37993 7392 38005 7395
rect 37516 7364 38005 7392
rect 37516 7352 37522 7364
rect 37993 7361 38005 7364
rect 38039 7361 38051 7395
rect 37993 7355 38051 7361
rect 38378 7352 38384 7404
rect 38436 7392 38442 7404
rect 42444 7392 42472 7500
rect 42518 7420 42524 7472
rect 42576 7460 42582 7472
rect 42797 7463 42855 7469
rect 42797 7460 42809 7463
rect 42576 7432 42809 7460
rect 42576 7420 42582 7432
rect 42797 7429 42809 7432
rect 42843 7460 42855 7463
rect 43349 7463 43407 7469
rect 43349 7460 43361 7463
rect 42843 7432 43361 7460
rect 42843 7429 42855 7432
rect 42797 7423 42855 7429
rect 43349 7429 43361 7432
rect 43395 7429 43407 7463
rect 43349 7423 43407 7429
rect 42610 7392 42616 7404
rect 38436 7364 42472 7392
rect 42571 7364 42616 7392
rect 38436 7352 38442 7364
rect 42610 7352 42616 7364
rect 42668 7352 42674 7404
rect 42702 7352 42708 7404
rect 42760 7392 42766 7404
rect 42760 7364 42805 7392
rect 42760 7352 42766 7364
rect 42886 7352 42892 7404
rect 42944 7401 42950 7404
rect 42944 7395 42973 7401
rect 42961 7361 42973 7395
rect 43548 7392 43576 7500
rect 45922 7488 45928 7540
rect 45980 7528 45986 7540
rect 54846 7528 54852 7540
rect 45980 7500 46428 7528
rect 54807 7500 54852 7528
rect 45980 7488 45986 7500
rect 46198 7460 46204 7472
rect 46159 7432 46204 7460
rect 46198 7420 46204 7432
rect 46256 7420 46262 7472
rect 44361 7395 44419 7401
rect 44361 7392 44373 7395
rect 43548 7364 44373 7392
rect 42944 7355 42973 7361
rect 44361 7361 44373 7364
rect 44407 7361 44419 7395
rect 44542 7392 44548 7404
rect 44503 7364 44548 7392
rect 44361 7355 44419 7361
rect 42944 7352 42950 7355
rect 32582 7324 32588 7336
rect 27856 7296 32260 7324
rect 32543 7296 32588 7324
rect 27856 7284 27862 7296
rect 32582 7284 32588 7296
rect 32640 7284 32646 7336
rect 33134 7284 33140 7336
rect 33192 7324 33198 7336
rect 37734 7324 37740 7336
rect 33192 7296 37228 7324
rect 37695 7296 37740 7324
rect 33192 7284 33198 7296
rect 25332 7228 26188 7256
rect 24305 7191 24363 7197
rect 24305 7157 24317 7191
rect 24351 7157 24363 7191
rect 24486 7188 24492 7200
rect 24447 7160 24492 7188
rect 24305 7151 24363 7157
rect 24486 7148 24492 7160
rect 24544 7148 24550 7200
rect 24670 7148 24676 7200
rect 24728 7188 24734 7200
rect 25332 7188 25360 7228
rect 26234 7216 26240 7268
rect 26292 7256 26298 7268
rect 29914 7256 29920 7268
rect 26292 7228 29920 7256
rect 26292 7216 26298 7228
rect 29914 7216 29920 7228
rect 29972 7216 29978 7268
rect 30374 7216 30380 7268
rect 30432 7256 30438 7268
rect 32493 7259 32551 7265
rect 32493 7256 32505 7259
rect 30432 7228 32505 7256
rect 30432 7216 30438 7228
rect 32493 7225 32505 7228
rect 32539 7225 32551 7259
rect 37090 7256 37096 7268
rect 32493 7219 32551 7225
rect 35452 7228 37096 7256
rect 24728 7160 25360 7188
rect 24728 7148 24734 7160
rect 25406 7148 25412 7200
rect 25464 7188 25470 7200
rect 25869 7191 25927 7197
rect 25869 7188 25881 7191
rect 25464 7160 25881 7188
rect 25464 7148 25470 7160
rect 25869 7157 25881 7160
rect 25915 7188 25927 7191
rect 27798 7188 27804 7200
rect 25915 7160 27804 7188
rect 25915 7157 25927 7160
rect 25869 7151 25927 7157
rect 27798 7148 27804 7160
rect 27856 7148 27862 7200
rect 27890 7148 27896 7200
rect 27948 7188 27954 7200
rect 27985 7191 28043 7197
rect 27985 7188 27997 7191
rect 27948 7160 27997 7188
rect 27948 7148 27954 7160
rect 27985 7157 27997 7160
rect 28031 7157 28043 7191
rect 28166 7188 28172 7200
rect 28127 7160 28172 7188
rect 27985 7151 28043 7157
rect 28166 7148 28172 7160
rect 28224 7148 28230 7200
rect 28718 7148 28724 7200
rect 28776 7188 28782 7200
rect 28905 7191 28963 7197
rect 28905 7188 28917 7191
rect 28776 7160 28917 7188
rect 28776 7148 28782 7160
rect 28905 7157 28917 7160
rect 28951 7157 28963 7191
rect 29086 7188 29092 7200
rect 29047 7160 29092 7188
rect 28905 7151 28963 7157
rect 29086 7148 29092 7160
rect 29144 7148 29150 7200
rect 29178 7148 29184 7200
rect 29236 7188 29242 7200
rect 35452 7188 35480 7228
rect 37090 7216 37096 7228
rect 37148 7216 37154 7268
rect 35618 7188 35624 7200
rect 29236 7160 35480 7188
rect 35579 7160 35624 7188
rect 29236 7148 29242 7160
rect 35618 7148 35624 7160
rect 35676 7148 35682 7200
rect 37200 7188 37228 7296
rect 37734 7284 37740 7296
rect 37792 7284 37798 7336
rect 42426 7284 42432 7336
rect 42484 7324 42490 7336
rect 43073 7327 43131 7333
rect 43073 7324 43085 7327
rect 42484 7296 43085 7324
rect 42484 7284 42490 7296
rect 43073 7293 43085 7296
rect 43119 7293 43131 7327
rect 44376 7324 44404 7355
rect 44542 7352 44548 7364
rect 44600 7352 44606 7404
rect 44634 7352 44640 7404
rect 44692 7392 44698 7404
rect 44775 7395 44833 7401
rect 44692 7364 44737 7392
rect 44692 7352 44698 7364
rect 44775 7361 44787 7395
rect 44821 7392 44833 7395
rect 45922 7392 45928 7404
rect 44821 7364 45928 7392
rect 44821 7361 44833 7364
rect 44775 7355 44833 7361
rect 45922 7352 45928 7364
rect 45980 7352 45986 7404
rect 46014 7352 46020 7404
rect 46072 7392 46078 7404
rect 46400 7401 46428 7500
rect 54846 7488 54852 7500
rect 54904 7488 54910 7540
rect 49145 7463 49203 7469
rect 49145 7429 49157 7463
rect 49191 7460 49203 7463
rect 50310 7463 50368 7469
rect 50310 7460 50322 7463
rect 49191 7432 50322 7460
rect 49191 7429 49203 7432
rect 49145 7423 49203 7429
rect 50310 7429 50322 7432
rect 50356 7429 50368 7463
rect 50310 7423 50368 7429
rect 52546 7420 52552 7472
rect 52604 7460 52610 7472
rect 53714 7463 53772 7469
rect 53714 7460 53726 7463
rect 52604 7432 53726 7460
rect 52604 7420 52610 7432
rect 53714 7429 53726 7432
rect 53760 7429 53772 7463
rect 53714 7423 53772 7429
rect 46293 7395 46351 7401
rect 46072 7364 46165 7392
rect 46072 7352 46078 7364
rect 46293 7361 46305 7395
rect 46339 7361 46351 7395
rect 46293 7355 46351 7361
rect 46385 7395 46443 7401
rect 46385 7361 46397 7395
rect 46431 7361 46443 7395
rect 46385 7355 46443 7361
rect 46032 7324 46060 7352
rect 44376 7296 46060 7324
rect 43073 7287 43131 7293
rect 46308 7256 46336 7355
rect 48774 7352 48780 7404
rect 48832 7392 48838 7404
rect 49326 7392 49332 7404
rect 48832 7364 49332 7392
rect 48832 7352 48838 7364
rect 49326 7352 49332 7364
rect 49384 7352 49390 7404
rect 49418 7352 49424 7404
rect 49476 7392 49482 7404
rect 49513 7395 49571 7401
rect 49513 7392 49525 7395
rect 49476 7364 49525 7392
rect 49476 7352 49482 7364
rect 49513 7361 49525 7364
rect 49559 7361 49571 7395
rect 51534 7392 51540 7404
rect 49513 7355 49571 7361
rect 50080 7364 51540 7392
rect 49602 7324 49608 7336
rect 49563 7296 49608 7324
rect 49602 7284 49608 7296
rect 49660 7284 49666 7336
rect 49878 7284 49884 7336
rect 49936 7324 49942 7336
rect 50080 7333 50108 7364
rect 51534 7352 51540 7364
rect 51592 7392 51598 7404
rect 53098 7392 53104 7404
rect 51592 7364 53104 7392
rect 51592 7352 51598 7364
rect 53098 7352 53104 7364
rect 53156 7392 53162 7404
rect 53469 7395 53527 7401
rect 53469 7392 53481 7395
rect 53156 7364 53481 7392
rect 53156 7352 53162 7364
rect 53469 7361 53481 7364
rect 53515 7361 53527 7395
rect 53469 7355 53527 7361
rect 50065 7327 50123 7333
rect 50065 7324 50077 7327
rect 49936 7296 50077 7324
rect 49936 7284 49942 7296
rect 50065 7293 50077 7296
rect 50111 7293 50123 7327
rect 50065 7287 50123 7293
rect 38672 7228 46336 7256
rect 38672 7188 38700 7228
rect 39114 7188 39120 7200
rect 37200 7160 38700 7188
rect 39075 7160 39120 7188
rect 39114 7148 39120 7160
rect 39172 7148 39178 7200
rect 42429 7191 42487 7197
rect 42429 7157 42441 7191
rect 42475 7188 42487 7191
rect 43070 7188 43076 7200
rect 42475 7160 43076 7188
rect 42475 7157 42487 7160
rect 42429 7151 42487 7157
rect 43070 7148 43076 7160
rect 43128 7148 43134 7200
rect 44913 7191 44971 7197
rect 44913 7157 44925 7191
rect 44959 7188 44971 7191
rect 45278 7188 45284 7200
rect 44959 7160 45284 7188
rect 44959 7157 44971 7160
rect 44913 7151 44971 7157
rect 45278 7148 45284 7160
rect 45336 7148 45342 7200
rect 46569 7191 46627 7197
rect 46569 7157 46581 7191
rect 46615 7188 46627 7191
rect 47210 7188 47216 7200
rect 46615 7160 47216 7188
rect 46615 7157 46627 7160
rect 46569 7151 46627 7157
rect 47210 7148 47216 7160
rect 47268 7148 47274 7200
rect 51445 7191 51503 7197
rect 51445 7157 51457 7191
rect 51491 7188 51503 7191
rect 51534 7188 51540 7200
rect 51491 7160 51540 7188
rect 51491 7157 51503 7160
rect 51445 7151 51503 7157
rect 51534 7148 51540 7160
rect 51592 7148 51598 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 14182 6984 14188 6996
rect 1636 6956 14188 6984
rect 1636 6944 1642 6956
rect 14182 6944 14188 6956
rect 14240 6944 14246 6996
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17184 6956 17264 6984
rect 17184 6944 17190 6956
rect 5644 6888 6500 6916
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 5644 6848 5672 6888
rect 1719 6820 5672 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 6472 6848 6500 6888
rect 15194 6876 15200 6928
rect 15252 6916 15258 6928
rect 15252 6888 17172 6916
rect 15252 6876 15258 6888
rect 11882 6848 11888 6860
rect 5776 6820 6408 6848
rect 6472 6820 11888 6848
rect 5776 6808 5782 6820
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 2866 6780 2872 6792
rect 2827 6752 2872 6780
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6270 6780 6276 6792
rect 6231 6752 6276 6780
rect 6089 6743 6147 6749
rect 3510 6672 3516 6724
rect 3568 6712 3574 6724
rect 6104 6712 6132 6743
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6380 6789 6408 6820
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 15102 6848 15108 6860
rect 14568 6820 15108 6848
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 8168 6752 9413 6780
rect 8168 6740 8174 6752
rect 9401 6749 9413 6752
rect 9447 6780 9459 6783
rect 9582 6780 9588 6792
rect 9447 6752 9588 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6780 14335 6783
rect 14458 6780 14464 6792
rect 14323 6752 14464 6780
rect 14323 6749 14335 6752
rect 14277 6743 14335 6749
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 14568 6789 14596 6820
rect 15102 6808 15108 6820
rect 15160 6808 15166 6860
rect 15654 6848 15660 6860
rect 15615 6820 15660 6848
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 17144 6857 17172 6888
rect 17236 6857 17264 6956
rect 19702 6944 19708 6996
rect 19760 6984 19766 6996
rect 19760 6956 23244 6984
rect 19760 6944 19766 6956
rect 23216 6928 23244 6956
rect 23382 6944 23388 6996
rect 23440 6984 23446 6996
rect 23477 6987 23535 6993
rect 23477 6984 23489 6987
rect 23440 6956 23489 6984
rect 23440 6944 23446 6956
rect 23477 6953 23489 6956
rect 23523 6953 23535 6987
rect 23477 6947 23535 6953
rect 23750 6944 23756 6996
rect 23808 6984 23814 6996
rect 27798 6984 27804 6996
rect 23808 6956 27804 6984
rect 23808 6944 23814 6956
rect 27798 6944 27804 6956
rect 27856 6944 27862 6996
rect 27890 6944 27896 6996
rect 27948 6984 27954 6996
rect 27985 6987 28043 6993
rect 27985 6984 27997 6987
rect 27948 6956 27997 6984
rect 27948 6944 27954 6956
rect 27985 6953 27997 6956
rect 28031 6953 28043 6987
rect 34514 6984 34520 6996
rect 27985 6947 28043 6953
rect 28092 6956 34520 6984
rect 19426 6876 19432 6928
rect 19484 6916 19490 6928
rect 21726 6916 21732 6928
rect 19484 6888 21732 6916
rect 19484 6876 19490 6888
rect 21726 6876 21732 6888
rect 21784 6876 21790 6928
rect 23198 6876 23204 6928
rect 23256 6916 23262 6928
rect 28092 6916 28120 6956
rect 34514 6944 34520 6956
rect 34572 6944 34578 6996
rect 34790 6944 34796 6996
rect 34848 6984 34854 6996
rect 35802 6984 35808 6996
rect 34848 6956 35808 6984
rect 34848 6944 34854 6956
rect 35802 6944 35808 6956
rect 35860 6944 35866 6996
rect 37458 6984 37464 6996
rect 37419 6956 37464 6984
rect 37458 6944 37464 6956
rect 37516 6944 37522 6996
rect 37734 6944 37740 6996
rect 37792 6984 37798 6996
rect 40034 6984 40040 6996
rect 37792 6956 40040 6984
rect 37792 6944 37798 6956
rect 40034 6944 40040 6956
rect 40092 6944 40098 6996
rect 45370 6984 45376 6996
rect 44284 6956 45376 6984
rect 30650 6916 30656 6928
rect 23256 6888 28120 6916
rect 28966 6888 30656 6916
rect 23256 6876 23262 6888
rect 17129 6851 17187 6857
rect 17129 6817 17141 6851
rect 17175 6817 17187 6851
rect 17129 6811 17187 6817
rect 17221 6851 17279 6857
rect 17221 6817 17233 6851
rect 17267 6817 17279 6851
rect 17402 6848 17408 6860
rect 17363 6820 17408 6848
rect 17221 6811 17279 6817
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 17494 6808 17500 6860
rect 17552 6848 17558 6860
rect 17552 6820 19840 6848
rect 17552 6808 17558 6820
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 15930 6780 15936 6792
rect 15891 6752 15936 6780
rect 14553 6743 14611 6749
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 19426 6780 19432 6792
rect 17368 6752 17413 6780
rect 19387 6752 19432 6780
rect 17368 6740 17374 6752
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 19702 6780 19708 6792
rect 19615 6752 19708 6780
rect 19702 6740 19708 6752
rect 19760 6740 19766 6792
rect 9122 6712 9128 6724
rect 3568 6684 6040 6712
rect 6104 6684 9128 6712
rect 3568 6672 3574 6684
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 2685 6647 2743 6653
rect 2685 6644 2697 6647
rect 2648 6616 2697 6644
rect 2648 6604 2654 6616
rect 2685 6613 2697 6616
rect 2731 6613 2743 6647
rect 5902 6644 5908 6656
rect 5863 6616 5908 6644
rect 2685 6607 2743 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6012 6644 6040 6684
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 19150 6672 19156 6724
rect 19208 6712 19214 6724
rect 19613 6715 19671 6721
rect 19613 6712 19625 6715
rect 19208 6684 19625 6712
rect 19208 6672 19214 6684
rect 19613 6681 19625 6684
rect 19659 6681 19671 6715
rect 19613 6675 19671 6681
rect 7466 6644 7472 6656
rect 6012 6616 7472 6644
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 11146 6644 11152 6656
rect 10284 6616 11152 6644
rect 10284 6604 10290 6616
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 14090 6644 14096 6656
rect 14051 6616 14096 6644
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14458 6644 14464 6656
rect 14419 6616 14464 6644
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 15378 6604 15384 6656
rect 15436 6644 15442 6656
rect 16945 6647 17003 6653
rect 16945 6644 16957 6647
rect 15436 6616 16957 6644
rect 15436 6604 15442 6616
rect 16945 6613 16957 6616
rect 16991 6613 17003 6647
rect 19242 6644 19248 6656
rect 19203 6616 19248 6644
rect 16945 6607 17003 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 19720 6644 19748 6740
rect 19812 6712 19840 6820
rect 25222 6808 25228 6860
rect 25280 6848 25286 6860
rect 26142 6848 26148 6860
rect 25280 6820 26148 6848
rect 25280 6808 25286 6820
rect 26142 6808 26148 6820
rect 26200 6808 26206 6860
rect 26326 6808 26332 6860
rect 26384 6848 26390 6860
rect 28966 6848 28994 6888
rect 30650 6876 30656 6888
rect 30708 6876 30714 6928
rect 31110 6876 31116 6928
rect 31168 6916 31174 6928
rect 31168 6888 32628 6916
rect 31168 6876 31174 6888
rect 26384 6820 28994 6848
rect 26384 6808 26390 6820
rect 30190 6808 30196 6860
rect 30248 6848 30254 6860
rect 32490 6848 32496 6860
rect 30248 6820 32496 6848
rect 30248 6808 30254 6820
rect 20622 6740 20628 6792
rect 20680 6780 20686 6792
rect 22097 6783 22155 6789
rect 22097 6780 22109 6783
rect 20680 6752 22109 6780
rect 20680 6740 20686 6752
rect 22097 6749 22109 6752
rect 22143 6749 22155 6783
rect 22097 6743 22155 6749
rect 22364 6783 22422 6789
rect 22364 6749 22376 6783
rect 22410 6780 22422 6783
rect 22738 6780 22744 6792
rect 22410 6752 22744 6780
rect 22410 6749 22422 6752
rect 22364 6743 22422 6749
rect 22738 6740 22744 6752
rect 22796 6740 22802 6792
rect 30484 6789 30512 6820
rect 32490 6808 32496 6820
rect 32548 6808 32554 6860
rect 32600 6848 32628 6888
rect 33410 6848 33416 6860
rect 32600 6820 33416 6848
rect 33410 6808 33416 6820
rect 33468 6808 33474 6860
rect 37093 6851 37151 6857
rect 37093 6817 37105 6851
rect 37139 6848 37151 6851
rect 37182 6848 37188 6860
rect 37139 6820 37188 6848
rect 37139 6817 37151 6820
rect 37093 6811 37151 6817
rect 37182 6808 37188 6820
rect 37240 6808 37246 6860
rect 37366 6848 37372 6860
rect 37292 6820 37372 6848
rect 30469 6783 30527 6789
rect 24780 6752 27844 6780
rect 24780 6712 24808 6752
rect 19812 6684 24808 6712
rect 24857 6715 24915 6721
rect 24857 6681 24869 6715
rect 24903 6712 24915 6715
rect 25590 6712 25596 6724
rect 24903 6684 25596 6712
rect 24903 6681 24915 6684
rect 24857 6675 24915 6681
rect 25590 6672 25596 6684
rect 25648 6672 25654 6724
rect 27816 6721 27844 6752
rect 30469 6749 30481 6783
rect 30515 6749 30527 6783
rect 32306 6780 32312 6792
rect 32267 6752 32312 6780
rect 30469 6743 30527 6749
rect 32306 6740 32312 6752
rect 32364 6740 32370 6792
rect 32585 6783 32643 6789
rect 32585 6780 32597 6783
rect 32416 6752 32597 6780
rect 27801 6715 27859 6721
rect 27801 6681 27813 6715
rect 27847 6681 27859 6715
rect 27801 6675 27859 6681
rect 28184 6684 30788 6712
rect 19392 6616 19748 6644
rect 19392 6604 19398 6616
rect 22830 6604 22836 6656
rect 22888 6644 22894 6656
rect 24949 6647 25007 6653
rect 24949 6644 24961 6647
rect 22888 6616 24961 6644
rect 22888 6604 22894 6616
rect 24949 6613 24961 6616
rect 24995 6644 25007 6647
rect 26418 6644 26424 6656
rect 24995 6616 26424 6644
rect 24995 6613 25007 6616
rect 24949 6607 25007 6613
rect 26418 6604 26424 6616
rect 26476 6644 26482 6656
rect 27522 6644 27528 6656
rect 26476 6616 27528 6644
rect 26476 6604 26482 6616
rect 27522 6604 27528 6616
rect 27580 6604 27586 6656
rect 27982 6604 27988 6656
rect 28040 6653 28046 6656
rect 28184 6653 28212 6684
rect 28040 6647 28059 6653
rect 28047 6613 28059 6647
rect 28040 6607 28059 6613
rect 28169 6647 28227 6653
rect 28169 6613 28181 6647
rect 28215 6613 28227 6647
rect 30760 6644 30788 6684
rect 30834 6672 30840 6724
rect 30892 6712 30898 6724
rect 32416 6712 32444 6752
rect 32585 6749 32597 6752
rect 32631 6749 32643 6783
rect 32585 6743 32643 6749
rect 32677 6783 32735 6789
rect 32677 6749 32689 6783
rect 32723 6780 32735 6783
rect 33318 6780 33324 6792
rect 32723 6752 33324 6780
rect 32723 6749 32735 6752
rect 32677 6743 32735 6749
rect 33318 6740 33324 6752
rect 33376 6740 33382 6792
rect 34698 6740 34704 6792
rect 34756 6780 34762 6792
rect 34793 6783 34851 6789
rect 34793 6780 34805 6783
rect 34756 6752 34805 6780
rect 34756 6740 34762 6752
rect 34793 6749 34805 6752
rect 34839 6749 34851 6783
rect 34793 6743 34851 6749
rect 35060 6783 35118 6789
rect 35060 6749 35072 6783
rect 35106 6780 35118 6783
rect 35618 6780 35624 6792
rect 35106 6752 35624 6780
rect 35106 6749 35118 6752
rect 35060 6743 35118 6749
rect 35618 6740 35624 6752
rect 35676 6740 35682 6792
rect 36538 6740 36544 6792
rect 36596 6780 36602 6792
rect 36725 6783 36783 6789
rect 36725 6780 36737 6783
rect 36596 6752 36737 6780
rect 36596 6740 36602 6752
rect 36725 6749 36737 6752
rect 36771 6749 36783 6783
rect 36906 6780 36912 6792
rect 36867 6752 36912 6780
rect 36725 6743 36783 6749
rect 36906 6740 36912 6752
rect 36964 6740 36970 6792
rect 37292 6789 37320 6820
rect 37366 6808 37372 6820
rect 37424 6808 37430 6860
rect 37458 6808 37464 6860
rect 37516 6848 37522 6860
rect 44174 6848 44180 6860
rect 37516 6820 44180 6848
rect 37516 6808 37522 6820
rect 44174 6808 44180 6820
rect 44232 6808 44238 6860
rect 37001 6783 37059 6789
rect 37001 6749 37013 6783
rect 37047 6749 37059 6783
rect 37001 6743 37059 6749
rect 37277 6783 37335 6789
rect 37277 6749 37289 6783
rect 37323 6749 37335 6783
rect 44284 6780 44312 6956
rect 45370 6944 45376 6956
rect 45428 6944 45434 6996
rect 45005 6851 45063 6857
rect 45005 6817 45017 6851
rect 45051 6817 45063 6851
rect 51534 6848 51540 6860
rect 45005 6811 45063 6817
rect 48884 6820 51540 6848
rect 37277 6743 37335 6749
rect 40604 6752 44312 6780
rect 45020 6780 45048 6811
rect 48884 6792 48912 6820
rect 51534 6808 51540 6820
rect 51592 6808 51598 6860
rect 52730 6848 52736 6860
rect 52656 6820 52736 6848
rect 46934 6780 46940 6792
rect 45020 6752 46940 6780
rect 30892 6684 32444 6712
rect 30892 6672 30898 6684
rect 32490 6672 32496 6724
rect 32548 6712 32554 6724
rect 32548 6684 32593 6712
rect 32692 6684 36308 6712
rect 32548 6672 32554 6684
rect 32692 6644 32720 6684
rect 32858 6644 32864 6656
rect 30760 6616 32720 6644
rect 32819 6616 32864 6644
rect 28169 6607 28227 6613
rect 28040 6604 28046 6607
rect 32858 6604 32864 6616
rect 32916 6604 32922 6656
rect 36170 6644 36176 6656
rect 36131 6616 36176 6644
rect 36170 6604 36176 6616
rect 36228 6604 36234 6656
rect 36280 6644 36308 6684
rect 36814 6672 36820 6724
rect 36872 6712 36878 6724
rect 37016 6712 37044 6743
rect 40604 6712 40632 6752
rect 46934 6740 46940 6752
rect 46992 6780 46998 6792
rect 47118 6780 47124 6792
rect 46992 6752 47124 6780
rect 46992 6740 46998 6752
rect 47118 6740 47124 6752
rect 47176 6740 47182 6792
rect 47210 6740 47216 6792
rect 47268 6780 47274 6792
rect 47377 6783 47435 6789
rect 47377 6780 47389 6783
rect 47268 6752 47389 6780
rect 47268 6740 47274 6752
rect 47377 6749 47389 6752
rect 47423 6749 47435 6783
rect 47377 6743 47435 6749
rect 48222 6740 48228 6792
rect 48280 6780 48286 6792
rect 48866 6780 48872 6792
rect 48280 6752 48872 6780
rect 48280 6740 48286 6752
rect 48866 6740 48872 6752
rect 48924 6740 48930 6792
rect 49326 6780 49332 6792
rect 49287 6752 49332 6780
rect 49326 6740 49332 6752
rect 49384 6740 49390 6792
rect 49513 6783 49571 6789
rect 49513 6749 49525 6783
rect 49559 6749 49571 6783
rect 49513 6743 49571 6749
rect 49605 6783 49663 6789
rect 49605 6749 49617 6783
rect 49651 6780 49663 6783
rect 50154 6780 50160 6792
rect 49651 6752 50160 6780
rect 49651 6749 49663 6752
rect 49605 6743 49663 6749
rect 36872 6684 37044 6712
rect 37108 6684 40632 6712
rect 36872 6672 36878 6684
rect 37108 6644 37136 6684
rect 40678 6672 40684 6724
rect 40736 6712 40742 6724
rect 45278 6721 45284 6724
rect 41325 6715 41383 6721
rect 41325 6712 41337 6715
rect 40736 6684 41337 6712
rect 40736 6672 40742 6684
rect 41325 6681 41337 6684
rect 41371 6681 41383 6715
rect 45272 6712 45284 6721
rect 45239 6684 45284 6712
rect 41325 6675 41383 6681
rect 45272 6675 45284 6684
rect 45278 6672 45284 6675
rect 45336 6672 45342 6724
rect 45370 6672 45376 6724
rect 45428 6712 45434 6724
rect 49528 6712 49556 6743
rect 50154 6740 50160 6752
rect 50212 6740 50218 6792
rect 52656 6789 52684 6820
rect 52730 6808 52736 6820
rect 52788 6808 52794 6860
rect 52641 6783 52699 6789
rect 52641 6749 52653 6783
rect 52687 6749 52699 6783
rect 52641 6743 52699 6749
rect 52825 6783 52883 6789
rect 52825 6749 52837 6783
rect 52871 6749 52883 6783
rect 52825 6743 52883 6749
rect 45428 6684 49556 6712
rect 45428 6672 45434 6684
rect 50062 6672 50068 6724
rect 50120 6712 50126 6724
rect 52840 6712 52868 6743
rect 52914 6740 52920 6792
rect 52972 6780 52978 6792
rect 52972 6752 53017 6780
rect 52972 6740 52978 6752
rect 50120 6684 52868 6712
rect 50120 6672 50126 6684
rect 36280 6616 37136 6644
rect 37366 6604 37372 6656
rect 37424 6644 37430 6656
rect 39114 6644 39120 6656
rect 37424 6616 39120 6644
rect 37424 6604 37430 6616
rect 39114 6604 39120 6616
rect 39172 6604 39178 6656
rect 41414 6604 41420 6656
rect 41472 6644 41478 6656
rect 41472 6616 41517 6644
rect 41472 6604 41478 6616
rect 45922 6604 45928 6656
rect 45980 6644 45986 6656
rect 46385 6647 46443 6653
rect 46385 6644 46397 6647
rect 45980 6616 46397 6644
rect 45980 6604 45986 6616
rect 46385 6613 46397 6616
rect 46431 6613 46443 6647
rect 46385 6607 46443 6613
rect 48406 6604 48412 6656
rect 48464 6644 48470 6656
rect 48501 6647 48559 6653
rect 48501 6644 48513 6647
rect 48464 6616 48513 6644
rect 48464 6604 48470 6616
rect 48501 6613 48513 6616
rect 48547 6613 48559 6647
rect 48501 6607 48559 6613
rect 49145 6647 49203 6653
rect 49145 6613 49157 6647
rect 49191 6644 49203 6647
rect 49694 6644 49700 6656
rect 49191 6616 49700 6644
rect 49191 6613 49203 6616
rect 49145 6607 49203 6613
rect 49694 6604 49700 6616
rect 49752 6604 49758 6656
rect 52457 6647 52515 6653
rect 52457 6613 52469 6647
rect 52503 6644 52515 6647
rect 53282 6644 53288 6656
rect 52503 6616 53288 6644
rect 52503 6613 52515 6616
rect 52457 6607 52515 6613
rect 53282 6604 53288 6616
rect 53340 6604 53346 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 2593 6443 2651 6449
rect 2593 6409 2605 6443
rect 2639 6440 2651 6443
rect 3326 6440 3332 6452
rect 2639 6412 3332 6440
rect 2639 6409 2651 6412
rect 2593 6403 2651 6409
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 15197 6443 15255 6449
rect 15197 6440 15209 6443
rect 5000 6412 15209 6440
rect 3510 6372 3516 6384
rect 2516 6344 3516 6372
rect 2516 6313 2544 6344
rect 3510 6332 3516 6344
rect 3568 6332 3574 6384
rect 5000 6313 5028 6412
rect 15197 6409 15209 6412
rect 15243 6409 15255 6443
rect 15197 6403 15255 6409
rect 15654 6400 15660 6452
rect 15712 6400 15718 6452
rect 17310 6400 17316 6452
rect 17368 6440 17374 6452
rect 23382 6440 23388 6452
rect 17368 6412 23388 6440
rect 17368 6400 17374 6412
rect 23382 6400 23388 6412
rect 23440 6400 23446 6452
rect 24578 6400 24584 6452
rect 24636 6440 24642 6452
rect 32674 6440 32680 6452
rect 24636 6412 32680 6440
rect 24636 6400 24642 6412
rect 32674 6400 32680 6412
rect 32732 6400 32738 6452
rect 33505 6443 33563 6449
rect 33505 6409 33517 6443
rect 33551 6440 33563 6443
rect 33594 6440 33600 6452
rect 33551 6412 33600 6440
rect 33551 6409 33563 6412
rect 33505 6403 33563 6409
rect 33594 6400 33600 6412
rect 33652 6400 33658 6452
rect 36633 6443 36691 6449
rect 36633 6409 36645 6443
rect 36679 6440 36691 6443
rect 36814 6440 36820 6452
rect 36679 6412 36820 6440
rect 36679 6409 36691 6412
rect 36633 6403 36691 6409
rect 36814 6400 36820 6412
rect 36872 6400 36878 6452
rect 38286 6400 38292 6452
rect 38344 6440 38350 6452
rect 44542 6440 44548 6452
rect 38344 6412 41414 6440
rect 44503 6412 44548 6440
rect 38344 6400 38350 6412
rect 5902 6332 5908 6384
rect 5960 6372 5966 6384
rect 6610 6375 6668 6381
rect 6610 6372 6622 6375
rect 5960 6344 6622 6372
rect 5960 6332 5966 6344
rect 6610 6341 6622 6344
rect 6656 6341 6668 6375
rect 6610 6335 6668 6341
rect 13348 6375 13406 6381
rect 13348 6341 13360 6375
rect 13394 6372 13406 6375
rect 14090 6372 14096 6384
rect 13394 6344 14096 6372
rect 13394 6341 13406 6344
rect 13348 6335 13406 6341
rect 14090 6332 14096 6344
rect 14148 6332 14154 6384
rect 15672 6372 15700 6400
rect 18500 6375 18558 6381
rect 15488 6344 15700 6372
rect 15856 6344 17172 6372
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6304 5319 6307
rect 5718 6304 5724 6316
rect 5307 6276 5724 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 1412 6168 1440 6267
rect 2682 6196 2688 6248
rect 2740 6236 2746 6248
rect 2740 6208 2785 6236
rect 2740 6196 2746 6208
rect 5184 6168 5212 6267
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6304 8907 6307
rect 10410 6304 10416 6316
rect 8895 6276 10416 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 10410 6264 10416 6276
rect 10468 6264 10474 6316
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 11020 6276 13093 6304
rect 11020 6264 11026 6276
rect 13081 6273 13093 6276
rect 13127 6304 13139 6307
rect 13814 6304 13820 6316
rect 13127 6276 13820 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 15378 6304 15384 6316
rect 15339 6276 15384 6304
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 15488 6313 15516 6344
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6273 15531 6307
rect 15473 6267 15531 6273
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6304 15715 6307
rect 15746 6304 15752 6316
rect 15703 6276 15752 6304
rect 15703 6273 15715 6276
rect 15657 6267 15715 6273
rect 15746 6264 15752 6276
rect 15804 6304 15810 6316
rect 15856 6304 15884 6344
rect 15804 6276 15884 6304
rect 15804 6264 15810 6276
rect 15930 6264 15936 6316
rect 15988 6304 15994 6316
rect 17144 6313 17172 6344
rect 18500 6341 18512 6375
rect 18546 6372 18558 6375
rect 19242 6372 19248 6384
rect 18546 6344 19248 6372
rect 18546 6341 18558 6344
rect 18500 6335 18558 6341
rect 19242 6332 19248 6344
rect 19300 6332 19306 6384
rect 22094 6332 22100 6384
rect 22152 6372 22158 6384
rect 22465 6375 22523 6381
rect 22465 6372 22477 6375
rect 22152 6344 22477 6372
rect 22152 6332 22158 6344
rect 22465 6341 22477 6344
rect 22511 6341 22523 6375
rect 22465 6335 22523 6341
rect 22554 6332 22560 6384
rect 22612 6332 22618 6384
rect 22649 6375 22707 6381
rect 22649 6341 22661 6375
rect 22695 6372 22707 6375
rect 28350 6372 28356 6384
rect 22695 6344 28356 6372
rect 22695 6341 22707 6344
rect 22649 6335 22707 6341
rect 28350 6332 28356 6344
rect 28408 6332 28414 6384
rect 29454 6372 29460 6384
rect 29415 6344 29460 6372
rect 29454 6332 29460 6344
rect 29512 6332 29518 6384
rect 29673 6375 29731 6381
rect 29673 6341 29685 6375
rect 29719 6372 29731 6375
rect 31294 6372 31300 6384
rect 29719 6344 31300 6372
rect 29719 6341 29731 6344
rect 29673 6335 29731 6341
rect 31294 6332 31300 6344
rect 31352 6332 31358 6384
rect 32392 6375 32450 6381
rect 32392 6341 32404 6375
rect 32438 6372 32450 6375
rect 32858 6372 32864 6384
rect 32438 6344 32864 6372
rect 32438 6341 32450 6344
rect 32392 6335 32450 6341
rect 32858 6332 32864 6344
rect 32916 6332 32922 6384
rect 41386 6372 41414 6412
rect 44542 6400 44548 6412
rect 44600 6400 44606 6452
rect 46198 6400 46204 6452
rect 46256 6440 46262 6452
rect 46753 6443 46811 6449
rect 46753 6440 46765 6443
rect 46256 6412 46765 6440
rect 46256 6400 46262 6412
rect 46753 6409 46765 6412
rect 46799 6409 46811 6443
rect 46753 6403 46811 6409
rect 46842 6400 46848 6452
rect 46900 6440 46906 6452
rect 49145 6443 49203 6449
rect 46900 6412 49096 6440
rect 46900 6400 46906 6412
rect 44174 6372 44180 6384
rect 33244 6344 40172 6372
rect 41386 6344 43852 6372
rect 44135 6344 44180 6372
rect 17037 6307 17095 6313
rect 17037 6304 17049 6307
rect 15988 6276 17049 6304
rect 15988 6264 15994 6276
rect 17037 6273 17049 6276
rect 17083 6273 17095 6307
rect 17037 6267 17095 6273
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6273 17187 6307
rect 17129 6267 17187 6273
rect 18138 6264 18144 6316
rect 18196 6304 18202 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 18196 6276 18245 6304
rect 18196 6264 18202 6276
rect 18233 6273 18245 6276
rect 18279 6304 18291 6307
rect 20622 6304 20628 6316
rect 18279 6276 20628 6304
rect 18279 6273 18291 6276
rect 18233 6267 18291 6273
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 21358 6264 21364 6316
rect 21416 6304 21422 6316
rect 22278 6304 22284 6316
rect 21416 6276 22284 6304
rect 21416 6264 21422 6276
rect 22278 6264 22284 6276
rect 22336 6264 22342 6316
rect 22373 6307 22431 6313
rect 22373 6273 22385 6307
rect 22419 6304 22431 6307
rect 22572 6304 22600 6332
rect 22419 6276 22600 6304
rect 22419 6273 22431 6276
rect 22373 6267 22431 6273
rect 25682 6264 25688 6316
rect 25740 6304 25746 6316
rect 33244 6304 33272 6344
rect 25740 6276 33272 6304
rect 25740 6264 25746 6276
rect 36262 6264 36268 6316
rect 36320 6304 36326 6316
rect 36449 6307 36507 6313
rect 36320 6276 36365 6304
rect 36320 6264 36326 6276
rect 36449 6273 36461 6307
rect 36495 6273 36507 6307
rect 36449 6267 36507 6273
rect 39945 6307 40003 6313
rect 39945 6273 39957 6307
rect 39991 6304 40003 6307
rect 40034 6304 40040 6316
rect 39991 6276 40040 6304
rect 39991 6273 40003 6276
rect 39945 6267 40003 6273
rect 5350 6196 5356 6248
rect 5408 6236 5414 6248
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5408 6208 6377 6236
rect 5408 6196 5414 6208
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 6365 6199 6423 6205
rect 8864 6208 9137 6236
rect 8864 6180 8892 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 15562 6236 15568 6248
rect 15523 6208 15568 6236
rect 9125 6199 9183 6205
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 16850 6236 16856 6248
rect 16811 6208 16856 6236
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 16942 6196 16948 6248
rect 17000 6236 17006 6248
rect 30834 6236 30840 6248
rect 17000 6208 17045 6236
rect 27724 6208 30840 6236
rect 17000 6196 17006 6208
rect 5442 6168 5448 6180
rect 1412 6140 5448 6168
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 8846 6128 8852 6180
rect 8904 6128 8910 6180
rect 9033 6171 9091 6177
rect 9033 6137 9045 6171
rect 9079 6168 9091 6171
rect 9214 6168 9220 6180
rect 9079 6140 9220 6168
rect 9079 6137 9091 6140
rect 9033 6131 9091 6137
rect 9214 6128 9220 6140
rect 9272 6128 9278 6180
rect 16669 6171 16727 6177
rect 16669 6168 16681 6171
rect 14384 6140 16681 6168
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2133 6103 2191 6109
rect 2133 6069 2145 6103
rect 2179 6100 2191 6103
rect 3602 6100 3608 6112
rect 2179 6072 3608 6100
rect 2179 6069 2191 6072
rect 2133 6063 2191 6069
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 4798 6100 4804 6112
rect 4759 6072 4804 6100
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 6328 6072 7757 6100
rect 6328 6060 6334 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 8665 6103 8723 6109
rect 8665 6069 8677 6103
rect 8711 6100 8723 6103
rect 8938 6100 8944 6112
rect 8711 6072 8944 6100
rect 8711 6069 8723 6072
rect 8665 6063 8723 6069
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 9122 6060 9128 6112
rect 9180 6100 9186 6112
rect 14384 6100 14412 6140
rect 16669 6137 16681 6140
rect 16715 6137 16727 6171
rect 16669 6131 16727 6137
rect 22097 6171 22155 6177
rect 22097 6137 22109 6171
rect 22143 6137 22155 6171
rect 22097 6131 22155 6137
rect 9180 6072 14412 6100
rect 9180 6060 9186 6072
rect 14458 6060 14464 6112
rect 14516 6100 14522 6112
rect 14516 6072 14561 6100
rect 14516 6060 14522 6072
rect 19150 6060 19156 6112
rect 19208 6100 19214 6112
rect 19613 6103 19671 6109
rect 19613 6100 19625 6103
rect 19208 6072 19625 6100
rect 19208 6060 19214 6072
rect 19613 6069 19625 6072
rect 19659 6069 19671 6103
rect 22112 6100 22140 6131
rect 23842 6128 23848 6180
rect 23900 6168 23906 6180
rect 27724 6168 27752 6208
rect 30834 6196 30840 6208
rect 30892 6196 30898 6248
rect 31846 6196 31852 6248
rect 31904 6236 31910 6248
rect 32125 6239 32183 6245
rect 32125 6236 32137 6239
rect 31904 6208 32137 6236
rect 31904 6196 31910 6208
rect 32125 6205 32137 6208
rect 32171 6205 32183 6239
rect 32125 6199 32183 6205
rect 36354 6196 36360 6248
rect 36412 6236 36418 6248
rect 36464 6236 36492 6267
rect 40034 6264 40040 6276
rect 40092 6264 40098 6316
rect 40144 6313 40172 6344
rect 40129 6307 40187 6313
rect 40129 6273 40141 6307
rect 40175 6273 40187 6307
rect 40129 6267 40187 6273
rect 41414 6264 41420 6316
rect 41472 6304 41478 6316
rect 42889 6307 42947 6313
rect 42889 6304 42901 6307
rect 41472 6276 42901 6304
rect 41472 6264 41478 6276
rect 42889 6273 42901 6276
rect 42935 6273 42947 6307
rect 43070 6304 43076 6316
rect 43031 6276 43076 6304
rect 42889 6267 42947 6273
rect 43070 6264 43076 6276
rect 43128 6264 43134 6316
rect 36412 6208 36492 6236
rect 36412 6196 36418 6208
rect 36630 6196 36636 6248
rect 36688 6236 36694 6248
rect 40221 6239 40279 6245
rect 36688 6208 40172 6236
rect 36688 6196 36694 6208
rect 23900 6140 27752 6168
rect 23900 6128 23906 6140
rect 28166 6128 28172 6180
rect 28224 6168 28230 6180
rect 39666 6168 39672 6180
rect 28224 6140 32168 6168
rect 28224 6128 28230 6140
rect 22278 6100 22284 6112
rect 22112 6072 22284 6100
rect 19613 6063 19671 6069
rect 22278 6060 22284 6072
rect 22336 6100 22342 6112
rect 24946 6100 24952 6112
rect 22336 6072 24952 6100
rect 22336 6060 22342 6072
rect 24946 6060 24952 6072
rect 25004 6060 25010 6112
rect 25774 6060 25780 6112
rect 25832 6100 25838 6112
rect 28718 6100 28724 6112
rect 25832 6072 28724 6100
rect 25832 6060 25838 6072
rect 28718 6060 28724 6072
rect 28776 6060 28782 6112
rect 28902 6060 28908 6112
rect 28960 6100 28966 6112
rect 29641 6103 29699 6109
rect 29641 6100 29653 6103
rect 28960 6072 29653 6100
rect 28960 6060 28966 6072
rect 29641 6069 29653 6072
rect 29687 6069 29699 6103
rect 29822 6100 29828 6112
rect 29783 6072 29828 6100
rect 29641 6063 29699 6069
rect 29822 6060 29828 6072
rect 29880 6060 29886 6112
rect 32140 6100 32168 6140
rect 33060 6140 39672 6168
rect 33060 6100 33088 6140
rect 39666 6128 39672 6140
rect 39724 6128 39730 6180
rect 40144 6168 40172 6208
rect 40221 6205 40233 6239
rect 40267 6236 40279 6239
rect 40586 6236 40592 6248
rect 40267 6208 40592 6236
rect 40267 6205 40279 6208
rect 40221 6199 40279 6205
rect 40586 6196 40592 6208
rect 40644 6196 40650 6248
rect 43162 6236 43168 6248
rect 43123 6208 43168 6236
rect 43162 6196 43168 6208
rect 43220 6196 43226 6248
rect 43824 6236 43852 6344
rect 44174 6332 44180 6344
rect 44232 6332 44238 6384
rect 44269 6375 44327 6381
rect 44269 6341 44281 6375
rect 44315 6372 44327 6375
rect 45922 6372 45928 6384
rect 44315 6344 45928 6372
rect 44315 6341 44327 6344
rect 44269 6335 44327 6341
rect 45922 6332 45928 6344
rect 45980 6332 45986 6384
rect 46385 6375 46443 6381
rect 46385 6372 46397 6375
rect 46124 6344 46397 6372
rect 43990 6304 43996 6316
rect 43951 6276 43996 6304
rect 43990 6264 43996 6276
rect 44048 6264 44054 6316
rect 44192 6236 44220 6332
rect 44358 6264 44364 6316
rect 44416 6304 44422 6316
rect 44416 6276 44461 6304
rect 44416 6264 44422 6276
rect 46124 6236 46152 6344
rect 46385 6341 46397 6344
rect 46431 6341 46443 6375
rect 46385 6335 46443 6341
rect 46477 6375 46535 6381
rect 46477 6341 46489 6375
rect 46523 6372 46535 6375
rect 48866 6372 48872 6384
rect 46523 6344 48314 6372
rect 48827 6344 48872 6372
rect 46523 6341 46535 6344
rect 46477 6335 46535 6341
rect 46201 6307 46259 6313
rect 46201 6273 46213 6307
rect 46247 6273 46259 6307
rect 46201 6267 46259 6273
rect 43824 6208 44128 6236
rect 44192 6208 46152 6236
rect 46216 6236 46244 6267
rect 46290 6264 46296 6316
rect 46348 6304 46354 6316
rect 46569 6307 46627 6313
rect 46569 6304 46581 6307
rect 46348 6276 46581 6304
rect 46348 6264 46354 6276
rect 46569 6273 46581 6276
rect 46615 6273 46627 6307
rect 48286 6304 48314 6344
rect 48866 6332 48872 6344
rect 48924 6332 48930 6384
rect 49068 6372 49096 6412
rect 49145 6409 49157 6443
rect 49191 6440 49203 6443
rect 49602 6440 49608 6452
rect 49191 6412 49608 6440
rect 49191 6409 49203 6412
rect 49145 6403 49203 6409
rect 49602 6400 49608 6412
rect 49660 6400 49666 6452
rect 50154 6440 50160 6452
rect 50115 6412 50160 6440
rect 50154 6400 50160 6412
rect 50212 6400 50218 6452
rect 53006 6400 53012 6452
rect 53064 6440 53070 6452
rect 53285 6443 53343 6449
rect 53285 6440 53297 6443
rect 53064 6412 53297 6440
rect 53064 6400 53070 6412
rect 53285 6409 53297 6412
rect 53331 6409 53343 6443
rect 53285 6403 53343 6409
rect 49881 6375 49939 6381
rect 49881 6372 49893 6375
rect 49068 6344 49893 6372
rect 49881 6341 49893 6344
rect 49927 6372 49939 6375
rect 50982 6372 50988 6384
rect 49927 6344 50988 6372
rect 49927 6341 49939 6344
rect 49881 6335 49939 6341
rect 50982 6332 50988 6344
rect 51040 6332 51046 6384
rect 52178 6332 52184 6384
rect 52236 6372 52242 6384
rect 52917 6375 52975 6381
rect 52917 6372 52929 6375
rect 52236 6344 52929 6372
rect 52236 6332 52242 6344
rect 52917 6341 52929 6344
rect 52963 6341 52975 6375
rect 54846 6372 54852 6384
rect 52917 6335 52975 6341
rect 53024 6344 54852 6372
rect 48406 6304 48412 6316
rect 48286 6276 48412 6304
rect 46569 6267 46627 6273
rect 48406 6264 48412 6276
rect 48464 6304 48470 6316
rect 48593 6307 48651 6313
rect 48593 6304 48605 6307
rect 48464 6276 48605 6304
rect 48464 6264 48470 6276
rect 48593 6273 48605 6276
rect 48639 6273 48651 6307
rect 48593 6267 48651 6273
rect 48774 6264 48780 6316
rect 48832 6304 48838 6316
rect 48961 6307 49019 6313
rect 48832 6276 48877 6304
rect 48832 6264 48838 6276
rect 48961 6273 48973 6307
rect 49007 6304 49019 6307
rect 49418 6304 49424 6316
rect 49007 6276 49424 6304
rect 49007 6273 49019 6276
rect 48961 6267 49019 6273
rect 49418 6264 49424 6276
rect 49476 6264 49482 6316
rect 49602 6304 49608 6316
rect 49563 6276 49608 6304
rect 49602 6264 49608 6276
rect 49660 6264 49666 6316
rect 49786 6313 49792 6316
rect 49743 6307 49792 6313
rect 49743 6273 49755 6307
rect 49789 6273 49792 6307
rect 49743 6267 49792 6273
rect 49786 6264 49792 6267
rect 49844 6264 49850 6316
rect 49973 6307 50031 6313
rect 49973 6273 49985 6307
rect 50019 6273 50031 6307
rect 52730 6304 52736 6316
rect 52691 6276 52736 6304
rect 49973 6267 50031 6273
rect 46474 6236 46480 6248
rect 46216 6208 46480 6236
rect 41874 6168 41880 6180
rect 40144 6140 41880 6168
rect 41874 6128 41880 6140
rect 41932 6168 41938 6180
rect 42610 6168 42616 6180
rect 41932 6140 42616 6168
rect 41932 6128 41938 6140
rect 42610 6128 42616 6140
rect 42668 6168 42674 6180
rect 42886 6168 42892 6180
rect 42668 6140 42892 6168
rect 42668 6128 42674 6140
rect 42886 6128 42892 6140
rect 42944 6128 42950 6180
rect 44100 6168 44128 6208
rect 46474 6196 46480 6208
rect 46532 6196 46538 6248
rect 48590 6168 48596 6180
rect 44100 6140 48596 6168
rect 48590 6128 48596 6140
rect 48648 6128 48654 6180
rect 49510 6128 49516 6180
rect 49568 6168 49574 6180
rect 49988 6168 50016 6267
rect 52730 6264 52736 6276
rect 52788 6264 52794 6316
rect 53024 6313 53052 6344
rect 54846 6332 54852 6344
rect 54904 6332 54910 6384
rect 53009 6307 53067 6313
rect 53009 6273 53021 6307
rect 53055 6273 53067 6307
rect 53009 6267 53067 6273
rect 53101 6307 53159 6313
rect 53101 6273 53113 6307
rect 53147 6273 53159 6307
rect 53101 6267 53159 6273
rect 53116 6236 53144 6267
rect 53024 6208 53144 6236
rect 52362 6168 52368 6180
rect 49568 6140 52368 6168
rect 49568 6128 49574 6140
rect 52362 6128 52368 6140
rect 52420 6168 52426 6180
rect 53024 6168 53052 6208
rect 52420 6140 53052 6168
rect 52420 6128 52426 6140
rect 32140 6072 33088 6100
rect 33134 6060 33140 6112
rect 33192 6100 33198 6112
rect 36998 6100 37004 6112
rect 33192 6072 37004 6100
rect 33192 6060 33198 6072
rect 36998 6060 37004 6072
rect 37056 6060 37062 6112
rect 39761 6103 39819 6109
rect 39761 6069 39773 6103
rect 39807 6100 39819 6103
rect 39942 6100 39948 6112
rect 39807 6072 39948 6100
rect 39807 6069 39819 6072
rect 39761 6063 39819 6069
rect 39942 6060 39948 6072
rect 40000 6060 40006 6112
rect 42705 6103 42763 6109
rect 42705 6069 42717 6103
rect 42751 6100 42763 6103
rect 43806 6100 43812 6112
rect 42751 6072 43812 6100
rect 42751 6069 42763 6072
rect 42705 6063 42763 6069
rect 43806 6060 43812 6072
rect 43864 6060 43870 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 5442 5896 5448 5908
rect 5403 5868 5448 5896
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 9122 5896 9128 5908
rect 8720 5868 9128 5896
rect 8720 5856 8726 5868
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 11974 5896 11980 5908
rect 10336 5868 11980 5896
rect 1854 5760 1860 5772
rect 1815 5732 1860 5760
rect 1854 5720 1860 5732
rect 1912 5720 1918 5772
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 10336 5769 10364 5868
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 12253 5899 12311 5905
rect 12253 5865 12265 5899
rect 12299 5896 12311 5899
rect 12342 5896 12348 5908
rect 12299 5868 12348 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 15197 5899 15255 5905
rect 15197 5865 15209 5899
rect 15243 5896 15255 5899
rect 16850 5896 16856 5908
rect 15243 5868 16856 5896
rect 15243 5865 15255 5868
rect 15197 5859 15255 5865
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 21266 5856 21272 5908
rect 21324 5896 21330 5908
rect 21453 5899 21511 5905
rect 21453 5896 21465 5899
rect 21324 5868 21465 5896
rect 21324 5856 21330 5868
rect 21453 5865 21465 5868
rect 21499 5865 21511 5899
rect 21453 5859 21511 5865
rect 27430 5856 27436 5908
rect 27488 5896 27494 5908
rect 27982 5896 27988 5908
rect 27488 5868 27988 5896
rect 27488 5856 27494 5868
rect 27982 5856 27988 5868
rect 28040 5896 28046 5908
rect 28534 5896 28540 5908
rect 28040 5868 28540 5896
rect 28040 5856 28046 5868
rect 28534 5856 28540 5868
rect 28592 5856 28598 5908
rect 28902 5856 28908 5908
rect 28960 5896 28966 5908
rect 29733 5899 29791 5905
rect 29733 5896 29745 5899
rect 28960 5868 29745 5896
rect 28960 5856 28966 5868
rect 29733 5865 29745 5868
rect 29779 5896 29791 5899
rect 31570 5896 31576 5908
rect 29779 5868 31576 5896
rect 29779 5865 29791 5868
rect 29733 5859 29791 5865
rect 31570 5856 31576 5868
rect 31628 5856 31634 5908
rect 38746 5896 38752 5908
rect 31956 5868 38752 5896
rect 15102 5788 15108 5840
rect 15160 5828 15166 5840
rect 19334 5828 19340 5840
rect 15160 5800 19340 5828
rect 15160 5788 15166 5800
rect 19334 5788 19340 5800
rect 19392 5788 19398 5840
rect 21085 5831 21143 5837
rect 21085 5797 21097 5831
rect 21131 5828 21143 5831
rect 22186 5828 22192 5840
rect 21131 5800 22192 5828
rect 21131 5797 21143 5800
rect 21085 5791 21143 5797
rect 22186 5788 22192 5800
rect 22244 5828 22250 5840
rect 22327 5831 22385 5837
rect 22327 5828 22339 5831
rect 22244 5800 22339 5828
rect 22244 5788 22250 5800
rect 22327 5797 22339 5800
rect 22373 5797 22385 5831
rect 26326 5828 26332 5840
rect 22327 5791 22385 5797
rect 25148 5800 26332 5828
rect 10137 5763 10195 5769
rect 10137 5760 10149 5763
rect 5592 5732 10149 5760
rect 5592 5720 5598 5732
rect 10137 5729 10149 5732
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 14458 5720 14464 5772
rect 14516 5760 14522 5772
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 14516 5732 15577 5760
rect 14516 5720 14522 5732
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 17402 5760 17408 5772
rect 15703 5732 17408 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 22002 5720 22008 5772
rect 22060 5760 22066 5772
rect 23753 5763 23811 5769
rect 23753 5760 23765 5763
rect 22060 5732 23765 5760
rect 22060 5720 22066 5732
rect 23753 5729 23765 5732
rect 23799 5729 23811 5763
rect 23753 5723 23811 5729
rect 2124 5695 2182 5701
rect 2124 5661 2136 5695
rect 2170 5692 2182 5695
rect 2590 5692 2596 5704
rect 2170 5664 2596 5692
rect 2170 5661 2182 5664
rect 2124 5655 2182 5661
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 2746 5664 4077 5692
rect 2038 5584 2044 5636
rect 2096 5624 2102 5636
rect 2746 5624 2774 5664
rect 4065 5661 4077 5664
rect 4111 5692 4123 5695
rect 4154 5692 4160 5704
rect 4111 5664 4160 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4332 5695 4390 5701
rect 4332 5661 4344 5695
rect 4378 5692 4390 5695
rect 4798 5692 4804 5704
rect 4378 5664 4804 5692
rect 4378 5661 4390 5664
rect 4332 5655 4390 5661
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 8938 5692 8944 5704
rect 8899 5664 8944 5692
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5692 9183 5695
rect 9766 5692 9772 5704
rect 9171 5664 9772 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 10873 5695 10931 5701
rect 10873 5661 10885 5695
rect 10919 5692 10931 5695
rect 10962 5692 10968 5704
rect 10919 5664 10968 5692
rect 10919 5661 10931 5664
rect 10873 5655 10931 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 11882 5652 11888 5704
rect 11940 5692 11946 5704
rect 15194 5692 15200 5704
rect 11940 5664 15200 5692
rect 11940 5652 11946 5664
rect 15194 5652 15200 5664
rect 15252 5692 15258 5704
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 15252 5664 15393 5692
rect 15252 5652 15258 5664
rect 15381 5661 15393 5664
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5692 15531 5695
rect 17126 5692 17132 5704
rect 15519 5664 17132 5692
rect 15519 5661 15531 5664
rect 15473 5655 15531 5661
rect 2096 5596 2774 5624
rect 2096 5584 2102 5596
rect 3326 5584 3332 5636
rect 3384 5624 3390 5636
rect 8110 5624 8116 5636
rect 3384 5596 8116 5624
rect 3384 5584 3390 5596
rect 8110 5584 8116 5596
rect 8168 5584 8174 5636
rect 11146 5633 11152 5636
rect 11140 5587 11152 5633
rect 11204 5624 11210 5636
rect 11204 5596 11240 5624
rect 11146 5584 11152 5587
rect 11204 5584 11210 5596
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 4890 5556 4896 5568
rect 3283 5528 4896 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 9033 5559 9091 5565
rect 9033 5556 9045 5559
rect 8628 5528 9045 5556
rect 8628 5516 8634 5528
rect 9033 5525 9045 5528
rect 9079 5525 9091 5559
rect 9674 5556 9680 5568
rect 9635 5528 9680 5556
rect 9033 5519 9091 5525
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 10045 5559 10103 5565
rect 10045 5525 10057 5559
rect 10091 5556 10103 5559
rect 15488 5556 15516 5655
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 22094 5652 22100 5704
rect 22152 5692 22158 5704
rect 22152 5664 22197 5692
rect 22152 5652 22158 5664
rect 23290 5652 23296 5704
rect 23348 5692 23354 5704
rect 25148 5702 25176 5800
rect 26326 5788 26332 5800
rect 26384 5788 26390 5840
rect 26970 5788 26976 5840
rect 27028 5828 27034 5840
rect 31956 5828 31984 5868
rect 38746 5856 38752 5868
rect 38804 5896 38810 5908
rect 52549 5899 52607 5905
rect 38804 5868 42472 5896
rect 38804 5856 38810 5868
rect 27028 5800 31984 5828
rect 32861 5831 32919 5837
rect 27028 5788 27034 5800
rect 25866 5760 25872 5772
rect 25516 5732 25872 5760
rect 25226 5705 25284 5711
rect 25226 5702 25238 5705
rect 23385 5695 23443 5701
rect 23385 5692 23397 5695
rect 23348 5664 23397 5692
rect 23348 5652 23354 5664
rect 23385 5661 23397 5664
rect 23431 5661 23443 5695
rect 25148 5674 25238 5702
rect 25226 5671 25238 5674
rect 25272 5671 25284 5705
rect 25226 5665 25284 5671
rect 25410 5695 25468 5701
rect 23385 5655 23443 5661
rect 25410 5661 25422 5695
rect 25456 5692 25468 5695
rect 25516 5692 25544 5732
rect 25866 5720 25872 5732
rect 25924 5720 25930 5772
rect 26786 5760 26792 5772
rect 26747 5732 26792 5760
rect 26786 5720 26792 5732
rect 26844 5720 26850 5772
rect 26878 5720 26884 5772
rect 26936 5760 26942 5772
rect 26936 5732 27660 5760
rect 26936 5720 26942 5732
rect 25456 5664 25544 5692
rect 25456 5661 25468 5664
rect 25410 5655 25468 5661
rect 25682 5652 25688 5704
rect 25740 5692 25746 5704
rect 26326 5692 26332 5704
rect 25740 5664 25785 5692
rect 26287 5664 26332 5692
rect 25740 5652 25746 5664
rect 26326 5652 26332 5664
rect 26384 5652 26390 5704
rect 27430 5692 27436 5704
rect 21450 5624 21456 5636
rect 21411 5596 21456 5624
rect 21450 5584 21456 5596
rect 21508 5584 21514 5636
rect 23569 5627 23627 5633
rect 23569 5593 23581 5627
rect 23615 5593 23627 5627
rect 25314 5624 25320 5636
rect 25275 5596 25320 5624
rect 23569 5587 23627 5593
rect 10091 5528 15516 5556
rect 21637 5559 21695 5565
rect 10091 5525 10103 5528
rect 10045 5519 10103 5525
rect 21637 5525 21649 5559
rect 21683 5556 21695 5559
rect 23584 5556 23612 5587
rect 25314 5584 25320 5596
rect 25372 5584 25378 5636
rect 25527 5627 25585 5633
rect 26418 5630 26424 5682
rect 26476 5630 26482 5682
rect 27391 5664 27436 5692
rect 27430 5652 27436 5664
rect 27488 5652 27494 5704
rect 27632 5701 27660 5732
rect 27750 5701 27778 5800
rect 32861 5797 32873 5831
rect 32907 5828 32919 5831
rect 33042 5828 33048 5840
rect 32907 5800 33048 5828
rect 32907 5797 32919 5800
rect 32861 5791 32919 5797
rect 33042 5788 33048 5800
rect 33100 5788 33106 5840
rect 38286 5828 38292 5840
rect 33336 5800 38292 5828
rect 33336 5760 33364 5800
rect 38286 5788 38292 5800
rect 38344 5788 38350 5840
rect 28828 5732 33364 5760
rect 27617 5695 27675 5701
rect 27617 5661 27629 5695
rect 27663 5661 27675 5695
rect 27617 5655 27675 5661
rect 27735 5695 27793 5701
rect 27735 5661 27747 5695
rect 27781 5661 27793 5695
rect 27890 5692 27896 5704
rect 27851 5664 27896 5692
rect 27735 5655 27793 5661
rect 27890 5652 27896 5664
rect 27948 5652 27954 5704
rect 28534 5692 28540 5704
rect 28495 5664 28540 5692
rect 28534 5652 28540 5664
rect 28592 5652 28598 5704
rect 28718 5692 28724 5704
rect 28679 5664 28724 5692
rect 28718 5652 28724 5664
rect 28776 5652 28782 5704
rect 28828 5701 28856 5732
rect 33410 5720 33416 5772
rect 33468 5760 33474 5772
rect 35529 5763 35587 5769
rect 35529 5760 35541 5763
rect 33468 5732 35541 5760
rect 33468 5720 33474 5732
rect 35529 5729 35541 5732
rect 35575 5729 35587 5763
rect 35529 5723 35587 5729
rect 35802 5720 35808 5772
rect 35860 5760 35866 5772
rect 36633 5763 36691 5769
rect 36633 5760 36645 5763
rect 35860 5732 36645 5760
rect 35860 5720 35866 5732
rect 36633 5729 36645 5732
rect 36679 5760 36691 5763
rect 37458 5760 37464 5772
rect 36679 5732 37464 5760
rect 36679 5729 36691 5732
rect 36633 5723 36691 5729
rect 37458 5720 37464 5732
rect 37516 5720 37522 5772
rect 39850 5760 39856 5772
rect 39811 5732 39856 5760
rect 39850 5720 39856 5732
rect 39908 5720 39914 5772
rect 41322 5720 41328 5772
rect 41380 5760 41386 5772
rect 42337 5763 42395 5769
rect 42337 5760 42349 5763
rect 41380 5732 42349 5760
rect 41380 5720 41386 5732
rect 42337 5729 42349 5732
rect 42383 5729 42395 5763
rect 42337 5723 42395 5729
rect 42444 5760 42472 5868
rect 52549 5865 52561 5899
rect 52595 5896 52607 5899
rect 52914 5896 52920 5908
rect 52595 5868 52920 5896
rect 52595 5865 52607 5868
rect 52549 5859 52607 5865
rect 52914 5856 52920 5868
rect 52972 5856 52978 5908
rect 42518 5788 42524 5840
rect 42576 5828 42582 5840
rect 50062 5828 50068 5840
rect 42576 5800 50068 5828
rect 42576 5788 42582 5800
rect 50062 5788 50068 5800
rect 50120 5788 50126 5840
rect 52454 5760 52460 5772
rect 42444 5732 43116 5760
rect 28828 5695 28897 5701
rect 28828 5664 28851 5695
rect 28839 5661 28851 5664
rect 28885 5661 28897 5695
rect 28839 5655 28897 5661
rect 28997 5695 29055 5701
rect 28997 5661 29009 5695
rect 29043 5661 29055 5695
rect 28997 5655 29055 5661
rect 25527 5593 25539 5627
rect 25573 5624 25585 5627
rect 26422 5627 26480 5630
rect 25573 5596 26280 5624
rect 25573 5593 25585 5596
rect 25527 5587 25585 5593
rect 25038 5556 25044 5568
rect 21683 5528 23612 5556
rect 24999 5528 25044 5556
rect 21683 5525 21695 5528
rect 21637 5519 21695 5525
rect 25038 5516 25044 5528
rect 25096 5516 25102 5568
rect 26142 5556 26148 5568
rect 26103 5528 26148 5556
rect 26142 5516 26148 5528
rect 26200 5516 26206 5568
rect 26252 5556 26280 5596
rect 26422 5593 26434 5627
rect 26468 5593 26480 5627
rect 26422 5587 26480 5593
rect 26510 5584 26516 5636
rect 26568 5624 26574 5636
rect 26651 5627 26709 5633
rect 26568 5596 26613 5624
rect 26568 5584 26574 5596
rect 26651 5593 26663 5627
rect 26697 5624 26709 5627
rect 26970 5624 26976 5636
rect 26697 5596 26976 5624
rect 26697 5593 26709 5596
rect 26651 5587 26709 5593
rect 26666 5556 26694 5587
rect 26970 5584 26976 5596
rect 27028 5584 27034 5636
rect 27522 5624 27528 5636
rect 27483 5596 27528 5624
rect 27522 5584 27528 5596
rect 27580 5624 27586 5636
rect 28629 5627 28687 5633
rect 28629 5624 28641 5627
rect 27580 5596 28641 5624
rect 27580 5584 27586 5596
rect 28629 5593 28641 5596
rect 28675 5593 28687 5627
rect 29012 5624 29040 5655
rect 29454 5652 29460 5704
rect 29512 5692 29518 5704
rect 32309 5695 32367 5701
rect 29512 5664 31754 5692
rect 29512 5652 29518 5664
rect 29546 5624 29552 5636
rect 29012 5596 29552 5624
rect 28629 5587 28687 5593
rect 29546 5584 29552 5596
rect 29604 5584 29610 5636
rect 29765 5627 29823 5633
rect 29765 5593 29777 5627
rect 29811 5624 29823 5627
rect 31294 5624 31300 5636
rect 29811 5596 31300 5624
rect 29811 5593 29823 5596
rect 29765 5587 29823 5593
rect 31294 5584 31300 5596
rect 31352 5584 31358 5636
rect 26252 5528 26694 5556
rect 27249 5559 27307 5565
rect 27249 5525 27261 5559
rect 27295 5556 27307 5559
rect 27982 5556 27988 5568
rect 27295 5528 27988 5556
rect 27295 5525 27307 5528
rect 27249 5519 27307 5525
rect 27982 5516 27988 5528
rect 28040 5516 28046 5568
rect 28353 5559 28411 5565
rect 28353 5525 28365 5559
rect 28399 5556 28411 5559
rect 28994 5556 29000 5568
rect 28399 5528 29000 5556
rect 28399 5525 28411 5528
rect 28353 5519 28411 5525
rect 28994 5516 29000 5528
rect 29052 5516 29058 5568
rect 29914 5556 29920 5568
rect 29875 5528 29920 5556
rect 29914 5516 29920 5528
rect 29972 5516 29978 5568
rect 31726 5556 31754 5664
rect 32309 5661 32321 5695
rect 32355 5661 32367 5695
rect 32309 5655 32367 5661
rect 32324 5556 32352 5655
rect 32398 5652 32404 5704
rect 32456 5692 32462 5704
rect 32677 5695 32735 5701
rect 32677 5692 32689 5695
rect 32456 5664 32689 5692
rect 32456 5652 32462 5664
rect 32677 5661 32689 5664
rect 32723 5661 32735 5695
rect 33594 5692 33600 5704
rect 32677 5655 32735 5661
rect 32968 5664 33600 5692
rect 32490 5624 32496 5636
rect 32451 5596 32496 5624
rect 32490 5584 32496 5596
rect 32548 5584 32554 5636
rect 32585 5627 32643 5633
rect 32585 5593 32597 5627
rect 32631 5624 32643 5627
rect 32968 5624 32996 5664
rect 33594 5652 33600 5664
rect 33652 5652 33658 5704
rect 35713 5695 35771 5701
rect 35713 5661 35725 5695
rect 35759 5692 35771 5695
rect 36262 5692 36268 5704
rect 35759 5664 36268 5692
rect 35759 5661 35771 5664
rect 35713 5655 35771 5661
rect 36262 5652 36268 5664
rect 36320 5652 36326 5704
rect 36446 5692 36452 5704
rect 36407 5664 36452 5692
rect 36446 5652 36452 5664
rect 36504 5652 36510 5704
rect 38105 5695 38163 5701
rect 38105 5661 38117 5695
rect 38151 5692 38163 5695
rect 38562 5692 38568 5704
rect 38151 5664 38568 5692
rect 38151 5661 38163 5664
rect 38105 5655 38163 5661
rect 38562 5652 38568 5664
rect 38620 5652 38626 5704
rect 39942 5652 39948 5704
rect 40000 5692 40006 5704
rect 40109 5695 40167 5701
rect 40109 5692 40121 5695
rect 40000 5664 40121 5692
rect 40000 5652 40006 5664
rect 40109 5661 40121 5664
rect 40155 5661 40167 5695
rect 41874 5692 41880 5704
rect 41835 5664 41880 5692
rect 40109 5655 40167 5661
rect 41874 5652 41880 5664
rect 41932 5652 41938 5704
rect 41966 5652 41972 5704
rect 42024 5692 42030 5704
rect 42199 5695 42257 5701
rect 42024 5664 42069 5692
rect 42024 5652 42030 5664
rect 42199 5661 42211 5695
rect 42245 5692 42257 5695
rect 42444 5692 42472 5732
rect 42245 5664 42472 5692
rect 42245 5661 42257 5664
rect 42199 5655 42257 5661
rect 42886 5652 42892 5704
rect 42944 5692 42950 5704
rect 42981 5695 43039 5701
rect 42981 5692 42993 5695
rect 42944 5664 42993 5692
rect 42944 5652 42950 5664
rect 42981 5661 42993 5664
rect 43027 5661 43039 5695
rect 43088 5692 43116 5732
rect 52012 5732 52460 5760
rect 43283 5695 43341 5701
rect 43283 5692 43295 5695
rect 43088 5664 43295 5692
rect 42981 5655 43039 5661
rect 43283 5661 43295 5664
rect 43329 5661 43341 5695
rect 43283 5655 43341 5661
rect 43441 5695 43499 5701
rect 43441 5661 43453 5695
rect 43487 5692 43499 5695
rect 46014 5692 46020 5704
rect 43487 5664 46020 5692
rect 43487 5661 43499 5664
rect 43441 5655 43499 5661
rect 46014 5652 46020 5664
rect 46072 5652 46078 5704
rect 52012 5701 52040 5732
rect 52454 5720 52460 5732
rect 52512 5720 52518 5772
rect 51997 5695 52055 5701
rect 51997 5661 52009 5695
rect 52043 5661 52055 5695
rect 52178 5692 52184 5704
rect 52139 5664 52184 5692
rect 51997 5655 52055 5661
rect 52178 5652 52184 5664
rect 52236 5652 52242 5704
rect 52362 5692 52368 5704
rect 52323 5664 52368 5692
rect 52362 5652 52368 5664
rect 52420 5652 52426 5704
rect 53009 5695 53067 5701
rect 53009 5661 53021 5695
rect 53055 5692 53067 5695
rect 53098 5692 53104 5704
rect 53055 5664 53104 5692
rect 53055 5661 53067 5664
rect 53009 5655 53067 5661
rect 53098 5652 53104 5664
rect 53156 5652 53162 5704
rect 53282 5701 53288 5704
rect 53276 5692 53288 5701
rect 53243 5664 53288 5692
rect 53276 5655 53288 5664
rect 53282 5652 53288 5655
rect 53340 5652 53346 5704
rect 42061 5627 42119 5633
rect 42061 5624 42073 5627
rect 32631 5596 32996 5624
rect 33152 5596 42073 5624
rect 32631 5593 32643 5596
rect 32585 5587 32643 5593
rect 31726 5528 32352 5556
rect 32674 5516 32680 5568
rect 32732 5556 32738 5568
rect 33152 5556 33180 5596
rect 42061 5593 42073 5596
rect 42107 5593 42119 5627
rect 42702 5624 42708 5636
rect 42061 5587 42119 5593
rect 42168 5596 42708 5624
rect 32732 5528 33180 5556
rect 32732 5516 32738 5528
rect 33318 5516 33324 5568
rect 33376 5556 33382 5568
rect 35710 5556 35716 5568
rect 33376 5528 35716 5556
rect 33376 5516 33382 5528
rect 35710 5516 35716 5528
rect 35768 5516 35774 5568
rect 35894 5556 35900 5568
rect 35855 5528 35900 5556
rect 35894 5516 35900 5528
rect 35952 5516 35958 5568
rect 39850 5516 39856 5568
rect 39908 5556 39914 5568
rect 40310 5556 40316 5568
rect 39908 5528 40316 5556
rect 39908 5516 39914 5528
rect 40310 5516 40316 5528
rect 40368 5516 40374 5568
rect 40402 5516 40408 5568
rect 40460 5556 40466 5568
rect 41233 5559 41291 5565
rect 41233 5556 41245 5559
rect 40460 5528 41245 5556
rect 40460 5516 40466 5528
rect 41233 5525 41245 5528
rect 41279 5556 41291 5559
rect 41322 5556 41328 5568
rect 41279 5528 41328 5556
rect 41279 5525 41291 5528
rect 41233 5519 41291 5525
rect 41322 5516 41328 5528
rect 41380 5516 41386 5568
rect 41690 5556 41696 5568
rect 41651 5528 41696 5556
rect 41690 5516 41696 5528
rect 41748 5516 41754 5568
rect 41966 5516 41972 5568
rect 42024 5556 42030 5568
rect 42168 5556 42196 5596
rect 42702 5584 42708 5596
rect 42760 5624 42766 5636
rect 43073 5627 43131 5633
rect 43073 5624 43085 5627
rect 42760 5596 43085 5624
rect 42760 5584 42766 5596
rect 43073 5593 43085 5596
rect 43119 5593 43131 5627
rect 43073 5587 43131 5593
rect 43165 5627 43223 5633
rect 43165 5593 43177 5627
rect 43211 5593 43223 5627
rect 43165 5587 43223 5593
rect 42794 5556 42800 5568
rect 42024 5528 42196 5556
rect 42755 5528 42800 5556
rect 42024 5516 42030 5528
rect 42794 5516 42800 5528
rect 42852 5516 42858 5568
rect 42978 5516 42984 5568
rect 43036 5556 43042 5568
rect 43180 5556 43208 5587
rect 45370 5584 45376 5636
rect 45428 5624 45434 5636
rect 46201 5627 46259 5633
rect 46201 5624 46213 5627
rect 45428 5596 46213 5624
rect 45428 5584 45434 5596
rect 46201 5593 46213 5596
rect 46247 5593 46259 5627
rect 46382 5624 46388 5636
rect 46343 5596 46388 5624
rect 46201 5587 46259 5593
rect 46382 5584 46388 5596
rect 46440 5624 46446 5636
rect 49510 5624 49516 5636
rect 46440 5596 49516 5624
rect 46440 5584 46446 5596
rect 49510 5584 49516 5596
rect 49568 5584 49574 5636
rect 52273 5627 52331 5633
rect 52273 5593 52285 5627
rect 52319 5593 52331 5627
rect 52273 5587 52331 5593
rect 43036 5528 43208 5556
rect 52288 5556 52316 5587
rect 52730 5556 52736 5568
rect 52288 5528 52736 5556
rect 43036 5516 43042 5528
rect 52730 5516 52736 5528
rect 52788 5556 52794 5568
rect 54386 5556 54392 5568
rect 52788 5528 54392 5556
rect 52788 5516 52794 5528
rect 54386 5516 54392 5528
rect 54444 5516 54450 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 4709 5355 4767 5361
rect 2700 5324 4660 5352
rect 1854 5284 1860 5296
rect 1815 5256 1860 5284
rect 1854 5244 1860 5256
rect 1912 5244 1918 5296
rect 2700 5225 2728 5324
rect 4632 5284 4660 5324
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 5534 5352 5540 5364
rect 4755 5324 5540 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 8846 5352 8852 5364
rect 8803 5324 8852 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 10781 5355 10839 5361
rect 10781 5321 10793 5355
rect 10827 5352 10839 5355
rect 11146 5352 11152 5364
rect 10827 5324 11152 5352
rect 10827 5321 10839 5324
rect 10781 5315 10839 5321
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 14826 5312 14832 5364
rect 14884 5352 14890 5364
rect 19426 5352 19432 5364
rect 14884 5324 19432 5352
rect 14884 5312 14890 5324
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22373 5355 22431 5361
rect 22373 5352 22385 5355
rect 22152 5324 22385 5352
rect 22152 5312 22158 5324
rect 22373 5321 22385 5324
rect 22419 5321 22431 5355
rect 22373 5315 22431 5321
rect 25682 5312 25688 5364
rect 25740 5352 25746 5364
rect 32306 5352 32312 5364
rect 25740 5324 32312 5352
rect 25740 5312 25746 5324
rect 32306 5312 32312 5324
rect 32364 5312 32370 5364
rect 32674 5312 32680 5364
rect 32732 5352 32738 5364
rect 32861 5355 32919 5361
rect 32861 5352 32873 5355
rect 32732 5324 32873 5352
rect 32732 5312 32738 5324
rect 32861 5321 32873 5324
rect 32907 5321 32919 5355
rect 32861 5315 32919 5321
rect 32950 5312 32956 5364
rect 33008 5312 33014 5364
rect 33134 5312 33140 5364
rect 33192 5352 33198 5364
rect 35986 5352 35992 5364
rect 33192 5324 35992 5352
rect 33192 5312 33198 5324
rect 35986 5312 35992 5324
rect 36044 5352 36050 5364
rect 36081 5355 36139 5361
rect 36081 5352 36093 5355
rect 36044 5324 36093 5352
rect 36044 5312 36050 5324
rect 36081 5321 36093 5324
rect 36127 5321 36139 5355
rect 36081 5315 36139 5321
rect 36541 5355 36599 5361
rect 36541 5321 36553 5355
rect 36587 5321 36599 5355
rect 38746 5352 38752 5364
rect 38707 5324 38752 5352
rect 36541 5315 36599 5321
rect 4632 5256 8432 5284
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5185 2743 5219
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 2685 5179 2743 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 4212 5188 4261 5216
rect 4212 5176 4218 5188
rect 4249 5185 4261 5188
rect 4295 5216 4307 5219
rect 4798 5216 4804 5228
rect 4295 5188 4804 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 4908 5148 4936 5179
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 7633 5219 7691 5225
rect 7633 5216 7645 5219
rect 7340 5188 7645 5216
rect 7340 5176 7346 5188
rect 7633 5185 7645 5188
rect 7679 5185 7691 5219
rect 7633 5179 7691 5185
rect 3844 5120 4936 5148
rect 7377 5151 7435 5157
rect 3844 5108 3850 5120
rect 7377 5117 7389 5151
rect 7423 5117 7435 5151
rect 8404 5148 8432 5256
rect 8478 5244 8484 5296
rect 8536 5284 8542 5296
rect 29914 5284 29920 5296
rect 8536 5256 25452 5284
rect 8536 5244 8542 5256
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 9732 5188 10977 5216
rect 9732 5176 9738 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 14826 5216 14832 5228
rect 14787 5188 14832 5216
rect 10965 5179 11023 5185
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 15010 5216 15016 5228
rect 14971 5188 15016 5216
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 15105 5219 15163 5225
rect 15105 5185 15117 5219
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 10870 5148 10876 5160
rect 8404 5120 10876 5148
rect 7377 5111 7435 5117
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 2866 5012 2872 5024
rect 2827 4984 2872 5012
rect 2866 4972 2872 4984
rect 2924 4972 2930 5024
rect 3418 5012 3424 5024
rect 3379 4984 3424 5012
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 4065 5015 4123 5021
rect 4065 5012 4077 5015
rect 3568 4984 4077 5012
rect 3568 4972 3574 4984
rect 4065 4981 4077 4984
rect 4111 4981 4123 5015
rect 4065 4975 4123 4981
rect 4798 4972 4804 5024
rect 4856 5012 4862 5024
rect 5258 5012 5264 5024
rect 4856 4984 5264 5012
rect 4856 4972 4862 4984
rect 5258 4972 5264 4984
rect 5316 5012 5322 5024
rect 7392 5012 7420 5111
rect 10870 5108 10876 5120
rect 10928 5108 10934 5160
rect 13630 5108 13636 5160
rect 13688 5148 13694 5160
rect 15120 5148 15148 5179
rect 18322 5176 18328 5228
rect 18380 5216 18386 5228
rect 18417 5219 18475 5225
rect 18417 5216 18429 5219
rect 18380 5188 18429 5216
rect 18380 5176 18386 5188
rect 18417 5185 18429 5188
rect 18463 5185 18475 5219
rect 18417 5179 18475 5185
rect 19061 5219 19119 5225
rect 19061 5185 19073 5219
rect 19107 5185 19119 5219
rect 19061 5179 19119 5185
rect 19245 5219 19303 5225
rect 19245 5185 19257 5219
rect 19291 5216 19303 5219
rect 20070 5216 20076 5228
rect 19291 5188 20076 5216
rect 19291 5185 19303 5188
rect 19245 5179 19303 5185
rect 13688 5120 15148 5148
rect 13688 5108 13694 5120
rect 18432 5080 18460 5179
rect 19076 5148 19104 5179
rect 20070 5176 20076 5188
rect 20128 5176 20134 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21928 5188 22017 5216
rect 20254 5148 20260 5160
rect 19076 5120 20260 5148
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 21818 5148 21824 5160
rect 21779 5120 21824 5148
rect 21818 5108 21824 5120
rect 21876 5108 21882 5160
rect 21634 5080 21640 5092
rect 18432 5052 21640 5080
rect 21634 5040 21640 5052
rect 21692 5080 21698 5092
rect 21928 5080 21956 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 22097 5219 22155 5225
rect 22097 5185 22109 5219
rect 22143 5185 22155 5219
rect 22097 5179 22155 5185
rect 21692 5052 21956 5080
rect 21692 5040 21698 5052
rect 8938 5012 8944 5024
rect 5316 4984 8944 5012
rect 5316 4972 5322 4984
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 14642 5012 14648 5024
rect 14603 4984 14648 5012
rect 14642 4972 14648 4984
rect 14700 4972 14706 5024
rect 18506 5012 18512 5024
rect 18467 4984 18512 5012
rect 18506 4972 18512 4984
rect 18564 4972 18570 5024
rect 19426 5012 19432 5024
rect 19387 4984 19432 5012
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 20070 4972 20076 5024
rect 20128 5012 20134 5024
rect 22112 5012 22140 5179
rect 22186 5176 22192 5228
rect 22244 5216 22250 5228
rect 25222 5216 25228 5228
rect 22244 5188 25228 5216
rect 22244 5176 22250 5188
rect 25222 5176 25228 5188
rect 25280 5176 25286 5228
rect 25424 5080 25452 5256
rect 25700 5256 27844 5284
rect 25498 5176 25504 5228
rect 25556 5216 25562 5228
rect 25700 5225 25728 5256
rect 25685 5219 25743 5225
rect 25685 5216 25697 5219
rect 25556 5188 25697 5216
rect 25556 5176 25562 5188
rect 25685 5185 25697 5188
rect 25731 5185 25743 5219
rect 25685 5179 25743 5185
rect 25869 5219 25927 5225
rect 25869 5185 25881 5219
rect 25915 5216 25927 5219
rect 26142 5216 26148 5228
rect 25915 5188 26148 5216
rect 25915 5185 25927 5188
rect 25869 5179 25927 5185
rect 26142 5176 26148 5188
rect 26200 5176 26206 5228
rect 27816 5225 27844 5256
rect 28092 5256 29920 5284
rect 27801 5219 27859 5225
rect 27801 5185 27813 5219
rect 27847 5185 27859 5219
rect 27982 5216 27988 5228
rect 27943 5188 27988 5216
rect 27801 5179 27859 5185
rect 25961 5151 26019 5157
rect 25961 5117 25973 5151
rect 26007 5148 26019 5151
rect 27522 5148 27528 5160
rect 26007 5120 27528 5148
rect 26007 5117 26019 5120
rect 25961 5111 26019 5117
rect 27522 5108 27528 5120
rect 27580 5108 27586 5160
rect 27816 5148 27844 5179
rect 27982 5176 27988 5188
rect 28040 5176 28046 5228
rect 28092 5225 28120 5256
rect 29914 5244 29920 5256
rect 29972 5244 29978 5296
rect 30466 5284 30472 5296
rect 30024 5256 30472 5284
rect 28077 5219 28135 5225
rect 28077 5185 28089 5219
rect 28123 5185 28135 5219
rect 28077 5179 28135 5185
rect 28813 5219 28871 5225
rect 28813 5185 28825 5219
rect 28859 5185 28871 5219
rect 28994 5216 29000 5228
rect 28955 5188 29000 5216
rect 28813 5179 28871 5185
rect 28828 5148 28856 5179
rect 28994 5176 29000 5188
rect 29052 5176 29058 5228
rect 29089 5219 29147 5225
rect 29089 5185 29101 5219
rect 29135 5216 29147 5219
rect 29822 5216 29828 5228
rect 29135 5188 29828 5216
rect 29135 5185 29147 5188
rect 29089 5179 29147 5185
rect 29822 5176 29828 5188
rect 29880 5176 29886 5228
rect 27816 5120 28856 5148
rect 28828 5080 28856 5120
rect 29917 5151 29975 5157
rect 29917 5117 29929 5151
rect 29963 5148 29975 5151
rect 30024 5148 30052 5256
rect 30466 5244 30472 5256
rect 30524 5284 30530 5296
rect 31110 5284 31116 5296
rect 30524 5256 31116 5284
rect 30524 5244 30530 5256
rect 31110 5244 31116 5256
rect 31168 5244 31174 5296
rect 31294 5284 31300 5296
rect 31255 5256 31300 5284
rect 31294 5244 31300 5256
rect 31352 5244 31358 5296
rect 32122 5244 32128 5296
rect 32180 5284 32186 5296
rect 32585 5287 32643 5293
rect 32180 5256 32352 5284
rect 32180 5244 32186 5256
rect 30098 5176 30104 5228
rect 30156 5216 30162 5228
rect 32324 5225 32352 5256
rect 32585 5253 32597 5287
rect 32631 5284 32643 5287
rect 32968 5284 32996 5312
rect 34146 5284 34152 5296
rect 32631 5256 34152 5284
rect 32631 5253 32643 5256
rect 32585 5247 32643 5253
rect 34146 5244 34152 5256
rect 34204 5244 34210 5296
rect 34968 5287 35026 5293
rect 34968 5253 34980 5287
rect 35014 5284 35026 5287
rect 36556 5284 36584 5315
rect 38746 5312 38752 5324
rect 38804 5312 38810 5364
rect 40586 5312 40592 5364
rect 40644 5352 40650 5364
rect 40681 5355 40739 5361
rect 40681 5352 40693 5355
rect 40644 5324 40693 5352
rect 40644 5312 40650 5324
rect 40681 5321 40693 5324
rect 40727 5321 40739 5355
rect 40681 5315 40739 5321
rect 40954 5312 40960 5364
rect 41012 5352 41018 5364
rect 43073 5355 43131 5361
rect 41012 5324 43024 5352
rect 41012 5312 41018 5324
rect 35014 5256 36584 5284
rect 35014 5253 35026 5256
rect 34968 5247 35026 5253
rect 38286 5244 38292 5296
rect 38344 5284 38350 5296
rect 40218 5284 40224 5296
rect 38344 5256 40224 5284
rect 38344 5244 38350 5256
rect 40218 5244 40224 5256
rect 40276 5284 40282 5296
rect 40313 5287 40371 5293
rect 40313 5284 40325 5287
rect 40276 5256 40325 5284
rect 40276 5244 40282 5256
rect 40313 5253 40325 5256
rect 40359 5253 40371 5287
rect 42702 5284 42708 5296
rect 42663 5256 42708 5284
rect 40313 5247 40371 5253
rect 42702 5244 42708 5256
rect 42760 5244 42766 5296
rect 42886 5244 42892 5296
rect 42944 5293 42950 5296
rect 42944 5287 42963 5293
rect 42951 5253 42963 5287
rect 42996 5284 43024 5324
rect 43073 5321 43085 5355
rect 43119 5352 43131 5355
rect 43162 5352 43168 5364
rect 43119 5324 43168 5352
rect 43119 5321 43131 5324
rect 43073 5315 43131 5321
rect 43162 5312 43168 5324
rect 43220 5312 43226 5364
rect 49878 5352 49884 5364
rect 49620 5324 49884 5352
rect 44358 5284 44364 5296
rect 42996 5256 44364 5284
rect 42944 5247 42963 5253
rect 42944 5244 42950 5247
rect 44358 5244 44364 5256
rect 44416 5284 44422 5296
rect 45370 5284 45376 5296
rect 44416 5256 45376 5284
rect 44416 5244 44422 5256
rect 45370 5244 45376 5256
rect 45428 5244 45434 5296
rect 32309 5219 32367 5225
rect 30156 5188 32260 5216
rect 30156 5176 30162 5188
rect 29963 5120 30052 5148
rect 30193 5151 30251 5157
rect 29963 5117 29975 5120
rect 29917 5111 29975 5117
rect 30193 5117 30205 5151
rect 30239 5117 30251 5151
rect 32232 5148 32260 5188
rect 32309 5185 32321 5219
rect 32355 5185 32367 5219
rect 32490 5216 32496 5228
rect 32451 5188 32496 5216
rect 32309 5179 32367 5185
rect 32490 5176 32496 5188
rect 32548 5176 32554 5228
rect 32677 5219 32735 5225
rect 32677 5185 32689 5219
rect 32723 5216 32735 5219
rect 32950 5216 32956 5228
rect 32723 5188 32956 5216
rect 32723 5185 32735 5188
rect 32677 5179 32735 5185
rect 32950 5176 32956 5188
rect 33008 5216 33014 5228
rect 33008 5188 35756 5216
rect 33008 5176 33014 5188
rect 32232 5120 34652 5148
rect 30193 5111 30251 5117
rect 30208 5080 30236 5111
rect 25424 5052 28764 5080
rect 28828 5052 30236 5080
rect 20128 4984 22140 5012
rect 25501 5015 25559 5021
rect 20128 4972 20134 4984
rect 25501 4981 25513 5015
rect 25547 5012 25559 5015
rect 26326 5012 26332 5024
rect 25547 4984 26332 5012
rect 25547 4981 25559 4984
rect 25501 4975 25559 4981
rect 26326 4972 26332 4984
rect 26384 4972 26390 5024
rect 27614 5012 27620 5024
rect 27575 4984 27620 5012
rect 27614 4972 27620 4984
rect 27672 4972 27678 5024
rect 28626 5012 28632 5024
rect 28587 4984 28632 5012
rect 28626 4972 28632 4984
rect 28684 4972 28690 5024
rect 28736 5012 28764 5052
rect 31202 5012 31208 5024
rect 28736 4984 31208 5012
rect 31202 4972 31208 4984
rect 31260 4972 31266 5024
rect 31294 4972 31300 5024
rect 31352 5012 31358 5024
rect 31389 5015 31447 5021
rect 31389 5012 31401 5015
rect 31352 4984 31401 5012
rect 31352 4972 31358 4984
rect 31389 4981 31401 4984
rect 31435 5012 31447 5015
rect 34514 5012 34520 5024
rect 31435 4984 34520 5012
rect 31435 4981 31447 4984
rect 31389 4975 31447 4981
rect 34514 4972 34520 4984
rect 34572 4972 34578 5024
rect 34624 5012 34652 5120
rect 34698 5108 34704 5160
rect 34756 5148 34762 5160
rect 35728 5148 35756 5188
rect 35894 5176 35900 5228
rect 35952 5216 35958 5228
rect 36725 5219 36783 5225
rect 36725 5216 36737 5219
rect 35952 5188 36737 5216
rect 35952 5176 35958 5188
rect 36725 5185 36737 5188
rect 36771 5185 36783 5219
rect 36725 5179 36783 5185
rect 38562 5176 38568 5228
rect 38620 5216 38626 5228
rect 38657 5219 38715 5225
rect 38657 5216 38669 5219
rect 38620 5188 38669 5216
rect 38620 5176 38626 5188
rect 38657 5185 38669 5188
rect 38703 5185 38715 5219
rect 40126 5216 40132 5228
rect 40087 5188 40132 5216
rect 38657 5179 38715 5185
rect 40126 5176 40132 5188
rect 40184 5176 40190 5228
rect 40402 5216 40408 5228
rect 40363 5188 40408 5216
rect 40402 5176 40408 5188
rect 40460 5176 40466 5228
rect 40494 5176 40500 5228
rect 40552 5225 40558 5228
rect 40552 5219 40579 5225
rect 40567 5185 40579 5219
rect 40552 5179 40579 5185
rect 46201 5219 46259 5225
rect 46201 5185 46213 5219
rect 46247 5216 46259 5219
rect 47118 5216 47124 5228
rect 46247 5188 47124 5216
rect 46247 5185 46259 5188
rect 46201 5179 46259 5185
rect 40552 5176 40558 5179
rect 47118 5176 47124 5188
rect 47176 5176 47182 5228
rect 36170 5148 36176 5160
rect 34756 5120 34801 5148
rect 35728 5120 36176 5148
rect 34756 5108 34762 5120
rect 36170 5108 36176 5120
rect 36228 5108 36234 5160
rect 36446 5108 36452 5160
rect 36504 5148 36510 5160
rect 37277 5151 37335 5157
rect 37277 5148 37289 5151
rect 36504 5120 37289 5148
rect 36504 5108 36510 5120
rect 37277 5117 37289 5120
rect 37323 5117 37335 5151
rect 37550 5148 37556 5160
rect 37511 5120 37556 5148
rect 37277 5111 37335 5117
rect 37550 5108 37556 5120
rect 37608 5108 37614 5160
rect 46474 5148 46480 5160
rect 39868 5120 43392 5148
rect 46435 5120 46480 5148
rect 39868 5080 39896 5120
rect 40494 5080 40500 5092
rect 35912 5052 39896 5080
rect 40052 5052 40500 5080
rect 35912 5012 35940 5052
rect 34624 4984 35940 5012
rect 36170 4972 36176 5024
rect 36228 5012 36234 5024
rect 40052 5012 40080 5052
rect 40494 5040 40500 5052
rect 40552 5080 40558 5092
rect 43364 5080 43392 5120
rect 46474 5108 46480 5120
rect 46532 5108 46538 5160
rect 48222 5108 48228 5160
rect 48280 5148 48286 5160
rect 49620 5157 49648 5324
rect 49878 5312 49884 5324
rect 49936 5312 49942 5364
rect 50982 5352 50988 5364
rect 50943 5324 50988 5352
rect 50982 5312 50988 5324
rect 51040 5312 51046 5364
rect 49694 5176 49700 5228
rect 49752 5216 49758 5228
rect 49861 5219 49919 5225
rect 49861 5216 49873 5219
rect 49752 5188 49873 5216
rect 49752 5176 49758 5188
rect 49861 5185 49873 5188
rect 49907 5185 49919 5219
rect 49861 5179 49919 5185
rect 49605 5151 49663 5157
rect 49605 5148 49617 5151
rect 48280 5120 49617 5148
rect 48280 5108 48286 5120
rect 49605 5117 49617 5120
rect 49651 5117 49663 5151
rect 49605 5111 49663 5117
rect 46385 5083 46443 5089
rect 46385 5080 46397 5083
rect 40552 5052 43300 5080
rect 43364 5052 46397 5080
rect 40552 5040 40558 5052
rect 36228 4984 40080 5012
rect 36228 4972 36234 4984
rect 40126 4972 40132 5024
rect 40184 5012 40190 5024
rect 41414 5012 41420 5024
rect 40184 4984 41420 5012
rect 40184 4972 40190 4984
rect 41414 4972 41420 4984
rect 41472 4972 41478 5024
rect 41598 4972 41604 5024
rect 41656 5012 41662 5024
rect 42610 5012 42616 5024
rect 41656 4984 42616 5012
rect 41656 4972 41662 4984
rect 42610 4972 42616 4984
rect 42668 5012 42674 5024
rect 42889 5015 42947 5021
rect 42889 5012 42901 5015
rect 42668 4984 42901 5012
rect 42668 4972 42674 4984
rect 42889 4981 42901 4984
rect 42935 4981 42947 5015
rect 43272 5012 43300 5052
rect 46385 5049 46397 5052
rect 46431 5049 46443 5083
rect 46385 5043 46443 5049
rect 45462 5012 45468 5024
rect 43272 4984 45468 5012
rect 42889 4975 42947 4981
rect 45462 4972 45468 4984
rect 45520 4972 45526 5024
rect 46017 5015 46075 5021
rect 46017 4981 46029 5015
rect 46063 5012 46075 5015
rect 46750 5012 46756 5024
rect 46063 4984 46756 5012
rect 46063 4981 46075 4984
rect 46017 4975 46075 4981
rect 46750 4972 46756 4984
rect 46808 4972 46814 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 2041 4811 2099 4817
rect 2041 4808 2053 4811
rect 1412 4780 2053 4808
rect 1412 4613 1440 4780
rect 2041 4777 2053 4780
rect 2087 4808 2099 4811
rect 7282 4808 7288 4820
rect 2087 4780 7144 4808
rect 7243 4780 7288 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 1578 4700 1584 4752
rect 1636 4740 1642 4752
rect 2317 4743 2375 4749
rect 2317 4740 2329 4743
rect 1636 4712 2329 4740
rect 1636 4700 1642 4712
rect 2317 4709 2329 4712
rect 2363 4709 2375 4743
rect 2317 4703 2375 4709
rect 3970 4700 3976 4752
rect 4028 4740 4034 4752
rect 5261 4743 5319 4749
rect 5261 4740 5273 4743
rect 4028 4712 5273 4740
rect 4028 4700 4034 4712
rect 5261 4709 5273 4712
rect 5307 4709 5319 4743
rect 7116 4740 7144 4780
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 10321 4811 10379 4817
rect 10321 4808 10333 4811
rect 10100 4780 10333 4808
rect 10100 4768 10106 4780
rect 10321 4777 10333 4780
rect 10367 4777 10379 4811
rect 10321 4771 10379 4777
rect 15010 4768 15016 4820
rect 15068 4808 15074 4820
rect 15473 4811 15531 4817
rect 15473 4808 15485 4811
rect 15068 4780 15485 4808
rect 15068 4768 15074 4780
rect 15473 4777 15485 4780
rect 15519 4777 15531 4811
rect 15473 4771 15531 4777
rect 20254 4768 20260 4820
rect 20312 4808 20318 4820
rect 21266 4808 21272 4820
rect 20312 4780 21128 4808
rect 21227 4780 21272 4808
rect 20312 4768 20318 4780
rect 8478 4740 8484 4752
rect 7116 4712 8484 4740
rect 5261 4703 5319 4709
rect 8478 4700 8484 4712
rect 8536 4700 8542 4752
rect 21100 4740 21128 4780
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 22186 4808 22192 4820
rect 21468 4780 22192 4808
rect 21468 4740 21496 4780
rect 22186 4768 22192 4780
rect 22244 4768 22250 4820
rect 24486 4768 24492 4820
rect 24544 4808 24550 4820
rect 24765 4811 24823 4817
rect 24765 4808 24777 4811
rect 24544 4780 24777 4808
rect 24544 4768 24550 4780
rect 24765 4777 24777 4780
rect 24811 4777 24823 4811
rect 24765 4771 24823 4777
rect 25038 4768 25044 4820
rect 25096 4808 25102 4820
rect 25685 4811 25743 4817
rect 25685 4808 25697 4811
rect 25096 4780 25697 4808
rect 25096 4768 25102 4780
rect 25685 4777 25697 4780
rect 25731 4777 25743 4811
rect 25685 4771 25743 4777
rect 26513 4811 26571 4817
rect 26513 4777 26525 4811
rect 26559 4808 26571 4811
rect 27341 4811 27399 4817
rect 26559 4780 27292 4808
rect 26559 4777 26571 4780
rect 26513 4771 26571 4777
rect 21100 4712 21496 4740
rect 2884 4644 6960 4672
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4604 2191 4607
rect 2682 4604 2688 4616
rect 2179 4576 2688 4604
rect 2179 4573 2191 4576
rect 2133 4567 2191 4573
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 2884 4613 2912 4644
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 2958 4564 2964 4616
rect 3016 4604 3022 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3016 4576 3985 4604
rect 3016 4564 3022 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 4798 4604 4804 4616
rect 4759 4576 4804 4604
rect 3973 4567 4031 4573
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 4908 4576 5457 4604
rect 3142 4496 3148 4548
rect 3200 4536 3206 4548
rect 4908 4536 4936 4576
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 3200 4508 4936 4536
rect 3200 4496 3206 4508
rect 5350 4496 5356 4548
rect 5408 4536 5414 4548
rect 6104 4536 6132 4567
rect 5408 4508 6132 4536
rect 6932 4536 6960 4644
rect 7098 4632 7104 4684
rect 7156 4672 7162 4684
rect 8570 4672 8576 4684
rect 7156 4644 8576 4672
rect 7156 4632 7162 4644
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 11609 4675 11667 4681
rect 11609 4672 11621 4675
rect 10744 4644 11621 4672
rect 10744 4632 10750 4644
rect 11609 4641 11621 4644
rect 11655 4641 11667 4675
rect 11609 4635 11667 4641
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 13872 4644 14105 4672
rect 13872 4632 13878 4644
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 15933 4675 15991 4681
rect 15933 4641 15945 4675
rect 15979 4672 15991 4675
rect 16114 4672 16120 4684
rect 15979 4644 16120 4672
rect 15979 4641 15991 4644
rect 15933 4635 15991 4641
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 19426 4672 19432 4684
rect 19387 4644 19432 4672
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 21468 4681 21496 4712
rect 19521 4675 19579 4681
rect 19521 4641 19533 4675
rect 19567 4672 19579 4675
rect 20349 4675 20407 4681
rect 20349 4672 20361 4675
rect 19567 4644 20361 4672
rect 19567 4641 19579 4644
rect 19521 4635 19579 4641
rect 20349 4641 20361 4644
rect 20395 4641 20407 4675
rect 20349 4635 20407 4641
rect 21453 4675 21511 4681
rect 21453 4641 21465 4675
rect 21499 4672 21511 4675
rect 21634 4672 21640 4684
rect 21499 4644 21533 4672
rect 21595 4644 21640 4672
rect 21499 4641 21511 4644
rect 21453 4635 21511 4641
rect 7561 4607 7619 4613
rect 7561 4573 7573 4607
rect 7607 4604 7619 4607
rect 7742 4604 7748 4616
rect 7607 4576 7748 4604
rect 7607 4573 7619 4576
rect 7561 4567 7619 4573
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 8938 4604 8944 4616
rect 7892 4576 8340 4604
rect 8899 4576 8944 4604
rect 7892 4564 7898 4576
rect 8312 4536 8340 4576
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 11882 4604 11888 4616
rect 11839 4576 11888 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 11882 4564 11888 4576
rect 11940 4564 11946 4616
rect 14360 4607 14418 4613
rect 14360 4573 14372 4607
rect 14406 4604 14418 4607
rect 14642 4604 14648 4616
rect 14406 4576 14648 4604
rect 14406 4573 14418 4576
rect 14360 4567 14418 4573
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4604 16267 4607
rect 16482 4604 16488 4616
rect 16255 4576 16488 4604
rect 16255 4573 16267 4576
rect 16209 4567 16267 4573
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 9186 4539 9244 4545
rect 9186 4536 9198 4539
rect 6932 4508 8248 4536
rect 8312 4508 9198 4536
rect 5408 4496 5414 4508
rect 1118 4428 1124 4480
rect 1176 4468 1182 4480
rect 1581 4471 1639 4477
rect 1581 4468 1593 4471
rect 1176 4440 1593 4468
rect 1176 4428 1182 4440
rect 1581 4437 1593 4440
rect 1627 4437 1639 4471
rect 1581 4431 1639 4437
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3053 4471 3111 4477
rect 3053 4468 3065 4471
rect 2832 4440 3065 4468
rect 2832 4428 2838 4440
rect 3053 4437 3065 4440
rect 3099 4437 3111 4471
rect 4614 4468 4620 4480
rect 4575 4440 4620 4468
rect 3053 4431 3111 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 4706 4428 4712 4480
rect 4764 4468 4770 4480
rect 5905 4471 5963 4477
rect 5905 4468 5917 4471
rect 4764 4440 5917 4468
rect 4764 4428 4770 4440
rect 5905 4437 5917 4440
rect 5951 4437 5963 4471
rect 7466 4468 7472 4480
rect 7427 4440 7472 4468
rect 5905 4431 5963 4437
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 8220 4468 8248 4508
rect 9186 4505 9198 4508
rect 9232 4505 9244 4539
rect 9186 4499 9244 4505
rect 18230 4496 18236 4548
rect 18288 4536 18294 4548
rect 18325 4539 18383 4545
rect 18325 4536 18337 4539
rect 18288 4508 18337 4536
rect 18288 4496 18294 4508
rect 18325 4505 18337 4508
rect 18371 4536 18383 4539
rect 19536 4536 19564 4635
rect 21634 4632 21640 4644
rect 21692 4632 21698 4684
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 19978 4604 19984 4616
rect 19751 4576 19984 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 18371 4508 19564 4536
rect 18371 4505 18383 4508
rect 18325 4499 18383 4505
rect 10594 4468 10600 4480
rect 8220 4440 10600 4468
rect 10594 4428 10600 4440
rect 10652 4428 10658 4480
rect 11977 4471 12035 4477
rect 11977 4437 11989 4471
rect 12023 4468 12035 4471
rect 12802 4468 12808 4480
rect 12023 4440 12808 4468
rect 12023 4437 12035 4440
rect 11977 4431 12035 4437
rect 12802 4428 12808 4440
rect 12860 4428 12866 4480
rect 18690 4468 18696 4480
rect 18651 4440 18696 4468
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 19242 4468 19248 4480
rect 19203 4440 19248 4468
rect 19242 4428 19248 4440
rect 19300 4428 19306 4480
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 19628 4468 19656 4567
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 20254 4604 20260 4616
rect 20215 4576 20260 4604
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 20441 4607 20499 4613
rect 20441 4573 20453 4607
rect 20487 4604 20499 4607
rect 21545 4607 21603 4613
rect 21545 4604 21557 4607
rect 20487 4576 21557 4604
rect 20487 4573 20499 4576
rect 20441 4567 20499 4573
rect 21545 4573 21557 4576
rect 21591 4573 21603 4607
rect 21545 4567 21603 4573
rect 21729 4607 21787 4613
rect 21729 4573 21741 4607
rect 21775 4604 21787 4607
rect 21818 4604 21824 4616
rect 21775 4576 21824 4604
rect 21775 4573 21787 4576
rect 21729 4567 21787 4573
rect 20070 4496 20076 4548
rect 20128 4536 20134 4548
rect 20456 4536 20484 4567
rect 21818 4564 21824 4576
rect 21876 4604 21882 4616
rect 23198 4604 23204 4616
rect 21876 4576 23204 4604
rect 21876 4564 21882 4576
rect 23198 4564 23204 4576
rect 23256 4564 23262 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4573 24639 4607
rect 24854 4604 24860 4616
rect 24815 4576 24860 4604
rect 24581 4567 24639 4573
rect 20128 4508 20484 4536
rect 24596 4536 24624 4567
rect 24854 4564 24860 4576
rect 24912 4564 24918 4616
rect 25498 4604 25504 4616
rect 25459 4576 25504 4604
rect 25498 4564 25504 4576
rect 25556 4564 25562 4616
rect 25777 4607 25835 4613
rect 25777 4573 25789 4607
rect 25823 4573 25835 4607
rect 26786 4604 26792 4616
rect 25777 4567 25835 4573
rect 26344 4576 26792 4604
rect 25516 4536 25544 4564
rect 24596 4508 25544 4536
rect 20128 4496 20134 4508
rect 20346 4468 20352 4480
rect 19484 4440 20352 4468
rect 19484 4428 19490 4440
rect 20346 4428 20352 4440
rect 20404 4428 20410 4480
rect 20530 4428 20536 4480
rect 20588 4468 20594 4480
rect 23106 4468 23112 4480
rect 20588 4440 23112 4468
rect 20588 4428 20594 4440
rect 23106 4428 23112 4440
rect 23164 4428 23170 4480
rect 24394 4468 24400 4480
rect 24355 4440 24400 4468
rect 24394 4428 24400 4440
rect 24452 4428 24458 4480
rect 24946 4428 24952 4480
rect 25004 4468 25010 4480
rect 25317 4471 25375 4477
rect 25317 4468 25329 4471
rect 25004 4440 25329 4468
rect 25004 4428 25010 4440
rect 25317 4437 25329 4440
rect 25363 4437 25375 4471
rect 25792 4468 25820 4567
rect 26234 4496 26240 4548
rect 26292 4536 26298 4548
rect 26344 4545 26372 4576
rect 26786 4564 26792 4576
rect 26844 4564 26850 4616
rect 27264 4604 27292 4780
rect 27341 4777 27353 4811
rect 27387 4777 27399 4811
rect 27522 4808 27528 4820
rect 27483 4780 27528 4808
rect 27341 4771 27399 4777
rect 27356 4740 27384 4771
rect 27522 4768 27528 4780
rect 27580 4768 27586 4820
rect 41598 4808 41604 4820
rect 29012 4780 41604 4808
rect 28902 4740 28908 4752
rect 27356 4712 28908 4740
rect 28902 4700 28908 4712
rect 28960 4700 28966 4752
rect 29012 4604 29040 4780
rect 41598 4768 41604 4780
rect 41656 4768 41662 4820
rect 41690 4768 41696 4820
rect 41748 4808 41754 4820
rect 42521 4811 42579 4817
rect 42521 4808 42533 4811
rect 41748 4780 42533 4808
rect 41748 4768 41754 4780
rect 42521 4777 42533 4780
rect 42567 4777 42579 4811
rect 42521 4771 42579 4777
rect 42794 4768 42800 4820
rect 42852 4808 42858 4820
rect 43441 4811 43499 4817
rect 43441 4808 43453 4811
rect 42852 4780 43453 4808
rect 42852 4768 42858 4780
rect 43441 4777 43453 4780
rect 43487 4777 43499 4811
rect 46474 4808 46480 4820
rect 46435 4780 46480 4808
rect 43441 4771 43499 4777
rect 46474 4768 46480 4780
rect 46532 4768 46538 4820
rect 47305 4743 47363 4749
rect 47305 4740 47317 4743
rect 31726 4712 47317 4740
rect 29086 4632 29092 4684
rect 29144 4672 29150 4684
rect 31726 4672 31754 4712
rect 47305 4709 47317 4712
rect 47351 4709 47363 4743
rect 47305 4703 47363 4709
rect 29144 4644 31754 4672
rect 29144 4632 29150 4644
rect 34514 4632 34520 4684
rect 34572 4672 34578 4684
rect 40586 4672 40592 4684
rect 34572 4644 40592 4672
rect 34572 4632 34578 4644
rect 40586 4632 40592 4644
rect 40644 4632 40650 4684
rect 40865 4675 40923 4681
rect 40865 4672 40877 4675
rect 40696 4644 40877 4672
rect 27264 4576 29040 4604
rect 32033 4607 32091 4613
rect 32033 4573 32045 4607
rect 32079 4604 32091 4607
rect 32122 4604 32128 4616
rect 32079 4576 32128 4604
rect 32079 4573 32091 4576
rect 32033 4567 32091 4573
rect 32122 4564 32128 4576
rect 32180 4564 32186 4616
rect 32306 4604 32312 4616
rect 32267 4576 32312 4604
rect 32306 4564 32312 4576
rect 32364 4564 32370 4616
rect 32401 4607 32459 4613
rect 32401 4573 32413 4607
rect 32447 4604 32459 4607
rect 32950 4604 32956 4616
rect 32447 4576 32956 4604
rect 32447 4573 32459 4576
rect 32401 4567 32459 4573
rect 32950 4564 32956 4576
rect 33008 4564 33014 4616
rect 35618 4604 35624 4616
rect 35579 4576 35624 4604
rect 35618 4564 35624 4576
rect 35676 4564 35682 4616
rect 35714 4607 35772 4613
rect 35714 4573 35726 4607
rect 35760 4573 35772 4607
rect 35986 4604 35992 4616
rect 35947 4576 35992 4604
rect 35714 4567 35772 4573
rect 26329 4539 26387 4545
rect 26329 4536 26341 4539
rect 26292 4508 26341 4536
rect 26292 4496 26298 4508
rect 26329 4505 26341 4508
rect 26375 4505 26387 4539
rect 26329 4499 26387 4505
rect 26545 4539 26603 4545
rect 26545 4505 26557 4539
rect 26591 4536 26603 4539
rect 27157 4539 27215 4545
rect 26591 4508 27108 4536
rect 26591 4505 26603 4508
rect 26545 4499 26603 4505
rect 26697 4471 26755 4477
rect 26697 4468 26709 4471
rect 25792 4440 26709 4468
rect 25317 4431 25375 4437
rect 26697 4437 26709 4440
rect 26743 4437 26755 4471
rect 27080 4468 27108 4508
rect 27157 4505 27169 4539
rect 27203 4536 27215 4539
rect 27982 4536 27988 4548
rect 27203 4508 27988 4536
rect 27203 4505 27215 4508
rect 27157 4499 27215 4505
rect 27982 4496 27988 4508
rect 28040 4496 28046 4548
rect 32217 4539 32275 4545
rect 32217 4505 32229 4539
rect 32263 4536 32275 4539
rect 32490 4536 32496 4548
rect 32263 4508 32496 4536
rect 32263 4505 32275 4508
rect 32217 4499 32275 4505
rect 32490 4496 32496 4508
rect 32548 4496 32554 4548
rect 35434 4496 35440 4548
rect 35492 4536 35498 4548
rect 35729 4536 35757 4567
rect 35986 4564 35992 4576
rect 36044 4564 36050 4616
rect 36170 4613 36176 4616
rect 36127 4607 36176 4613
rect 36127 4604 36139 4607
rect 36083 4576 36139 4604
rect 36127 4573 36139 4576
rect 36173 4573 36176 4607
rect 36127 4567 36176 4573
rect 36170 4564 36176 4567
rect 36228 4604 36234 4616
rect 36722 4604 36728 4616
rect 36228 4576 36728 4604
rect 36228 4564 36234 4576
rect 36722 4564 36728 4576
rect 36780 4604 36786 4616
rect 36817 4607 36875 4613
rect 36817 4604 36829 4607
rect 36780 4576 36829 4604
rect 36780 4564 36786 4576
rect 36817 4573 36829 4576
rect 36863 4573 36875 4607
rect 36998 4604 37004 4616
rect 36959 4576 37004 4604
rect 36817 4567 36875 4573
rect 36998 4564 37004 4576
rect 37056 4564 37062 4616
rect 37550 4564 37556 4616
rect 37608 4604 37614 4616
rect 38197 4607 38255 4613
rect 38197 4604 38209 4607
rect 37608 4576 38209 4604
rect 37608 4564 37614 4576
rect 38197 4573 38209 4576
rect 38243 4604 38255 4607
rect 38562 4604 38568 4616
rect 38243 4576 38568 4604
rect 38243 4573 38255 4576
rect 38197 4567 38255 4573
rect 38562 4564 38568 4576
rect 38620 4564 38626 4616
rect 40034 4564 40040 4616
rect 40092 4604 40098 4616
rect 40696 4604 40724 4644
rect 40865 4641 40877 4644
rect 40911 4672 40923 4675
rect 40911 4644 46934 4672
rect 40911 4641 40923 4644
rect 40865 4635 40923 4641
rect 42352 4613 42380 4644
rect 40092 4576 40724 4604
rect 42337 4607 42395 4613
rect 40092 4564 40098 4576
rect 42337 4573 42349 4607
rect 42383 4573 42395 4607
rect 42337 4567 42395 4573
rect 42613 4607 42671 4613
rect 42613 4573 42625 4607
rect 42659 4604 42671 4607
rect 42978 4604 42984 4616
rect 42659 4576 42984 4604
rect 42659 4573 42671 4576
rect 42613 4567 42671 4573
rect 42978 4564 42984 4576
rect 43036 4564 43042 4616
rect 43272 4613 43300 4644
rect 43257 4607 43315 4613
rect 43257 4573 43269 4607
rect 43303 4573 43315 4607
rect 43257 4567 43315 4573
rect 43530 4564 43536 4616
rect 43588 4604 43594 4616
rect 43588 4576 43633 4604
rect 43588 4564 43594 4576
rect 44910 4564 44916 4616
rect 44968 4604 44974 4616
rect 45925 4607 45983 4613
rect 45925 4604 45937 4607
rect 44968 4576 45937 4604
rect 44968 4564 44974 4576
rect 45925 4573 45937 4576
rect 45971 4573 45983 4607
rect 46106 4604 46112 4616
rect 45925 4567 45983 4573
rect 46032 4576 46112 4604
rect 35492 4508 35757 4536
rect 35897 4539 35955 4545
rect 35492 4496 35498 4508
rect 35897 4505 35909 4539
rect 35943 4505 35955 4539
rect 36446 4536 36452 4548
rect 35897 4499 35955 4505
rect 36142 4508 36452 4536
rect 27357 4471 27415 4477
rect 27357 4468 27369 4471
rect 27080 4440 27369 4468
rect 26697 4431 26755 4437
rect 27357 4437 27369 4440
rect 27403 4468 27415 4471
rect 31294 4468 31300 4480
rect 27403 4440 31300 4468
rect 27403 4437 27415 4440
rect 27357 4431 27415 4437
rect 31294 4428 31300 4440
rect 31352 4428 31358 4480
rect 32582 4468 32588 4480
rect 32543 4440 32588 4468
rect 32582 4428 32588 4440
rect 32640 4428 32646 4480
rect 35912 4468 35940 4499
rect 36142 4468 36170 4508
rect 36446 4496 36452 4508
rect 36504 4496 36510 4548
rect 37016 4536 37044 4564
rect 39022 4536 39028 4548
rect 37016 4508 39028 4536
rect 39022 4496 39028 4508
rect 39080 4496 39086 4548
rect 40126 4496 40132 4548
rect 40184 4536 40190 4548
rect 40678 4536 40684 4548
rect 40184 4508 40684 4536
rect 40184 4496 40190 4508
rect 40678 4496 40684 4508
rect 40736 4496 40742 4548
rect 46032 4536 46060 4576
rect 46106 4564 46112 4576
rect 46164 4604 46170 4616
rect 46293 4607 46351 4613
rect 46164 4576 46257 4604
rect 46164 4564 46170 4576
rect 46293 4573 46305 4607
rect 46339 4604 46351 4607
rect 46382 4604 46388 4616
rect 46339 4576 46388 4604
rect 46339 4573 46351 4576
rect 46293 4567 46351 4573
rect 46382 4564 46388 4576
rect 46440 4564 46446 4616
rect 46906 4604 46934 4644
rect 47118 4604 47124 4616
rect 46906 4576 47124 4604
rect 47118 4564 47124 4576
rect 47176 4564 47182 4616
rect 47394 4564 47400 4616
rect 47452 4604 47458 4616
rect 48222 4604 48228 4616
rect 47452 4576 47497 4604
rect 48183 4576 48228 4604
rect 47452 4564 47458 4576
rect 48222 4564 48228 4576
rect 48280 4564 48286 4616
rect 46198 4536 46204 4548
rect 41616 4508 46060 4536
rect 46159 4508 46204 4536
rect 36262 4468 36268 4480
rect 35912 4440 36170 4468
rect 36223 4440 36268 4468
rect 36262 4428 36268 4440
rect 36320 4428 36326 4480
rect 38286 4468 38292 4480
rect 38247 4440 38292 4468
rect 38286 4428 38292 4440
rect 38344 4428 38350 4480
rect 40218 4428 40224 4480
rect 40276 4468 40282 4480
rect 41616 4468 41644 4508
rect 46198 4496 46204 4508
rect 46256 4496 46262 4548
rect 46937 4539 46995 4545
rect 46937 4505 46949 4539
rect 46983 4536 46995 4539
rect 48470 4539 48528 4545
rect 48470 4536 48482 4539
rect 46983 4508 48482 4536
rect 46983 4505 46995 4508
rect 46937 4499 46995 4505
rect 48470 4505 48482 4508
rect 48516 4505 48528 4539
rect 48470 4499 48528 4505
rect 40276 4440 41644 4468
rect 42153 4471 42211 4477
rect 40276 4428 40282 4440
rect 42153 4437 42165 4471
rect 42199 4468 42211 4471
rect 42242 4468 42248 4480
rect 42199 4440 42248 4468
rect 42199 4437 42211 4440
rect 42153 4431 42211 4437
rect 42242 4428 42248 4440
rect 42300 4428 42306 4480
rect 43073 4471 43131 4477
rect 43073 4437 43085 4471
rect 43119 4468 43131 4471
rect 45370 4468 45376 4480
rect 43119 4440 45376 4468
rect 43119 4437 43131 4440
rect 43073 4431 43131 4437
rect 45370 4428 45376 4440
rect 45428 4428 45434 4480
rect 46842 4428 46848 4480
rect 46900 4468 46906 4480
rect 49605 4471 49663 4477
rect 49605 4468 49617 4471
rect 46900 4440 49617 4468
rect 46900 4428 46906 4440
rect 49605 4437 49617 4440
rect 49651 4437 49663 4471
rect 49605 4431 49663 4437
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 2130 4224 2136 4276
rect 2188 4264 2194 4276
rect 20530 4264 20536 4276
rect 2188 4236 20536 4264
rect 2188 4224 2194 4236
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 24854 4224 24860 4276
rect 24912 4264 24918 4276
rect 32582 4264 32588 4276
rect 24912 4236 32588 4264
rect 24912 4224 24918 4236
rect 32582 4224 32588 4236
rect 32640 4224 32646 4276
rect 35802 4224 35808 4276
rect 35860 4224 35866 4276
rect 37550 4264 37556 4276
rect 36004 4236 37556 4264
rect 8662 4156 8668 4208
rect 8720 4196 8726 4208
rect 9950 4196 9956 4208
rect 8720 4168 9956 4196
rect 8720 4156 8726 4168
rect 9950 4156 9956 4168
rect 10008 4156 10014 4208
rect 19334 4196 19340 4208
rect 11440 4168 12020 4196
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 1443 4100 2084 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 198 3884 204 3936
rect 256 3924 262 3936
rect 1581 3927 1639 3933
rect 1581 3924 1593 3927
rect 256 3896 1593 3924
rect 256 3884 262 3896
rect 1581 3893 1593 3896
rect 1627 3893 1639 3927
rect 2056 3924 2084 4100
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2400 4131 2458 4137
rect 2188 4100 2233 4128
rect 2188 4088 2194 4100
rect 2400 4097 2412 4131
rect 2446 4128 2458 4131
rect 3418 4128 3424 4140
rect 2446 4100 3424 4128
rect 2446 4097 2458 4100
rect 2400 4091 2458 4097
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4128 4215 4131
rect 4706 4128 4712 4140
rect 4203 4100 4712 4128
rect 4203 4097 4215 4100
rect 4157 4091 4215 4097
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 4798 4088 4804 4140
rect 4856 4128 4862 4140
rect 4856 4100 4901 4128
rect 4856 4088 4862 4100
rect 5074 4088 5080 4140
rect 5132 4128 5138 4140
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 5132 4100 5641 4128
rect 5132 4088 5138 4100
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 6564 4060 6592 4091
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 8067 4131 8125 4137
rect 8067 4128 8079 4131
rect 7524 4100 8079 4128
rect 7524 4088 7530 4100
rect 8067 4097 8079 4100
rect 8113 4097 8125 4131
rect 8202 4128 8208 4140
rect 8163 4100 8208 4128
rect 8067 4091 8125 4097
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8318 4131 8376 4137
rect 8318 4097 8330 4131
rect 8364 4128 8376 4131
rect 8364 4100 8432 4128
rect 8364 4097 8376 4100
rect 8318 4091 8376 4097
rect 7834 4060 7840 4072
rect 4120 4032 6592 4060
rect 7795 4032 7840 4060
rect 4120 4020 4126 4032
rect 7834 4020 7840 4032
rect 7892 4020 7898 4072
rect 8404 4060 8432 4100
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 8536 4100 8581 4128
rect 8536 4088 8542 4100
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9456 4100 9996 4128
rect 9456 4088 9462 4100
rect 9858 4060 9864 4072
rect 8404 4032 9864 4060
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 9968 4060 9996 4100
rect 10410 4088 10416 4140
rect 10468 4128 10474 4140
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 10468 4100 10701 4128
rect 10468 4088 10474 4100
rect 10689 4097 10701 4100
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 11440 4060 11468 4168
rect 11517 4131 11575 4137
rect 11517 4097 11529 4131
rect 11563 4128 11575 4131
rect 11882 4128 11888 4140
rect 11563 4100 11888 4128
rect 11563 4097 11575 4100
rect 11517 4091 11575 4097
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 11992 4128 12020 4168
rect 18064 4168 19340 4196
rect 16390 4128 16396 4140
rect 11992 4100 16396 4128
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4128 16727 4131
rect 18064 4128 18092 4168
rect 19334 4156 19340 4168
rect 19392 4156 19398 4208
rect 28528 4199 28586 4205
rect 28528 4165 28540 4199
rect 28574 4196 28586 4199
rect 28626 4196 28632 4208
rect 28574 4168 28632 4196
rect 28574 4165 28586 4168
rect 28528 4159 28586 4165
rect 28626 4156 28632 4168
rect 28684 4156 28690 4208
rect 35526 4196 35532 4208
rect 34983 4168 35532 4196
rect 18230 4128 18236 4140
rect 16715 4100 18092 4128
rect 18191 4100 18236 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 18417 4131 18475 4137
rect 18417 4097 18429 4131
rect 18463 4128 18475 4131
rect 18506 4128 18512 4140
rect 18463 4100 18512 4128
rect 18463 4097 18475 4100
rect 18417 4091 18475 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18690 4088 18696 4140
rect 18748 4128 18754 4140
rect 19153 4131 19211 4137
rect 19153 4128 19165 4131
rect 18748 4100 19165 4128
rect 18748 4088 18754 4100
rect 19153 4097 19165 4100
rect 19199 4097 19211 4131
rect 19426 4126 19432 4140
rect 19153 4091 19211 4097
rect 19260 4098 19432 4126
rect 11790 4060 11796 4072
rect 9968 4032 11468 4060
rect 11751 4032 11796 4060
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 15013 4063 15071 4069
rect 15013 4060 15025 4063
rect 13504 4032 15025 4060
rect 13504 4020 13510 4032
rect 15013 4029 15025 4032
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 15194 4020 15200 4072
rect 15252 4060 15258 4072
rect 15289 4063 15347 4069
rect 15289 4060 15301 4063
rect 15252 4032 15301 4060
rect 15252 4020 15258 4032
rect 15289 4029 15301 4032
rect 15335 4029 15347 4063
rect 15289 4023 15347 4029
rect 16022 4020 16028 4072
rect 16080 4060 16086 4072
rect 19260 4069 19288 4098
rect 19426 4088 19432 4098
rect 19484 4088 19490 4140
rect 22002 4128 22008 4140
rect 21963 4100 22008 4128
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 33134 4128 33140 4140
rect 27356 4100 33140 4128
rect 16945 4063 17003 4069
rect 16945 4060 16957 4063
rect 16080 4032 16957 4060
rect 16080 4020 16086 4032
rect 16945 4029 16957 4032
rect 16991 4029 17003 4063
rect 16945 4023 17003 4029
rect 18325 4063 18383 4069
rect 18325 4029 18337 4063
rect 18371 4060 18383 4063
rect 19061 4063 19119 4069
rect 19061 4060 19073 4063
rect 18371 4032 19073 4060
rect 18371 4029 18383 4032
rect 18325 4023 18383 4029
rect 19061 4029 19073 4032
rect 19107 4029 19119 4063
rect 19061 4023 19119 4029
rect 19245 4063 19303 4069
rect 19245 4029 19257 4063
rect 19291 4029 19303 4063
rect 19245 4023 19303 4029
rect 19337 4063 19395 4069
rect 19337 4029 19349 4063
rect 19383 4060 19395 4063
rect 20162 4060 20168 4072
rect 19383 4032 20168 4060
rect 19383 4029 19395 4032
rect 19337 4023 19395 4029
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 20254 4020 20260 4072
rect 20312 4060 20318 4072
rect 27356 4060 27384 4100
rect 33134 4088 33140 4100
rect 33192 4088 33198 4140
rect 33502 4088 33508 4140
rect 33560 4128 33566 4140
rect 34514 4128 34520 4140
rect 33560 4100 34520 4128
rect 33560 4088 33566 4100
rect 34514 4088 34520 4100
rect 34572 4088 34578 4140
rect 34698 4128 34704 4140
rect 34659 4100 34704 4128
rect 34698 4088 34704 4100
rect 34756 4088 34762 4140
rect 34885 4131 34943 4137
rect 34885 4097 34897 4131
rect 34931 4126 34943 4131
rect 34983 4126 35011 4168
rect 35526 4156 35532 4168
rect 35584 4156 35590 4208
rect 34931 4098 35011 4126
rect 35069 4131 35127 4137
rect 34931 4097 34943 4098
rect 34885 4091 34943 4097
rect 35069 4097 35081 4131
rect 35115 4097 35127 4131
rect 35069 4091 35127 4097
rect 20312 4032 27384 4060
rect 20312 4020 20318 4032
rect 28258 4020 28264 4072
rect 28316 4060 28322 4072
rect 28316 4032 28361 4060
rect 28316 4020 28322 4032
rect 33686 4020 33692 4072
rect 33744 4060 33750 4072
rect 34716 4060 34744 4088
rect 33744 4032 34744 4060
rect 34793 4063 34851 4069
rect 33744 4020 33750 4032
rect 34793 4029 34805 4063
rect 34839 4029 34851 4063
rect 35084 4060 35112 4091
rect 35618 4088 35624 4140
rect 35676 4128 35682 4140
rect 35820 4137 35848 4224
rect 36004 4205 36032 4236
rect 37550 4224 37556 4236
rect 37608 4224 37614 4276
rect 39022 4224 39028 4276
rect 39080 4264 39086 4276
rect 40954 4264 40960 4276
rect 39080 4236 40960 4264
rect 39080 4224 39086 4236
rect 40954 4224 40960 4236
rect 41012 4224 41018 4276
rect 41046 4224 41052 4276
rect 41104 4264 41110 4276
rect 42794 4264 42800 4276
rect 42852 4273 42858 4276
rect 42852 4267 42871 4273
rect 41104 4236 42800 4264
rect 41104 4224 41110 4236
rect 42794 4224 42800 4236
rect 42859 4233 42871 4267
rect 42978 4264 42984 4276
rect 42939 4236 42984 4264
rect 42852 4227 42871 4233
rect 42852 4224 42858 4227
rect 42978 4224 42984 4236
rect 43036 4224 43042 4276
rect 43530 4224 43536 4276
rect 43588 4264 43594 4276
rect 43809 4267 43867 4273
rect 43809 4264 43821 4267
rect 43588 4236 43821 4264
rect 43588 4224 43594 4236
rect 43809 4233 43821 4236
rect 43855 4233 43867 4267
rect 43809 4227 43867 4233
rect 35989 4199 36047 4205
rect 35989 4165 36001 4199
rect 36035 4165 36047 4199
rect 35989 4159 36047 4165
rect 36538 4156 36544 4208
rect 36596 4196 36602 4208
rect 42613 4199 42671 4205
rect 36596 4168 42564 4196
rect 36596 4156 36602 4168
rect 35713 4131 35771 4137
rect 35713 4128 35725 4131
rect 35676 4100 35725 4128
rect 35676 4088 35682 4100
rect 35713 4097 35725 4100
rect 35759 4097 35771 4131
rect 35713 4091 35771 4097
rect 35806 4131 35864 4137
rect 35806 4097 35818 4131
rect 35852 4097 35864 4131
rect 35806 4091 35864 4097
rect 36081 4131 36139 4137
rect 36081 4097 36093 4131
rect 36127 4097 36139 4131
rect 36081 4091 36139 4097
rect 35434 4060 35440 4072
rect 35084 4032 35440 4060
rect 34793 4023 34851 4029
rect 4614 3992 4620 4004
rect 3436 3964 4620 3992
rect 3436 3924 3464 3964
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 6270 3992 6276 4004
rect 4724 3964 6276 3992
rect 2056 3896 3464 3924
rect 3513 3927 3571 3933
rect 1581 3887 1639 3893
rect 3513 3893 3525 3927
rect 3559 3924 3571 3927
rect 3602 3924 3608 3936
rect 3559 3896 3608 3924
rect 3559 3893 3571 3896
rect 3513 3887 3571 3893
rect 3602 3884 3608 3896
rect 3660 3884 3666 3936
rect 4065 3927 4123 3933
rect 4065 3893 4077 3927
rect 4111 3924 4123 3927
rect 4724 3924 4752 3964
rect 6270 3952 6276 3964
rect 6328 3952 6334 4004
rect 6365 3995 6423 4001
rect 6365 3961 6377 3995
rect 6411 3992 6423 3995
rect 7466 3992 7472 4004
rect 6411 3964 7472 3992
rect 6411 3961 6423 3964
rect 6365 3955 6423 3961
rect 7466 3952 7472 3964
rect 7524 3952 7530 4004
rect 7558 3952 7564 4004
rect 7616 3992 7622 4004
rect 27246 3992 27252 4004
rect 7616 3964 27252 3992
rect 7616 3952 7622 3964
rect 27246 3952 27252 3964
rect 27304 3952 27310 4004
rect 29380 3964 29960 3992
rect 4111 3896 4752 3924
rect 5445 3927 5503 3933
rect 4111 3893 4123 3896
rect 4065 3887 4123 3893
rect 5445 3893 5457 3927
rect 5491 3924 5503 3927
rect 6546 3924 6552 3936
rect 5491 3896 6552 3924
rect 5491 3893 5503 3896
rect 5445 3887 5503 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 9214 3924 9220 3936
rect 6696 3896 9220 3924
rect 6696 3884 6702 3896
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 13446 3924 13452 3936
rect 10551 3896 13452 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 13998 3884 14004 3936
rect 14056 3924 14062 3936
rect 18782 3924 18788 3936
rect 14056 3896 18788 3924
rect 14056 3884 14062 3896
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 18877 3927 18935 3933
rect 18877 3893 18889 3927
rect 18923 3924 18935 3927
rect 19426 3924 19432 3936
rect 18923 3896 19432 3924
rect 18923 3893 18935 3896
rect 18877 3887 18935 3893
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 21542 3924 21548 3936
rect 19576 3896 21548 3924
rect 19576 3884 19582 3896
rect 21542 3884 21548 3896
rect 21600 3884 21606 3936
rect 21821 3927 21879 3933
rect 21821 3893 21833 3927
rect 21867 3924 21879 3927
rect 22646 3924 22652 3936
rect 21867 3896 22652 3924
rect 21867 3893 21879 3896
rect 21821 3887 21879 3893
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 23474 3884 23480 3936
rect 23532 3924 23538 3936
rect 28166 3924 28172 3936
rect 23532 3896 28172 3924
rect 23532 3884 23538 3896
rect 28166 3884 28172 3896
rect 28224 3884 28230 3936
rect 28442 3884 28448 3936
rect 28500 3924 28506 3936
rect 29380 3924 29408 3964
rect 28500 3896 29408 3924
rect 28500 3884 28506 3896
rect 29454 3884 29460 3936
rect 29512 3924 29518 3936
rect 29641 3927 29699 3933
rect 29641 3924 29653 3927
rect 29512 3896 29653 3924
rect 29512 3884 29518 3896
rect 29641 3893 29653 3896
rect 29687 3893 29699 3927
rect 29932 3924 29960 3964
rect 30006 3952 30012 4004
rect 30064 3992 30070 4004
rect 33410 3992 33416 4004
rect 30064 3964 33416 3992
rect 30064 3952 30070 3964
rect 33410 3952 33416 3964
rect 33468 3952 33474 4004
rect 34808 3992 34836 4023
rect 35434 4020 35440 4032
rect 35492 4020 35498 4072
rect 36096 3992 36124 4091
rect 36170 4088 36176 4140
rect 36228 4137 36234 4140
rect 36228 4128 36236 4137
rect 38470 4128 38476 4140
rect 36228 4100 36273 4128
rect 38431 4100 38476 4128
rect 36228 4091 36236 4100
rect 36228 4088 36234 4091
rect 38470 4088 38476 4100
rect 38528 4088 38534 4140
rect 38566 4131 38624 4137
rect 38566 4097 38578 4131
rect 38612 4097 38624 4131
rect 38566 4091 38624 4097
rect 34624 3964 36124 3992
rect 31570 3924 31576 3936
rect 29932 3896 31576 3924
rect 29641 3887 29699 3893
rect 31570 3884 31576 3896
rect 31628 3924 31634 3936
rect 34624 3924 34652 3964
rect 37366 3952 37372 4004
rect 37424 3992 37430 4004
rect 38580 3992 38608 4091
rect 38654 4088 38660 4140
rect 38712 4128 38718 4140
rect 38749 4131 38807 4137
rect 38749 4128 38761 4131
rect 38712 4100 38761 4128
rect 38712 4088 38718 4100
rect 38749 4097 38761 4100
rect 38795 4097 38807 4131
rect 38749 4091 38807 4097
rect 38838 4088 38844 4140
rect 38896 4128 38902 4140
rect 39022 4137 39028 4140
rect 38979 4131 39028 4137
rect 38896 4100 38941 4128
rect 38896 4088 38902 4100
rect 38979 4097 38991 4131
rect 39025 4097 39028 4131
rect 38979 4091 39028 4097
rect 39022 4088 39028 4091
rect 39080 4088 39086 4140
rect 40037 4131 40095 4137
rect 40037 4097 40049 4131
rect 40083 4128 40095 4131
rect 40218 4128 40224 4140
rect 40083 4100 40224 4128
rect 40083 4097 40095 4100
rect 40037 4091 40095 4097
rect 40218 4088 40224 4100
rect 40276 4088 40282 4140
rect 40586 4088 40592 4140
rect 40644 4128 40650 4140
rect 41046 4128 41052 4140
rect 40644 4100 41052 4128
rect 40644 4088 40650 4100
rect 41046 4088 41052 4100
rect 41104 4088 41110 4140
rect 41233 4131 41291 4137
rect 41233 4097 41245 4131
rect 41279 4128 41291 4131
rect 41322 4128 41328 4140
rect 41279 4100 41328 4128
rect 41279 4097 41291 4100
rect 41233 4091 41291 4097
rect 41322 4088 41328 4100
rect 41380 4088 41386 4140
rect 42536 4060 42564 4168
rect 42613 4165 42625 4199
rect 42659 4165 42671 4199
rect 42613 4159 42671 4165
rect 42628 4128 42656 4159
rect 42702 4156 42708 4208
rect 42760 4196 42766 4208
rect 43441 4199 43499 4205
rect 43441 4196 43453 4199
rect 42760 4156 42774 4196
rect 42746 4128 42774 4156
rect 42628 4100 42774 4128
rect 42812 4168 43453 4196
rect 42812 4060 42840 4168
rect 43441 4165 43453 4168
rect 43487 4165 43499 4199
rect 46106 4196 46112 4208
rect 43441 4159 43499 4165
rect 43671 4165 43729 4171
rect 46067 4168 46112 4196
rect 43671 4162 43683 4165
rect 43661 4131 43683 4162
rect 43717 4131 43729 4165
rect 46106 4156 46112 4168
rect 46164 4156 46170 4208
rect 46842 4196 46848 4208
rect 46216 4168 46848 4196
rect 43661 4125 43729 4131
rect 45922 4128 45928 4140
rect 42536 4032 42840 4060
rect 37424 3964 38608 3992
rect 42812 3992 42840 4032
rect 42886 4020 42892 4072
rect 42944 4060 42950 4072
rect 43661 4060 43689 4125
rect 45883 4100 45928 4128
rect 45922 4088 45928 4100
rect 45980 4088 45986 4140
rect 46014 4088 46020 4140
rect 46072 4128 46078 4140
rect 46216 4137 46244 4168
rect 46842 4156 46848 4168
rect 46900 4156 46906 4208
rect 46934 4156 46940 4208
rect 46992 4196 46998 4208
rect 48222 4196 48228 4208
rect 46992 4168 48228 4196
rect 46992 4156 46998 4168
rect 48222 4156 48228 4168
rect 48280 4156 48286 4208
rect 46201 4131 46259 4137
rect 46201 4128 46213 4131
rect 46072 4100 46213 4128
rect 46072 4088 46078 4100
rect 46201 4097 46213 4100
rect 46247 4097 46259 4131
rect 46201 4091 46259 4097
rect 46290 4088 46296 4140
rect 46348 4128 46354 4140
rect 46348 4100 46441 4128
rect 46348 4088 46354 4100
rect 46474 4088 46480 4140
rect 46532 4128 46538 4140
rect 46952 4128 46980 4156
rect 46532 4100 46980 4128
rect 46532 4088 46538 4100
rect 42944 4032 43689 4060
rect 42944 4020 42950 4032
rect 45462 4020 45468 4072
rect 45520 4060 45526 4072
rect 46308 4060 46336 4088
rect 45520 4032 46336 4060
rect 45520 4020 45526 4032
rect 45830 3992 45836 4004
rect 42812 3964 45836 3992
rect 37424 3952 37430 3964
rect 45830 3952 45836 3964
rect 45888 3952 45894 4004
rect 46477 3995 46535 4001
rect 46477 3961 46489 3995
rect 46523 3992 46535 3995
rect 47394 3992 47400 4004
rect 46523 3964 47400 3992
rect 46523 3961 46535 3964
rect 46477 3955 46535 3961
rect 47394 3952 47400 3964
rect 47452 3952 47458 4004
rect 31628 3896 34652 3924
rect 31628 3884 31634 3896
rect 34698 3884 34704 3936
rect 34756 3924 34762 3936
rect 35253 3927 35311 3933
rect 35253 3924 35265 3927
rect 34756 3896 35265 3924
rect 34756 3884 34762 3896
rect 35253 3893 35265 3896
rect 35299 3893 35311 3927
rect 36354 3924 36360 3936
rect 36315 3896 36360 3924
rect 35253 3887 35311 3893
rect 36354 3884 36360 3896
rect 36412 3884 36418 3936
rect 39114 3924 39120 3936
rect 39075 3896 39120 3924
rect 39114 3884 39120 3896
rect 39172 3884 39178 3936
rect 39850 3924 39856 3936
rect 39811 3896 39856 3924
rect 39850 3884 39856 3896
rect 39908 3884 39914 3936
rect 41138 3884 41144 3936
rect 41196 3924 41202 3936
rect 41417 3927 41475 3933
rect 41417 3924 41429 3927
rect 41196 3896 41429 3924
rect 41196 3884 41202 3896
rect 41417 3893 41429 3896
rect 41463 3893 41475 3927
rect 41417 3887 41475 3893
rect 42610 3884 42616 3936
rect 42668 3924 42674 3936
rect 42797 3927 42855 3933
rect 42797 3924 42809 3927
rect 42668 3896 42809 3924
rect 42668 3884 42674 3896
rect 42797 3893 42809 3896
rect 42843 3924 42855 3927
rect 43625 3927 43683 3933
rect 43625 3924 43637 3927
rect 42843 3896 43637 3924
rect 42843 3893 42855 3896
rect 42797 3887 42855 3893
rect 43625 3893 43637 3896
rect 43671 3893 43683 3927
rect 43625 3887 43683 3893
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 2130 3680 2136 3732
rect 2188 3720 2194 3732
rect 4798 3720 4804 3732
rect 2188 3692 4804 3720
rect 2188 3680 2194 3692
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 7558 3720 7564 3732
rect 5040 3692 7564 3720
rect 5040 3680 5046 3692
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8202 3720 8208 3732
rect 7668 3692 8208 3720
rect 4890 3652 4896 3664
rect 4448 3624 4896 3652
rect 4448 3593 4476 3624
rect 4890 3612 4896 3624
rect 4948 3612 4954 3664
rect 7668 3652 7696 3692
rect 8202 3680 8208 3692
rect 8260 3720 8266 3732
rect 11146 3720 11152 3732
rect 8260 3692 11152 3720
rect 8260 3680 8266 3692
rect 11146 3680 11152 3692
rect 11204 3720 11210 3732
rect 11790 3720 11796 3732
rect 11204 3692 11796 3720
rect 11204 3680 11210 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12066 3680 12072 3732
rect 12124 3720 12130 3732
rect 21910 3720 21916 3732
rect 12124 3692 21916 3720
rect 12124 3680 12130 3692
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 22066 3692 27200 3720
rect 7300 3624 7696 3652
rect 7929 3655 7987 3661
rect 4433 3587 4491 3593
rect 3620 3556 4108 3584
rect 1854 3516 1860 3528
rect 1815 3488 1860 3516
rect 1854 3476 1860 3488
rect 1912 3476 1918 3528
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 3510 3516 3516 3528
rect 2731 3488 3516 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 2225 3451 2283 3457
rect 2225 3417 2237 3451
rect 2271 3448 2283 3451
rect 3620 3448 3648 3556
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3936 3488 3985 3516
rect 3936 3476 3942 3488
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 4080 3516 4108 3556
rect 4433 3553 4445 3587
rect 4479 3553 4491 3587
rect 4801 3587 4859 3593
rect 4433 3547 4491 3553
rect 4540 3556 4752 3584
rect 4540 3516 4568 3556
rect 4080 3488 4568 3516
rect 4617 3519 4675 3525
rect 3973 3479 4031 3485
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4724 3516 4752 3556
rect 4801 3553 4813 3587
rect 4847 3584 4859 3587
rect 5074 3584 5080 3596
rect 4847 3556 5080 3584
rect 4847 3553 4859 3556
rect 4801 3547 4859 3553
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 5258 3584 5264 3596
rect 5219 3556 5264 3584
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6788 3556 7113 3584
rect 6788 3544 6794 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 7101 3547 7159 3553
rect 6914 3516 6920 3528
rect 4724 3488 6920 3516
rect 4617 3479 4675 3485
rect 2271 3420 3648 3448
rect 2271 3417 2283 3420
rect 2225 3411 2283 3417
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 4632 3448 4660 3479
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7300 3525 7328 3624
rect 7929 3621 7941 3655
rect 7975 3652 7987 3655
rect 13357 3655 13415 3661
rect 7975 3624 12434 3652
rect 7975 3621 7987 3624
rect 7929 3615 7987 3621
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 9916 3556 10364 3584
rect 9916 3544 9922 3556
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3485 7343 3519
rect 7466 3516 7472 3528
rect 7427 3488 7472 3516
rect 7285 3479 7343 3485
rect 3752 3420 4660 3448
rect 3752 3408 3758 3420
rect 658 3340 664 3392
rect 716 3380 722 3392
rect 2869 3383 2927 3389
rect 2869 3380 2881 3383
rect 716 3352 2881 3380
rect 716 3340 722 3352
rect 2869 3349 2881 3352
rect 2915 3349 2927 3383
rect 3786 3380 3792 3392
rect 3747 3352 3792 3380
rect 2869 3343 2927 3349
rect 3786 3340 3792 3352
rect 3844 3340 3850 3392
rect 4632 3380 4660 3420
rect 5528 3451 5586 3457
rect 5528 3417 5540 3451
rect 5574 3448 5586 3451
rect 6362 3448 6368 3460
rect 5574 3420 6368 3448
rect 5574 3417 5586 3420
rect 5528 3411 5586 3417
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 7300 3448 7328 3479
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7558 3476 7564 3528
rect 7616 3516 7622 3528
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 7616 3488 8125 3516
rect 7616 3476 7622 3488
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3516 10103 3519
rect 10226 3516 10232 3528
rect 10091 3488 10232 3516
rect 10091 3485 10103 3488
rect 10045 3479 10103 3485
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10336 3525 10364 3556
rect 10428 3556 11284 3584
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 10428 3448 10456 3556
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 10594 3516 10600 3528
rect 10551 3488 10600 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 10744 3488 10977 3516
rect 10744 3476 10750 3488
rect 10965 3485 10977 3488
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3485 11207 3519
rect 11256 3516 11284 3556
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 12066 3584 12072 3596
rect 11388 3556 12072 3584
rect 11388 3544 11394 3556
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 12406 3584 12434 3624
rect 13357 3621 13369 3655
rect 13403 3652 13415 3655
rect 15102 3652 15108 3664
rect 13403 3624 15108 3652
rect 13403 3621 13415 3624
rect 13357 3615 13415 3621
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 15562 3612 15568 3664
rect 15620 3652 15626 3664
rect 15620 3624 15665 3652
rect 15620 3612 15626 3624
rect 16390 3612 16396 3664
rect 16448 3652 16454 3664
rect 22066 3652 22094 3692
rect 23658 3652 23664 3664
rect 16448 3624 22094 3652
rect 23619 3624 23664 3652
rect 16448 3612 16454 3624
rect 23658 3612 23664 3624
rect 23716 3612 23722 3664
rect 25777 3655 25835 3661
rect 25777 3621 25789 3655
rect 25823 3652 25835 3655
rect 26234 3652 26240 3664
rect 25823 3624 26240 3652
rect 25823 3621 25835 3624
rect 25777 3615 25835 3621
rect 26234 3612 26240 3624
rect 26292 3612 26298 3664
rect 27172 3652 27200 3692
rect 27246 3680 27252 3732
rect 27304 3720 27310 3732
rect 33318 3720 33324 3732
rect 27304 3692 33324 3720
rect 27304 3680 27310 3692
rect 33318 3680 33324 3692
rect 33376 3680 33382 3732
rect 33410 3680 33416 3732
rect 33468 3720 33474 3732
rect 35115 3723 35173 3729
rect 35115 3720 35127 3723
rect 33468 3692 35127 3720
rect 33468 3680 33474 3692
rect 35115 3689 35127 3692
rect 35161 3689 35173 3723
rect 35115 3683 35173 3689
rect 35526 3680 35532 3732
rect 35584 3720 35590 3732
rect 37458 3720 37464 3732
rect 35584 3692 37464 3720
rect 35584 3680 35590 3692
rect 37458 3680 37464 3692
rect 37516 3680 37522 3732
rect 40218 3720 40224 3732
rect 40179 3692 40224 3720
rect 40218 3680 40224 3692
rect 40276 3680 40282 3732
rect 41386 3692 55214 3720
rect 33042 3652 33048 3664
rect 27172 3624 33048 3652
rect 33042 3612 33048 3624
rect 33100 3612 33106 3664
rect 33520 3624 33732 3652
rect 12406 3556 15332 3584
rect 11793 3519 11851 3525
rect 11793 3516 11805 3519
rect 11256 3488 11805 3516
rect 11149 3479 11207 3485
rect 11793 3485 11805 3488
rect 11839 3485 11851 3519
rect 11793 3479 11851 3485
rect 6472 3420 7328 3448
rect 7392 3420 10456 3448
rect 6472 3380 6500 3420
rect 6638 3380 6644 3392
rect 4632 3352 6500 3380
rect 6599 3352 6644 3380
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7392 3380 7420 3420
rect 11164 3392 11192 3479
rect 11882 3476 11888 3528
rect 11940 3516 11946 3528
rect 11977 3519 12035 3525
rect 11977 3516 11989 3519
rect 11940 3488 11989 3516
rect 11940 3476 11946 3488
rect 11977 3485 11989 3488
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 13354 3476 13360 3528
rect 13412 3516 13418 3528
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13412 3488 13553 3516
rect 13412 3476 13418 3488
rect 13541 3485 13553 3488
rect 13587 3485 13599 3519
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 13541 3479 13599 3485
rect 14753 3488 14933 3516
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 12621 3451 12679 3457
rect 12621 3448 12633 3451
rect 11296 3420 12633 3448
rect 11296 3408 11302 3420
rect 12621 3417 12633 3420
rect 12667 3417 12679 3451
rect 12621 3411 12679 3417
rect 12894 3408 12900 3460
rect 12952 3448 12958 3460
rect 13998 3448 14004 3460
rect 12952 3420 14004 3448
rect 12952 3408 12958 3420
rect 13998 3408 14004 3420
rect 14056 3408 14062 3460
rect 9858 3380 9864 3392
rect 6880 3352 7420 3380
rect 9819 3352 9864 3380
rect 6880 3340 6886 3352
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 11146 3340 11152 3392
rect 11204 3340 11210 3392
rect 11333 3383 11391 3389
rect 11333 3349 11345 3383
rect 11379 3380 11391 3383
rect 11698 3380 11704 3392
rect 11379 3352 11704 3380
rect 11379 3349 11391 3352
rect 11333 3343 11391 3349
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 12158 3380 12164 3392
rect 12119 3352 12164 3380
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 13814 3340 13820 3392
rect 13872 3380 13878 3392
rect 14093 3383 14151 3389
rect 14093 3380 14105 3383
rect 13872 3352 14105 3380
rect 13872 3340 13878 3352
rect 14093 3349 14105 3352
rect 14139 3349 14151 3383
rect 14093 3343 14151 3349
rect 14550 3340 14556 3392
rect 14608 3380 14614 3392
rect 14753 3380 14781 3488
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 14921 3479 14979 3485
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 15304 3525 15332 3556
rect 16298 3544 16304 3596
rect 16356 3584 16362 3596
rect 16356 3556 17356 3584
rect 16356 3544 16362 3556
rect 15289 3519 15347 3525
rect 15068 3488 15113 3516
rect 15068 3476 15074 3488
rect 15289 3485 15301 3519
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 15427 3519 15485 3525
rect 15427 3485 15439 3519
rect 15473 3516 15485 3519
rect 15562 3516 15568 3528
rect 15473 3488 15568 3516
rect 15473 3485 15485 3488
rect 15427 3479 15485 3485
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 16022 3516 16028 3528
rect 15983 3488 16028 3516
rect 16022 3476 16028 3488
rect 16080 3476 16086 3528
rect 16206 3525 16212 3528
rect 16173 3519 16212 3525
rect 16173 3485 16185 3519
rect 16173 3479 16212 3485
rect 16206 3476 16212 3479
rect 16264 3476 16270 3528
rect 16482 3476 16488 3528
rect 16540 3525 16546 3528
rect 16540 3516 16548 3525
rect 17126 3516 17132 3528
rect 16540 3488 17132 3516
rect 16540 3479 16548 3488
rect 16540 3476 16546 3479
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 17328 3525 17356 3556
rect 17402 3544 17408 3596
rect 17460 3584 17466 3596
rect 17460 3556 21496 3584
rect 17460 3544 17466 3556
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3485 17371 3519
rect 17313 3479 17371 3485
rect 18690 3476 18696 3528
rect 18748 3516 18754 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 18748 3488 19441 3516
rect 18748 3476 18754 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 20254 3516 20260 3528
rect 20215 3488 20260 3516
rect 19429 3479 19487 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21361 3519 21419 3525
rect 21361 3516 21373 3519
rect 21140 3488 21373 3516
rect 21140 3476 21146 3488
rect 21361 3485 21373 3488
rect 21407 3485 21419 3519
rect 21468 3516 21496 3556
rect 21542 3544 21548 3596
rect 21600 3584 21606 3596
rect 22554 3584 22560 3596
rect 21600 3556 22560 3584
rect 21600 3544 21606 3556
rect 22554 3544 22560 3556
rect 22612 3544 22618 3596
rect 28166 3544 28172 3596
rect 28224 3584 28230 3596
rect 30558 3584 30564 3596
rect 28224 3556 30564 3584
rect 28224 3544 28230 3556
rect 30558 3544 30564 3556
rect 30616 3544 30622 3596
rect 31481 3587 31539 3593
rect 31481 3584 31493 3587
rect 30668 3556 31493 3584
rect 23474 3516 23480 3528
rect 21468 3488 23480 3516
rect 21361 3479 21419 3485
rect 23474 3476 23480 3488
rect 23532 3476 23538 3528
rect 23566 3476 23572 3528
rect 23624 3516 23630 3528
rect 23845 3519 23903 3525
rect 23845 3516 23857 3519
rect 23624 3488 23857 3516
rect 23624 3476 23630 3488
rect 23845 3485 23857 3488
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 24397 3519 24455 3525
rect 24397 3485 24409 3519
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 24664 3519 24722 3525
rect 24664 3485 24676 3519
rect 24710 3516 24722 3519
rect 24946 3516 24952 3528
rect 24710 3488 24952 3516
rect 24710 3485 24722 3488
rect 24664 3479 24722 3485
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 15194 3448 15200 3460
rect 14884 3420 15200 3448
rect 14884 3408 14890 3420
rect 15194 3408 15200 3420
rect 15252 3448 15258 3460
rect 16301 3451 16359 3457
rect 16301 3448 16313 3451
rect 15252 3420 16313 3448
rect 15252 3408 15258 3420
rect 16301 3417 16313 3420
rect 16347 3417 16359 3451
rect 16301 3411 16359 3417
rect 16393 3451 16451 3457
rect 16393 3417 16405 3451
rect 16439 3448 16451 3451
rect 16439 3420 17172 3448
rect 16439 3417 16451 3420
rect 16393 3411 16451 3417
rect 16022 3380 16028 3392
rect 14608 3352 16028 3380
rect 14608 3340 14614 3352
rect 16022 3340 16028 3352
rect 16080 3340 16086 3392
rect 16316 3380 16344 3411
rect 16482 3380 16488 3392
rect 16316 3352 16488 3380
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 16574 3340 16580 3392
rect 16632 3380 16638 3392
rect 17144 3389 17172 3420
rect 19150 3408 19156 3460
rect 19208 3448 19214 3460
rect 21818 3448 21824 3460
rect 19208 3420 21824 3448
rect 19208 3408 19214 3420
rect 21818 3408 21824 3420
rect 21876 3448 21882 3460
rect 23658 3448 23664 3460
rect 21876 3420 23664 3448
rect 21876 3408 21882 3420
rect 23658 3408 23664 3420
rect 23716 3448 23722 3460
rect 24412 3448 24440 3479
rect 24946 3476 24952 3488
rect 25004 3476 25010 3528
rect 26142 3516 26148 3528
rect 25056 3488 26148 3516
rect 25056 3448 25084 3488
rect 26142 3476 26148 3488
rect 26200 3516 26206 3528
rect 26237 3519 26295 3525
rect 26237 3516 26249 3519
rect 26200 3488 26249 3516
rect 26200 3476 26206 3488
rect 26237 3485 26249 3488
rect 26283 3485 26295 3519
rect 26237 3479 26295 3485
rect 26326 3476 26332 3528
rect 26384 3516 26390 3528
rect 26493 3519 26551 3525
rect 26493 3516 26505 3519
rect 26384 3488 26505 3516
rect 26384 3476 26390 3488
rect 26493 3485 26505 3488
rect 26539 3485 26551 3519
rect 26493 3479 26551 3485
rect 27430 3476 27436 3528
rect 27488 3516 27494 3528
rect 30668 3525 30696 3556
rect 31481 3553 31493 3556
rect 31527 3553 31539 3587
rect 31481 3547 31539 3553
rect 33134 3544 33140 3596
rect 33192 3584 33198 3596
rect 33520 3584 33548 3624
rect 33704 3593 33732 3624
rect 34054 3612 34060 3664
rect 34112 3652 34118 3664
rect 41386 3652 41414 3692
rect 34112 3624 41414 3652
rect 43533 3655 43591 3661
rect 34112 3612 34118 3624
rect 43533 3621 43545 3655
rect 43579 3652 43591 3655
rect 43990 3652 43996 3664
rect 43579 3624 43996 3652
rect 43579 3621 43591 3624
rect 43533 3615 43591 3621
rect 33192 3556 33548 3584
rect 33689 3587 33747 3593
rect 33192 3544 33198 3556
rect 33689 3553 33701 3587
rect 33735 3553 33747 3587
rect 33689 3547 33747 3553
rect 33781 3587 33839 3593
rect 33781 3553 33793 3587
rect 33827 3584 33839 3587
rect 35526 3584 35532 3596
rect 33827 3556 35532 3584
rect 33827 3553 33839 3556
rect 33781 3547 33839 3553
rect 35526 3544 35532 3556
rect 35584 3544 35590 3596
rect 36906 3544 36912 3596
rect 36964 3584 36970 3596
rect 37369 3587 37427 3593
rect 36964 3556 37320 3584
rect 36964 3544 36970 3556
rect 28261 3519 28319 3525
rect 28261 3516 28273 3519
rect 27488 3488 28273 3516
rect 27488 3476 27494 3488
rect 28261 3485 28273 3488
rect 28307 3485 28319 3519
rect 28261 3479 28319 3485
rect 30653 3519 30711 3525
rect 30653 3485 30665 3519
rect 30699 3485 30711 3519
rect 31110 3516 31116 3528
rect 31071 3488 31116 3516
rect 30653 3479 30711 3485
rect 31110 3476 31116 3488
rect 31168 3476 31174 3528
rect 31294 3516 31300 3528
rect 31255 3488 31300 3516
rect 31294 3476 31300 3488
rect 31352 3476 31358 3528
rect 33410 3516 33416 3528
rect 33371 3488 33416 3516
rect 33410 3476 33416 3488
rect 33468 3476 33474 3528
rect 33601 3519 33659 3525
rect 33601 3518 33613 3519
rect 33520 3490 33613 3518
rect 23716 3420 25084 3448
rect 23716 3408 23722 3420
rect 25406 3408 25412 3460
rect 25464 3448 25470 3460
rect 33318 3448 33324 3460
rect 25464 3420 33324 3448
rect 25464 3408 25470 3420
rect 33318 3408 33324 3420
rect 33376 3408 33382 3460
rect 16669 3383 16727 3389
rect 16669 3380 16681 3383
rect 16632 3352 16681 3380
rect 16632 3340 16638 3352
rect 16669 3349 16681 3352
rect 16715 3349 16727 3383
rect 16669 3343 16727 3349
rect 17129 3383 17187 3389
rect 17129 3349 17141 3383
rect 17175 3349 17187 3383
rect 17129 3343 17187 3349
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 19245 3383 19303 3389
rect 19245 3380 19257 3383
rect 17552 3352 19257 3380
rect 17552 3340 17558 3352
rect 19245 3349 19257 3352
rect 19291 3349 19303 3383
rect 19245 3343 19303 3349
rect 20162 3340 20168 3392
rect 20220 3380 20226 3392
rect 20441 3383 20499 3389
rect 20441 3380 20453 3383
rect 20220 3352 20453 3380
rect 20220 3340 20226 3352
rect 20441 3349 20453 3352
rect 20487 3349 20499 3383
rect 21174 3380 21180 3392
rect 21135 3352 21180 3380
rect 20441 3343 20499 3349
rect 21174 3340 21180 3352
rect 21232 3340 21238 3392
rect 22186 3340 22192 3392
rect 22244 3380 22250 3392
rect 22830 3380 22836 3392
rect 22244 3352 22836 3380
rect 22244 3340 22250 3352
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 27617 3383 27675 3389
rect 27617 3349 27629 3383
rect 27663 3380 27675 3383
rect 27982 3380 27988 3392
rect 27663 3352 27988 3380
rect 27663 3349 27675 3352
rect 27617 3343 27675 3349
rect 27982 3340 27988 3352
rect 28040 3340 28046 3392
rect 28074 3340 28080 3392
rect 28132 3380 28138 3392
rect 30466 3380 30472 3392
rect 28132 3352 28177 3380
rect 30427 3352 30472 3380
rect 28132 3340 28138 3352
rect 30466 3340 30472 3352
rect 30524 3340 30530 3392
rect 33520 3380 33548 3490
rect 33592 3488 33613 3490
rect 33601 3485 33613 3488
rect 33647 3485 33659 3519
rect 33965 3519 34023 3525
rect 33965 3512 33977 3519
rect 33601 3479 33659 3485
rect 33888 3485 33977 3512
rect 34011 3485 34023 3519
rect 33888 3484 34023 3485
rect 33686 3380 33692 3392
rect 33520 3352 33692 3380
rect 33686 3340 33692 3352
rect 33744 3340 33750 3392
rect 33778 3340 33784 3392
rect 33836 3380 33842 3392
rect 33888 3380 33916 3484
rect 33965 3479 34023 3484
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34848 3488 34897 3516
rect 34848 3476 34854 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 34885 3479 34943 3485
rect 35342 3476 35348 3528
rect 35400 3516 35406 3528
rect 36173 3519 36231 3525
rect 36173 3516 36185 3519
rect 35400 3488 36185 3516
rect 35400 3476 35406 3488
rect 36173 3485 36185 3488
rect 36219 3485 36231 3519
rect 36173 3479 36231 3485
rect 37093 3519 37151 3525
rect 37093 3485 37105 3519
rect 37139 3516 37151 3519
rect 37182 3516 37188 3528
rect 37139 3488 37188 3516
rect 37139 3485 37151 3488
rect 37093 3479 37151 3485
rect 37182 3476 37188 3488
rect 37240 3476 37246 3528
rect 37292 3525 37320 3556
rect 37369 3553 37381 3587
rect 37415 3584 37427 3587
rect 37550 3584 37556 3596
rect 37415 3556 37556 3584
rect 37415 3553 37427 3556
rect 37369 3547 37427 3553
rect 37550 3544 37556 3556
rect 37608 3584 37614 3596
rect 38838 3584 38844 3596
rect 37608 3556 38844 3584
rect 37608 3544 37614 3556
rect 38838 3544 38844 3556
rect 38896 3544 38902 3596
rect 39114 3544 39120 3596
rect 39172 3584 39178 3596
rect 39172 3556 40080 3584
rect 39172 3544 39178 3556
rect 37277 3519 37335 3525
rect 37277 3485 37289 3519
rect 37323 3485 37335 3519
rect 37458 3516 37464 3528
rect 37419 3488 37464 3516
rect 37277 3479 37335 3485
rect 37458 3476 37464 3488
rect 37516 3476 37522 3528
rect 37645 3519 37703 3525
rect 37645 3485 37657 3519
rect 37691 3516 37703 3519
rect 37734 3516 37740 3528
rect 37691 3488 37740 3516
rect 37691 3485 37703 3488
rect 37645 3479 37703 3485
rect 37734 3476 37740 3488
rect 37792 3476 37798 3528
rect 38286 3516 38292 3528
rect 38247 3488 38292 3516
rect 38286 3476 38292 3488
rect 38344 3476 38350 3528
rect 38378 3476 38384 3528
rect 38436 3516 38442 3528
rect 39853 3519 39911 3525
rect 39853 3516 39865 3519
rect 38436 3488 39865 3516
rect 38436 3476 38442 3488
rect 39853 3485 39865 3488
rect 39899 3516 39911 3519
rect 39942 3516 39948 3528
rect 39899 3488 39948 3516
rect 39899 3485 39911 3488
rect 39853 3479 39911 3485
rect 39942 3476 39948 3488
rect 40000 3476 40006 3528
rect 40052 3525 40080 3556
rect 40037 3519 40095 3525
rect 40037 3485 40049 3519
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 41414 3476 41420 3528
rect 41472 3516 41478 3528
rect 42150 3516 42156 3528
rect 41472 3488 41517 3516
rect 42111 3488 42156 3516
rect 41472 3476 41478 3488
rect 42150 3476 42156 3488
rect 42208 3476 42214 3528
rect 42242 3476 42248 3528
rect 42300 3516 42306 3528
rect 42409 3519 42467 3525
rect 42409 3516 42421 3519
rect 42300 3488 42421 3516
rect 42300 3476 42306 3488
rect 42409 3485 42421 3488
rect 42455 3485 42467 3519
rect 42409 3479 42467 3485
rect 42702 3476 42708 3528
rect 42760 3516 42766 3528
rect 43548 3516 43576 3615
rect 43990 3612 43996 3624
rect 44048 3612 44054 3664
rect 55186 3652 55214 3692
rect 57146 3652 57152 3664
rect 55186 3624 57152 3652
rect 57146 3612 57152 3624
rect 57204 3612 57210 3664
rect 45738 3544 45744 3596
rect 45796 3584 45802 3596
rect 46474 3584 46480 3596
rect 45796 3556 46480 3584
rect 45796 3544 45802 3556
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 42760 3488 43576 3516
rect 45557 3519 45615 3525
rect 42760 3476 42766 3488
rect 45557 3485 45569 3519
rect 45603 3516 45615 3519
rect 46014 3516 46020 3528
rect 45603 3488 46020 3516
rect 45603 3485 45615 3488
rect 45557 3479 45615 3485
rect 46014 3476 46020 3488
rect 46072 3476 46078 3528
rect 57701 3519 57759 3525
rect 46584 3488 55214 3516
rect 34330 3408 34336 3460
rect 34388 3448 34394 3460
rect 46584 3448 46612 3488
rect 46750 3457 46756 3460
rect 46744 3448 46756 3457
rect 34388 3420 46612 3448
rect 46711 3420 46756 3448
rect 34388 3408 34394 3420
rect 46744 3411 46756 3420
rect 46750 3408 46756 3411
rect 46808 3408 46814 3460
rect 55186 3448 55214 3488
rect 57701 3485 57713 3519
rect 57747 3516 57759 3519
rect 58158 3516 58164 3528
rect 57747 3488 58164 3516
rect 57747 3485 57759 3488
rect 57701 3479 57759 3485
rect 58158 3476 58164 3488
rect 58216 3476 58222 3528
rect 57977 3451 58035 3457
rect 57977 3448 57989 3451
rect 55186 3420 57989 3448
rect 57977 3417 57989 3420
rect 58023 3417 58035 3451
rect 57977 3411 58035 3417
rect 33836 3352 33916 3380
rect 33836 3340 33842 3352
rect 34054 3340 34060 3392
rect 34112 3380 34118 3392
rect 34149 3383 34207 3389
rect 34149 3380 34161 3383
rect 34112 3352 34161 3380
rect 34112 3340 34118 3352
rect 34149 3349 34161 3352
rect 34195 3349 34207 3383
rect 34149 3343 34207 3349
rect 35342 3340 35348 3392
rect 35400 3380 35406 3392
rect 36357 3383 36415 3389
rect 36357 3380 36369 3383
rect 35400 3352 36369 3380
rect 35400 3340 35406 3352
rect 36357 3349 36369 3352
rect 36403 3349 36415 3383
rect 37826 3380 37832 3392
rect 37787 3352 37832 3380
rect 36357 3343 36415 3349
rect 37826 3340 37832 3352
rect 37884 3340 37890 3392
rect 38194 3340 38200 3392
rect 38252 3380 38258 3392
rect 38473 3383 38531 3389
rect 38473 3380 38485 3383
rect 38252 3352 38485 3380
rect 38252 3340 38258 3352
rect 38473 3349 38485 3352
rect 38519 3349 38531 3383
rect 38473 3343 38531 3349
rect 39666 3340 39672 3392
rect 39724 3380 39730 3392
rect 41601 3383 41659 3389
rect 41601 3380 41613 3383
rect 39724 3352 41613 3380
rect 39724 3340 39730 3352
rect 41601 3349 41613 3352
rect 41647 3349 41659 3383
rect 41601 3343 41659 3349
rect 45462 3340 45468 3392
rect 45520 3380 45526 3392
rect 45741 3383 45799 3389
rect 45741 3380 45753 3383
rect 45520 3352 45753 3380
rect 45520 3340 45526 3352
rect 45741 3349 45753 3352
rect 45787 3349 45799 3383
rect 45741 3343 45799 3349
rect 46198 3340 46204 3392
rect 46256 3380 46262 3392
rect 47857 3383 47915 3389
rect 47857 3380 47869 3383
rect 46256 3352 47869 3380
rect 46256 3340 46262 3352
rect 47857 3349 47869 3352
rect 47903 3349 47915 3383
rect 47857 3343 47915 3349
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 3326 3176 3332 3188
rect 1627 3148 3332 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 3878 3176 3884 3188
rect 3839 3148 3884 3176
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4709 3179 4767 3185
rect 4709 3145 4721 3179
rect 4755 3145 4767 3179
rect 6362 3176 6368 3188
rect 6323 3148 6368 3176
rect 4709 3139 4767 3145
rect 3602 3068 3608 3120
rect 3660 3108 3666 3120
rect 4724 3108 4752 3139
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 21634 3176 21640 3188
rect 7300 3148 21640 3176
rect 3660 3080 4752 3108
rect 5184 3080 7236 3108
rect 3660 3068 3666 3080
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3040 2743 3043
rect 2731 3012 3648 3040
rect 2731 3009 2743 3012
rect 2685 3003 2743 3009
rect 3510 2972 3516 2984
rect 3471 2944 3516 2972
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 3620 2972 3648 3012
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 4249 3043 4307 3049
rect 3752 3012 3797 3040
rect 3752 3000 3758 3012
rect 4249 3009 4261 3043
rect 4295 3040 4307 3043
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 4295 3012 4537 3040
rect 4295 3009 4307 3012
rect 4249 3003 4307 3009
rect 4525 3009 4537 3012
rect 4571 3040 4583 3043
rect 4982 3040 4988 3052
rect 4571 3012 4988 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 5184 2972 5212 3080
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 7098 3040 7104 3052
rect 6595 3012 7104 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 3620 2944 5212 2972
rect 5276 2972 5304 3003
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 6638 2972 6644 2984
rect 5276 2944 6644 2972
rect 6638 2932 6644 2944
rect 6696 2972 6702 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6696 2944 6837 2972
rect 6696 2932 6702 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 7208 2972 7236 3080
rect 7300 3049 7328 3148
rect 21634 3136 21640 3148
rect 21692 3136 21698 3188
rect 33502 3176 33508 3188
rect 21836 3148 32352 3176
rect 33415 3148 33508 3176
rect 9858 3117 9864 3120
rect 9852 3108 9864 3117
rect 7392 3080 8432 3108
rect 9819 3080 9864 3108
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7392 2972 7420 3080
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 8297 3043 8355 3049
rect 8297 3040 8309 3043
rect 7524 3012 8309 3040
rect 7524 3000 7530 3012
rect 8297 3009 8309 3012
rect 8343 3009 8355 3043
rect 8404 3040 8432 3080
rect 9852 3071 9864 3080
rect 9858 3068 9864 3071
rect 9916 3068 9922 3120
rect 10870 3068 10876 3120
rect 10928 3108 10934 3120
rect 11238 3108 11244 3120
rect 10928 3080 11244 3108
rect 10928 3068 10934 3080
rect 11238 3068 11244 3080
rect 11296 3068 11302 3120
rect 12158 3068 12164 3120
rect 12216 3108 12222 3120
rect 14458 3108 14464 3120
rect 12216 3080 13492 3108
rect 14371 3080 14464 3108
rect 12216 3068 12222 3080
rect 11698 3040 11704 3052
rect 8404 3012 11560 3040
rect 11659 3012 11704 3040
rect 8297 3003 8355 3009
rect 7208 2944 7420 2972
rect 6825 2935 6883 2941
rect 7926 2932 7932 2984
rect 7984 2972 7990 2984
rect 8757 2975 8815 2981
rect 8757 2972 8769 2975
rect 7984 2944 8769 2972
rect 7984 2932 7990 2944
rect 8757 2941 8769 2944
rect 8803 2941 8815 2975
rect 8757 2935 8815 2941
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 8996 2944 9597 2972
rect 8996 2932 9002 2944
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 11532 2972 11560 3012
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 12802 3040 12808 3052
rect 12763 3012 12808 3040
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 13464 3049 13492 3080
rect 14458 3068 14464 3080
rect 14516 3108 14522 3120
rect 14516 3080 14780 3108
rect 14516 3068 14522 3080
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3009 13507 3043
rect 13906 3040 13912 3052
rect 13867 3012 13912 3040
rect 13449 3003 13507 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14476 2972 14504 3068
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 14752 3049 14780 3080
rect 14918 3068 14924 3120
rect 14976 3108 14982 3120
rect 14976 3080 15021 3108
rect 14976 3068 14982 3080
rect 16482 3068 16488 3120
rect 16540 3108 16546 3120
rect 16540 3080 16988 3108
rect 16540 3068 16546 3080
rect 14652 3043 14710 3049
rect 14652 3040 14664 3043
rect 14608 3012 14664 3040
rect 14608 3000 14614 3012
rect 14652 3009 14664 3012
rect 14698 3009 14710 3043
rect 14752 3043 14823 3049
rect 14752 3012 14777 3043
rect 14652 3003 14710 3009
rect 14765 3009 14777 3012
rect 14811 3009 14823 3043
rect 14765 3003 14823 3009
rect 15010 3000 15016 3052
rect 15068 3040 15074 3052
rect 15151 3043 15209 3049
rect 15068 3012 15113 3040
rect 15068 3000 15074 3012
rect 15151 3009 15163 3043
rect 15197 3009 15209 3043
rect 15151 3003 15209 3009
rect 11532 2944 14504 2972
rect 15166 2972 15194 3003
rect 15286 3000 15292 3052
rect 15344 3040 15350 3052
rect 15749 3043 15807 3049
rect 15749 3040 15761 3043
rect 15344 3012 15761 3040
rect 15344 3000 15350 3012
rect 15749 3009 15761 3012
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 16022 3000 16028 3052
rect 16080 3040 16086 3052
rect 16676 3043 16734 3049
rect 16676 3040 16688 3043
rect 16080 3012 16688 3040
rect 16080 3000 16086 3012
rect 16676 3009 16688 3012
rect 16722 3009 16734 3043
rect 16676 3003 16734 3009
rect 16762 3043 16820 3049
rect 16762 3009 16774 3043
rect 16808 3040 16820 3043
rect 16850 3040 16856 3052
rect 16808 3012 16856 3040
rect 16808 3009 16820 3012
rect 16762 3003 16820 3009
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 16960 3049 16988 3080
rect 18138 3068 18144 3120
rect 18196 3108 18202 3120
rect 18782 3108 18788 3120
rect 18196 3080 18788 3108
rect 18196 3068 18202 3080
rect 18782 3068 18788 3080
rect 18840 3068 18846 3120
rect 18960 3111 19018 3117
rect 18960 3077 18972 3111
rect 19006 3108 19018 3111
rect 19242 3108 19248 3120
rect 19006 3080 19248 3108
rect 19006 3077 19018 3080
rect 18960 3071 19018 3077
rect 19242 3068 19248 3080
rect 19300 3068 19306 3120
rect 21836 3108 21864 3148
rect 20548 3080 21864 3108
rect 22088 3111 22146 3117
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3009 17003 3043
rect 16945 3003 17003 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 15562 2972 15568 2984
rect 15166 2944 15568 2972
rect 9585 2935 9643 2941
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 17052 2972 17080 3003
rect 17126 3000 17132 3052
rect 17184 3049 17190 3052
rect 17184 3040 17192 3049
rect 17773 3043 17831 3049
rect 17184 3012 17229 3040
rect 17184 3003 17192 3012
rect 17773 3009 17785 3043
rect 17819 3040 17831 3043
rect 20548 3040 20576 3080
rect 22088 3077 22100 3111
rect 22134 3108 22146 3111
rect 22646 3108 22652 3120
rect 22134 3080 22652 3108
rect 22134 3077 22146 3080
rect 22088 3071 22146 3077
rect 22646 3068 22652 3080
rect 22704 3068 22710 3120
rect 23928 3111 23986 3117
rect 23928 3077 23940 3111
rect 23974 3108 23986 3111
rect 24394 3108 24400 3120
rect 23974 3080 24400 3108
rect 23974 3077 23986 3080
rect 23928 3071 23986 3077
rect 24394 3068 24400 3080
rect 24452 3068 24458 3120
rect 27614 3117 27620 3120
rect 27608 3108 27620 3117
rect 27575 3080 27620 3108
rect 27608 3071 27620 3080
rect 27614 3068 27620 3071
rect 27672 3068 27678 3120
rect 28258 3068 28264 3120
rect 28316 3068 28322 3120
rect 30466 3117 30472 3120
rect 30460 3108 30472 3117
rect 30427 3080 30472 3108
rect 30460 3071 30472 3080
rect 30466 3068 30472 3071
rect 30524 3068 30530 3120
rect 17819 3012 20576 3040
rect 20625 3043 20683 3049
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 20625 3009 20637 3043
rect 20671 3009 20683 3043
rect 23658 3040 23664 3052
rect 23619 3012 23664 3040
rect 20625 3003 20683 3009
rect 17184 3000 17190 3003
rect 17494 2972 17500 2984
rect 17052 2944 17500 2972
rect 17494 2932 17500 2944
rect 17552 2932 17558 2984
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 18693 2975 18751 2981
rect 18693 2972 18705 2975
rect 18196 2944 18705 2972
rect 18196 2932 18202 2944
rect 18693 2941 18705 2944
rect 18739 2941 18751 2975
rect 18693 2935 18751 2941
rect 20438 2932 20444 2984
rect 20496 2972 20502 2984
rect 20640 2972 20668 3003
rect 23658 3000 23664 3012
rect 23716 3000 23722 3052
rect 23768 3012 25728 3040
rect 21818 2972 21824 2984
rect 20496 2944 20668 2972
rect 21779 2944 21824 2972
rect 20496 2932 20502 2944
rect 21818 2932 21824 2944
rect 21876 2932 21882 2984
rect 22830 2932 22836 2984
rect 22888 2972 22894 2984
rect 23768 2972 23796 3012
rect 22888 2944 23796 2972
rect 22888 2932 22894 2944
rect 4062 2864 4068 2916
rect 4120 2904 4126 2916
rect 5445 2907 5503 2913
rect 5445 2904 5457 2907
rect 4120 2876 5457 2904
rect 4120 2864 4126 2876
rect 5445 2873 5457 2876
rect 5491 2873 5503 2907
rect 5445 2867 5503 2873
rect 6454 2864 6460 2916
rect 6512 2904 6518 2916
rect 7469 2907 7527 2913
rect 7469 2904 7481 2907
rect 6512 2876 7481 2904
rect 6512 2864 6518 2876
rect 7469 2873 7481 2876
rect 7515 2873 7527 2907
rect 7469 2867 7527 2873
rect 7650 2864 7656 2916
rect 7708 2904 7714 2916
rect 7708 2876 9628 2904
rect 7708 2864 7714 2876
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 2869 2839 2927 2845
rect 2869 2836 2881 2839
rect 2648 2808 2881 2836
rect 2648 2796 2654 2808
rect 2869 2805 2881 2808
rect 2915 2805 2927 2839
rect 2869 2799 2927 2805
rect 6733 2839 6791 2845
rect 6733 2805 6745 2839
rect 6779 2836 6791 2839
rect 7742 2836 7748 2848
rect 6779 2808 7748 2836
rect 6779 2805 6791 2808
rect 6733 2799 6791 2805
rect 7742 2796 7748 2808
rect 7800 2796 7806 2848
rect 8113 2839 8171 2845
rect 8113 2805 8125 2839
rect 8159 2836 8171 2839
rect 9490 2836 9496 2848
rect 8159 2808 9496 2836
rect 8159 2805 8171 2808
rect 8113 2799 8171 2805
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 9600 2836 9628 2876
rect 10594 2864 10600 2916
rect 10652 2904 10658 2916
rect 10965 2907 11023 2913
rect 10965 2904 10977 2907
rect 10652 2876 10977 2904
rect 10652 2864 10658 2876
rect 10965 2873 10977 2876
rect 11011 2873 11023 2907
rect 10965 2867 11023 2873
rect 12621 2907 12679 2913
rect 12621 2873 12633 2907
rect 12667 2904 12679 2907
rect 12894 2904 12900 2916
rect 12667 2876 12900 2904
rect 12667 2873 12679 2876
rect 12621 2867 12679 2873
rect 12894 2864 12900 2876
rect 12952 2864 12958 2916
rect 13265 2907 13323 2913
rect 13265 2873 13277 2907
rect 13311 2904 13323 2907
rect 14734 2904 14740 2916
rect 13311 2876 14740 2904
rect 13311 2873 13323 2876
rect 13265 2867 13323 2873
rect 14734 2864 14740 2876
rect 14792 2864 14798 2916
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 15933 2907 15991 2913
rect 15933 2904 15945 2907
rect 14884 2876 15945 2904
rect 14884 2864 14890 2876
rect 15933 2873 15945 2876
rect 15979 2873 15991 2907
rect 15933 2867 15991 2873
rect 17218 2864 17224 2916
rect 17276 2904 17282 2916
rect 17313 2907 17371 2913
rect 17313 2904 17325 2907
rect 17276 2876 17325 2904
rect 17276 2864 17282 2876
rect 17313 2873 17325 2876
rect 17359 2873 17371 2907
rect 25041 2907 25099 2913
rect 17313 2867 17371 2873
rect 19996 2876 20944 2904
rect 10686 2836 10692 2848
rect 9600 2808 10692 2836
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 12066 2836 12072 2848
rect 11563 2808 12072 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 14093 2839 14151 2845
rect 14093 2805 14105 2839
rect 14139 2836 14151 2839
rect 15194 2836 15200 2848
rect 14139 2808 15200 2836
rect 14139 2805 14151 2808
rect 14093 2799 14151 2805
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 15289 2839 15347 2845
rect 15289 2805 15301 2839
rect 15335 2836 15347 2839
rect 16942 2836 16948 2848
rect 15335 2808 16948 2836
rect 15335 2805 15347 2808
rect 15289 2799 15347 2805
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 17678 2796 17684 2848
rect 17736 2836 17742 2848
rect 17957 2839 18015 2845
rect 17957 2836 17969 2839
rect 17736 2808 17969 2836
rect 17736 2796 17742 2808
rect 17957 2805 17969 2808
rect 18003 2805 18015 2839
rect 17957 2799 18015 2805
rect 18046 2796 18052 2848
rect 18104 2836 18110 2848
rect 19996 2836 20024 2876
rect 18104 2808 20024 2836
rect 18104 2796 18110 2808
rect 20070 2796 20076 2848
rect 20128 2836 20134 2848
rect 20128 2808 20173 2836
rect 20128 2796 20134 2808
rect 20254 2796 20260 2848
rect 20312 2836 20318 2848
rect 20809 2839 20867 2845
rect 20809 2836 20821 2839
rect 20312 2808 20821 2836
rect 20312 2796 20318 2808
rect 20809 2805 20821 2808
rect 20855 2805 20867 2839
rect 20916 2836 20944 2876
rect 23124 2876 23428 2904
rect 23124 2836 23152 2876
rect 20916 2808 23152 2836
rect 20809 2799 20867 2805
rect 23198 2796 23204 2848
rect 23256 2836 23262 2848
rect 23400 2836 23428 2876
rect 25041 2873 25053 2907
rect 25087 2904 25099 2907
rect 25590 2904 25596 2916
rect 25087 2876 25596 2904
rect 25087 2873 25099 2876
rect 25041 2867 25099 2873
rect 25590 2864 25596 2876
rect 25648 2864 25654 2916
rect 24854 2836 24860 2848
rect 23256 2808 23301 2836
rect 23400 2808 24860 2836
rect 23256 2796 23262 2808
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 25700 2836 25728 3012
rect 25958 3000 25964 3052
rect 26016 3040 26022 3052
rect 26237 3043 26295 3049
rect 26237 3040 26249 3043
rect 26016 3012 26249 3040
rect 26016 3000 26022 3012
rect 26237 3009 26249 3012
rect 26283 3009 26295 3043
rect 28276 3040 28304 3068
rect 26237 3003 26295 3009
rect 27356 3012 28304 3040
rect 30193 3043 30251 3049
rect 26142 2932 26148 2984
rect 26200 2972 26206 2984
rect 27356 2981 27384 3012
rect 30193 3009 30205 3043
rect 30239 3040 30251 3043
rect 31846 3040 31852 3052
rect 30239 3012 31852 3040
rect 30239 3009 30251 3012
rect 30193 3003 30251 3009
rect 31846 3000 31852 3012
rect 31904 3040 31910 3052
rect 32122 3040 32128 3052
rect 31904 3012 32128 3040
rect 31904 3000 31910 3012
rect 32122 3000 32128 3012
rect 32180 3000 32186 3052
rect 32324 3040 32352 3148
rect 33502 3136 33508 3148
rect 33560 3176 33566 3188
rect 33778 3176 33784 3188
rect 33560 3148 33784 3176
rect 33560 3136 33566 3148
rect 33778 3136 33784 3148
rect 33836 3136 33842 3188
rect 34146 3136 34152 3188
rect 34204 3176 34210 3188
rect 34204 3148 34836 3176
rect 34204 3136 34210 3148
rect 32392 3111 32450 3117
rect 32392 3077 32404 3111
rect 32438 3108 32450 3111
rect 34054 3108 34060 3120
rect 32438 3080 34060 3108
rect 32438 3077 32450 3080
rect 32392 3071 32450 3077
rect 34054 3068 34060 3080
rect 34112 3068 34118 3120
rect 34698 3117 34704 3120
rect 34692 3108 34704 3117
rect 34659 3080 34704 3108
rect 34692 3071 34704 3080
rect 34698 3068 34704 3071
rect 34756 3068 34762 3120
rect 34808 3108 34836 3148
rect 35802 3136 35808 3188
rect 35860 3176 35866 3188
rect 37734 3176 37740 3188
rect 35860 3148 37740 3176
rect 35860 3136 35866 3148
rect 37734 3136 37740 3148
rect 37792 3176 37798 3188
rect 38749 3179 38807 3185
rect 38749 3176 38761 3179
rect 37792 3148 38761 3176
rect 37792 3136 37798 3148
rect 38749 3145 38761 3148
rect 38795 3145 38807 3179
rect 38749 3139 38807 3145
rect 38838 3136 38844 3188
rect 38896 3176 38902 3188
rect 41141 3179 41199 3185
rect 41141 3176 41153 3179
rect 38896 3148 41153 3176
rect 38896 3136 38902 3148
rect 41141 3145 41153 3148
rect 41187 3145 41199 3179
rect 41141 3139 41199 3145
rect 44082 3136 44088 3188
rect 44140 3176 44146 3188
rect 47765 3179 47823 3185
rect 47765 3176 47777 3179
rect 44140 3148 47777 3176
rect 44140 3136 44146 3148
rect 47765 3145 47777 3148
rect 47811 3145 47823 3179
rect 47765 3139 47823 3145
rect 54846 3136 54852 3188
rect 54904 3176 54910 3188
rect 54904 3148 57928 3176
rect 54904 3136 54910 3148
rect 37636 3111 37694 3117
rect 34808 3080 36308 3108
rect 32324 3012 33916 3040
rect 27341 2975 27399 2981
rect 27341 2972 27353 2975
rect 26200 2944 27353 2972
rect 26200 2932 26206 2944
rect 27341 2941 27353 2944
rect 27387 2941 27399 2975
rect 33888 2972 33916 3012
rect 34330 3000 34336 3052
rect 34388 3040 34394 3052
rect 34425 3043 34483 3049
rect 34425 3040 34437 3043
rect 34388 3012 34437 3040
rect 34388 3000 34394 3012
rect 34425 3009 34437 3012
rect 34471 3009 34483 3043
rect 35434 3040 35440 3052
rect 34425 3003 34483 3009
rect 34532 3012 35440 3040
rect 34532 2972 34560 3012
rect 35434 3000 35440 3012
rect 35492 3040 35498 3052
rect 35710 3040 35716 3052
rect 35492 3012 35716 3040
rect 35492 3000 35498 3012
rect 35710 3000 35716 3012
rect 35768 3000 35774 3052
rect 36280 3049 36308 3080
rect 37636 3077 37648 3111
rect 37682 3108 37694 3111
rect 37826 3108 37832 3120
rect 37682 3080 37832 3108
rect 37682 3077 37694 3080
rect 37636 3071 37694 3077
rect 37826 3068 37832 3080
rect 37884 3068 37890 3120
rect 39850 3068 39856 3120
rect 39908 3108 39914 3120
rect 40006 3111 40064 3117
rect 40006 3108 40018 3111
rect 39908 3080 40018 3108
rect 39908 3068 39914 3080
rect 40006 3077 40018 3080
rect 40052 3077 40064 3111
rect 40006 3071 40064 3077
rect 41414 3068 41420 3120
rect 41472 3108 41478 3120
rect 43806 3117 43812 3120
rect 43800 3108 43812 3117
rect 41472 3080 42932 3108
rect 43767 3080 43812 3108
rect 41472 3068 41478 3080
rect 36265 3043 36323 3049
rect 36265 3009 36277 3043
rect 36311 3009 36323 3043
rect 36265 3003 36323 3009
rect 37369 3043 37427 3049
rect 37369 3009 37381 3043
rect 37415 3040 37427 3043
rect 39761 3043 39819 3049
rect 39761 3040 39773 3043
rect 37415 3012 39773 3040
rect 37415 3009 37427 3012
rect 37369 3003 37427 3009
rect 39761 3009 39773 3012
rect 39807 3040 39819 3043
rect 40310 3040 40316 3052
rect 39807 3012 40316 3040
rect 39807 3009 39819 3012
rect 39761 3003 39819 3009
rect 40310 3000 40316 3012
rect 40368 3040 40374 3052
rect 42150 3040 42156 3052
rect 40368 3012 42156 3040
rect 40368 3000 40374 3012
rect 42150 3000 42156 3012
rect 42208 3000 42214 3052
rect 42702 3040 42708 3052
rect 42663 3012 42708 3040
rect 42702 3000 42708 3012
rect 42760 3000 42766 3052
rect 42904 3040 42932 3080
rect 43800 3071 43812 3080
rect 43806 3068 43812 3071
rect 43864 3068 43870 3120
rect 45370 3068 45376 3120
rect 45428 3108 45434 3120
rect 45802 3111 45860 3117
rect 45802 3108 45814 3111
rect 45428 3080 45814 3108
rect 45428 3068 45434 3080
rect 45802 3077 45814 3080
rect 45848 3077 45860 3111
rect 45802 3071 45860 3077
rect 45922 3068 45928 3120
rect 45980 3108 45986 3120
rect 45980 3080 47624 3108
rect 45980 3068 45986 3080
rect 46198 3040 46204 3052
rect 42904 3012 46204 3040
rect 46198 3000 46204 3012
rect 46256 3000 46262 3052
rect 47596 3049 47624 3080
rect 48406 3068 48412 3120
rect 48464 3108 48470 3120
rect 48464 3080 51580 3108
rect 48464 3068 48470 3080
rect 47581 3043 47639 3049
rect 47581 3009 47593 3043
rect 47627 3009 47639 3043
rect 47581 3003 47639 3009
rect 48317 3043 48375 3049
rect 48317 3009 48329 3043
rect 48363 3009 48375 3043
rect 48317 3003 48375 3009
rect 33888 2944 34560 2972
rect 27341 2935 27399 2941
rect 35526 2932 35532 2984
rect 35584 2972 35590 2984
rect 37274 2972 37280 2984
rect 35584 2944 37280 2972
rect 35584 2932 35590 2944
rect 37274 2932 37280 2944
rect 37332 2932 37338 2984
rect 42168 2972 42196 3000
rect 43533 2975 43591 2981
rect 43533 2972 43545 2975
rect 42168 2944 43545 2972
rect 43533 2941 43545 2944
rect 43579 2941 43591 2975
rect 43533 2935 43591 2941
rect 45557 2975 45615 2981
rect 45557 2941 45569 2975
rect 45603 2941 45615 2975
rect 48332 2972 48360 3003
rect 49602 3000 49608 3052
rect 49660 3040 49666 3052
rect 49973 3043 50031 3049
rect 49973 3040 49985 3043
rect 49660 3012 49985 3040
rect 49660 3000 49666 3012
rect 49973 3009 49985 3012
rect 50019 3009 50031 3043
rect 49973 3003 50031 3009
rect 50982 3000 50988 3052
rect 51040 3040 51046 3052
rect 51445 3043 51503 3049
rect 51445 3040 51457 3043
rect 51040 3012 51457 3040
rect 51040 3000 51046 3012
rect 51445 3009 51457 3012
rect 51491 3009 51503 3043
rect 51552 3040 51580 3080
rect 52454 3068 52460 3120
rect 52512 3108 52518 3120
rect 57146 3108 57152 3120
rect 52512 3080 55214 3108
rect 57107 3080 57152 3108
rect 52512 3068 52518 3080
rect 52917 3043 52975 3049
rect 52917 3040 52929 3043
rect 51552 3012 52929 3040
rect 51445 3003 51503 3009
rect 52917 3009 52929 3012
rect 52963 3009 52975 3043
rect 52917 3003 52975 3009
rect 54389 3043 54447 3049
rect 54389 3009 54401 3043
rect 54435 3009 54447 3043
rect 55186 3040 55214 3080
rect 57146 3068 57152 3080
rect 57204 3068 57210 3120
rect 57900 3049 57928 3148
rect 55861 3043 55919 3049
rect 55861 3040 55873 3043
rect 55186 3012 55873 3040
rect 54389 3003 54447 3009
rect 55861 3009 55873 3012
rect 55907 3009 55919 3043
rect 55861 3003 55919 3009
rect 56873 3043 56931 3049
rect 56873 3009 56885 3043
rect 56919 3009 56931 3043
rect 56873 3003 56931 3009
rect 57885 3043 57943 3049
rect 57885 3009 57897 3043
rect 57931 3009 57943 3043
rect 57885 3003 57943 3009
rect 45557 2935 45615 2941
rect 46952 2944 48360 2972
rect 26050 2904 26056 2916
rect 26011 2876 26056 2904
rect 26050 2864 26056 2876
rect 26108 2864 26114 2916
rect 28721 2907 28779 2913
rect 28721 2873 28733 2907
rect 28767 2904 28779 2907
rect 29546 2904 29552 2916
rect 28767 2876 29552 2904
rect 28767 2873 28779 2876
rect 28721 2867 28779 2873
rect 29546 2864 29552 2876
rect 29604 2864 29610 2916
rect 34330 2904 34336 2916
rect 31128 2876 32168 2904
rect 31128 2836 31156 2876
rect 31570 2836 31576 2848
rect 25700 2808 31156 2836
rect 31531 2808 31576 2836
rect 31570 2796 31576 2808
rect 31628 2796 31634 2848
rect 32140 2836 32168 2876
rect 33704 2876 34336 2904
rect 33704 2836 33732 2876
rect 34330 2864 34336 2876
rect 34388 2864 34394 2916
rect 36449 2907 36507 2913
rect 36449 2904 36461 2907
rect 35360 2876 36461 2904
rect 32140 2808 33732 2836
rect 33778 2796 33784 2848
rect 33836 2836 33842 2848
rect 35360 2836 35388 2876
rect 36449 2873 36461 2876
rect 36495 2873 36507 2907
rect 36449 2867 36507 2873
rect 33836 2808 35388 2836
rect 33836 2796 33842 2808
rect 35710 2796 35716 2848
rect 35768 2836 35774 2848
rect 35805 2839 35863 2845
rect 35805 2836 35817 2839
rect 35768 2808 35817 2836
rect 35768 2796 35774 2808
rect 35805 2805 35817 2808
rect 35851 2805 35863 2839
rect 35805 2799 35863 2805
rect 36722 2796 36728 2848
rect 36780 2836 36786 2848
rect 38654 2836 38660 2848
rect 36780 2808 38660 2836
rect 36780 2796 36786 2808
rect 38654 2796 38660 2808
rect 38712 2796 38718 2848
rect 42610 2796 42616 2848
rect 42668 2836 42674 2848
rect 42889 2839 42947 2845
rect 42889 2836 42901 2839
rect 42668 2808 42901 2836
rect 42668 2796 42674 2808
rect 42889 2805 42901 2808
rect 42935 2805 42947 2839
rect 43548 2836 43576 2935
rect 44910 2904 44916 2916
rect 44871 2876 44916 2904
rect 44910 2864 44916 2876
rect 44968 2864 44974 2916
rect 45572 2836 45600 2935
rect 45738 2836 45744 2848
rect 43548 2808 45744 2836
rect 42889 2799 42947 2805
rect 45738 2796 45744 2808
rect 45796 2796 45802 2848
rect 45830 2796 45836 2848
rect 45888 2836 45894 2848
rect 46952 2845 46980 2944
rect 51534 2932 51540 2984
rect 51592 2972 51598 2984
rect 54404 2972 54432 3003
rect 51592 2944 54432 2972
rect 56888 2972 56916 3003
rect 59630 2972 59636 2984
rect 56888 2944 59636 2972
rect 51592 2932 51598 2944
rect 59630 2932 59636 2944
rect 59688 2932 59694 2984
rect 47026 2864 47032 2916
rect 47084 2904 47090 2916
rect 48501 2907 48559 2913
rect 48501 2904 48513 2907
rect 47084 2876 48513 2904
rect 47084 2864 47090 2876
rect 48501 2873 48513 2876
rect 48547 2873 48559 2907
rect 48501 2867 48559 2873
rect 46937 2839 46995 2845
rect 46937 2836 46949 2839
rect 45888 2808 46949 2836
rect 45888 2796 45894 2808
rect 46937 2805 46949 2808
rect 46983 2805 46995 2839
rect 46937 2799 46995 2805
rect 49878 2796 49884 2848
rect 49936 2836 49942 2848
rect 50157 2839 50215 2845
rect 50157 2836 50169 2839
rect 49936 2808 50169 2836
rect 49936 2796 49942 2808
rect 50157 2805 50169 2808
rect 50203 2805 50215 2839
rect 50157 2799 50215 2805
rect 51350 2796 51356 2848
rect 51408 2836 51414 2848
rect 51629 2839 51687 2845
rect 51629 2836 51641 2839
rect 51408 2808 51641 2836
rect 51408 2796 51414 2808
rect 51629 2805 51641 2808
rect 51675 2805 51687 2839
rect 51629 2799 51687 2805
rect 52822 2796 52828 2848
rect 52880 2836 52886 2848
rect 53101 2839 53159 2845
rect 53101 2836 53113 2839
rect 52880 2808 53113 2836
rect 52880 2796 52886 2808
rect 53101 2805 53113 2808
rect 53147 2805 53159 2839
rect 53101 2799 53159 2805
rect 54294 2796 54300 2848
rect 54352 2836 54358 2848
rect 54573 2839 54631 2845
rect 54573 2836 54585 2839
rect 54352 2808 54585 2836
rect 54352 2796 54358 2808
rect 54573 2805 54585 2808
rect 54619 2805 54631 2839
rect 54573 2799 54631 2805
rect 55766 2796 55772 2848
rect 55824 2836 55830 2848
rect 56045 2839 56103 2845
rect 56045 2836 56057 2839
rect 55824 2808 56057 2836
rect 55824 2796 55830 2808
rect 56045 2805 56057 2808
rect 56091 2805 56103 2839
rect 56045 2799 56103 2805
rect 58069 2839 58127 2845
rect 58069 2805 58081 2839
rect 58115 2836 58127 2839
rect 58710 2836 58716 2848
rect 58115 2808 58716 2836
rect 58115 2805 58127 2808
rect 58069 2799 58127 2805
rect 58710 2796 58716 2808
rect 58768 2796 58774 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 2038 2592 2044 2644
rect 2096 2632 2102 2644
rect 2777 2635 2835 2641
rect 2777 2632 2789 2635
rect 2096 2604 2789 2632
rect 2096 2592 2102 2604
rect 2777 2601 2789 2604
rect 2823 2601 2835 2635
rect 2777 2595 2835 2601
rect 3050 2592 3056 2644
rect 3108 2632 3114 2644
rect 5442 2632 5448 2644
rect 3108 2604 5448 2632
rect 3108 2592 3114 2604
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 13262 2632 13268 2644
rect 7064 2604 13268 2632
rect 7064 2592 7070 2604
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 15289 2635 15347 2641
rect 15289 2601 15301 2635
rect 15335 2632 15347 2635
rect 15378 2632 15384 2644
rect 15335 2604 15384 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 18414 2592 18420 2644
rect 18472 2632 18478 2644
rect 21358 2632 21364 2644
rect 18472 2604 21364 2632
rect 18472 2592 18478 2604
rect 21358 2592 21364 2604
rect 21416 2592 21422 2644
rect 28810 2632 28816 2644
rect 28771 2604 28816 2632
rect 28810 2592 28816 2604
rect 28868 2592 28874 2644
rect 29362 2592 29368 2644
rect 29420 2632 29426 2644
rect 29822 2632 29828 2644
rect 29420 2604 29828 2632
rect 29420 2592 29426 2604
rect 29822 2592 29828 2604
rect 29880 2592 29886 2644
rect 30282 2632 30288 2644
rect 30243 2604 30288 2632
rect 30282 2592 30288 2604
rect 30340 2592 30346 2644
rect 32858 2592 32864 2644
rect 32916 2632 32922 2644
rect 38013 2635 38071 2641
rect 38013 2632 38025 2635
rect 32916 2604 38025 2632
rect 32916 2592 32922 2604
rect 38013 2601 38025 2604
rect 38059 2601 38071 2635
rect 38013 2595 38071 2601
rect 38654 2592 38660 2644
rect 38712 2632 38718 2644
rect 38749 2635 38807 2641
rect 38749 2632 38761 2635
rect 38712 2604 38761 2632
rect 38712 2592 38718 2604
rect 38749 2601 38761 2604
rect 38795 2601 38807 2635
rect 38749 2595 38807 2601
rect 5994 2524 6000 2576
rect 6052 2564 6058 2576
rect 7285 2567 7343 2573
rect 7285 2564 7297 2567
rect 6052 2536 7297 2564
rect 6052 2524 6058 2536
rect 7285 2533 7297 2536
rect 7331 2533 7343 2567
rect 7285 2527 7343 2533
rect 9398 2524 9404 2576
rect 9456 2564 9462 2576
rect 10597 2567 10655 2573
rect 10597 2564 10609 2567
rect 9456 2536 10609 2564
rect 9456 2524 9462 2536
rect 10597 2533 10609 2536
rect 10643 2533 10655 2567
rect 10597 2527 10655 2533
rect 12342 2524 12348 2576
rect 12400 2564 12406 2576
rect 13173 2567 13231 2573
rect 13173 2564 13185 2567
rect 12400 2536 13185 2564
rect 12400 2524 12406 2536
rect 13173 2533 13185 2536
rect 13219 2533 13231 2567
rect 16850 2564 16856 2576
rect 13173 2527 13231 2533
rect 13924 2536 16856 2564
rect 13722 2496 13728 2508
rect 6380 2468 13728 2496
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 6380 2437 6408 2468
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 1486 2360 1492 2372
rect 1447 2332 1492 2360
rect 1486 2320 1492 2332
rect 1544 2320 1550 2372
rect 4908 2360 4936 2391
rect 6546 2388 6552 2440
rect 6604 2428 6610 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6604 2400 7113 2428
rect 6604 2388 6610 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 8938 2428 8944 2440
rect 8899 2400 8944 2428
rect 7101 2391 7159 2397
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9490 2428 9496 2440
rect 9451 2400 9496 2428
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 10137 2431 10195 2437
rect 10137 2397 10149 2431
rect 10183 2428 10195 2431
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 10183 2400 10425 2428
rect 10183 2397 10195 2400
rect 10137 2391 10195 2397
rect 10413 2397 10425 2400
rect 10459 2428 10471 2431
rect 10502 2428 10508 2440
rect 10459 2400 10508 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 12066 2428 12072 2440
rect 12027 2400 12072 2428
rect 11517 2391 11575 2397
rect 7006 2360 7012 2372
rect 4908 2332 7012 2360
rect 7006 2320 7012 2332
rect 7064 2320 7070 2372
rect 7837 2363 7895 2369
rect 7837 2360 7849 2363
rect 7208 2332 7849 2360
rect 3050 2252 3056 2304
rect 3108 2292 3114 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3108 2264 3985 2292
rect 3108 2252 3114 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 5592 2264 6561 2292
rect 5592 2252 5598 2264
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 6549 2255 6607 2261
rect 6638 2252 6644 2304
rect 6696 2292 6702 2304
rect 7208 2292 7236 2332
rect 7837 2329 7849 2332
rect 7883 2329 7895 2363
rect 11532 2360 11560 2391
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 12986 2428 12992 2440
rect 12759 2400 12992 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 13924 2360 13952 2536
rect 16850 2524 16856 2536
rect 16908 2564 16914 2576
rect 18322 2564 18328 2576
rect 16908 2536 18328 2564
rect 16908 2524 16914 2536
rect 18322 2524 18328 2536
rect 18380 2564 18386 2576
rect 18380 2536 18736 2564
rect 18380 2524 18386 2536
rect 14550 2388 14556 2440
rect 14608 2428 14614 2440
rect 14645 2431 14703 2437
rect 14645 2428 14657 2431
rect 14608 2400 14657 2428
rect 14608 2388 14614 2400
rect 14645 2397 14657 2400
rect 14691 2397 14703 2431
rect 14645 2391 14703 2397
rect 14793 2431 14851 2437
rect 14793 2397 14805 2431
rect 14839 2397 14851 2431
rect 14918 2428 14924 2440
rect 14879 2400 14924 2428
rect 14793 2391 14851 2397
rect 14808 2360 14836 2391
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 15010 2388 15016 2440
rect 15068 2428 15074 2440
rect 15151 2431 15209 2437
rect 15068 2400 15113 2428
rect 15068 2388 15074 2400
rect 15151 2397 15163 2431
rect 15197 2428 15209 2431
rect 15562 2428 15568 2440
rect 15197 2400 15568 2428
rect 15197 2397 15209 2400
rect 15151 2391 15209 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15746 2428 15752 2440
rect 15707 2400 15752 2428
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16850 2428 16856 2440
rect 16811 2400 16856 2428
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17586 2428 17592 2440
rect 17547 2400 17592 2428
rect 17586 2388 17592 2400
rect 17644 2388 17650 2440
rect 18414 2388 18420 2440
rect 18472 2428 18478 2440
rect 18708 2428 18736 2536
rect 25038 2524 25044 2576
rect 25096 2564 25102 2576
rect 26053 2567 26111 2573
rect 26053 2564 26065 2567
rect 25096 2536 26065 2564
rect 25096 2524 25102 2536
rect 26053 2533 26065 2536
rect 26099 2533 26111 2567
rect 26053 2527 26111 2533
rect 29638 2524 29644 2576
rect 29696 2564 29702 2576
rect 29696 2536 35020 2564
rect 29696 2524 29702 2536
rect 18782 2456 18788 2508
rect 18840 2496 18846 2508
rect 19242 2496 19248 2508
rect 18840 2468 19248 2496
rect 18840 2456 18846 2468
rect 19242 2456 19248 2468
rect 19300 2456 19306 2508
rect 29454 2456 29460 2508
rect 29512 2496 29518 2508
rect 29512 2468 30972 2496
rect 29512 2456 29518 2468
rect 19518 2437 19524 2440
rect 18472 2400 18517 2428
rect 18708 2400 19380 2428
rect 18472 2388 18478 2400
rect 19242 2360 19248 2372
rect 11532 2332 13952 2360
rect 14016 2332 19248 2360
rect 7837 2323 7895 2329
rect 6696 2264 7236 2292
rect 6696 2252 6702 2264
rect 8478 2252 8484 2304
rect 8536 2292 8542 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8536 2264 9137 2292
rect 8536 2252 8542 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 9214 2252 9220 2304
rect 9272 2292 9278 2304
rect 9677 2295 9735 2301
rect 9677 2292 9689 2295
rect 9272 2264 9689 2292
rect 9272 2252 9278 2264
rect 9677 2261 9689 2264
rect 9723 2261 9735 2295
rect 9677 2255 9735 2261
rect 11330 2252 11336 2304
rect 11388 2292 11394 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11388 2264 11713 2292
rect 11388 2252 11394 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 12253 2295 12311 2301
rect 12253 2292 12265 2295
rect 11940 2264 12265 2292
rect 11940 2252 11946 2264
rect 12253 2261 12265 2264
rect 12299 2261 12311 2295
rect 12253 2255 12311 2261
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 14016 2292 14044 2332
rect 19242 2320 19248 2332
rect 19300 2320 19306 2372
rect 13780 2264 14044 2292
rect 13780 2252 13786 2264
rect 14274 2252 14280 2304
rect 14332 2292 14338 2304
rect 15933 2295 15991 2301
rect 15933 2292 15945 2295
rect 14332 2264 15945 2292
rect 14332 2252 14338 2264
rect 15933 2261 15945 2264
rect 15979 2261 15991 2295
rect 15933 2255 15991 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 17218 2252 17224 2304
rect 17276 2292 17282 2304
rect 17773 2295 17831 2301
rect 17773 2292 17785 2295
rect 17276 2264 17785 2292
rect 17276 2252 17282 2264
rect 17773 2261 17785 2264
rect 17819 2261 17831 2295
rect 17773 2255 17831 2261
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2292 18659 2295
rect 19150 2292 19156 2304
rect 18647 2264 19156 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 19150 2252 19156 2264
rect 19208 2252 19214 2304
rect 19352 2292 19380 2400
rect 19512 2391 19524 2437
rect 19576 2428 19582 2440
rect 21821 2431 21879 2437
rect 19576 2400 19612 2428
rect 19518 2388 19524 2391
rect 19576 2388 19582 2400
rect 21821 2397 21833 2431
rect 21867 2428 21879 2431
rect 22278 2428 22284 2440
rect 21867 2400 22284 2428
rect 21867 2397 21879 2400
rect 21821 2391 21879 2397
rect 22278 2388 22284 2400
rect 22336 2388 22342 2440
rect 22554 2428 22560 2440
rect 22515 2400 22560 2428
rect 22554 2388 22560 2400
rect 22612 2388 22618 2440
rect 23290 2428 23296 2440
rect 23251 2400 23296 2428
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2428 24455 2431
rect 24762 2428 24768 2440
rect 24443 2400 24768 2428
rect 24443 2397 24455 2400
rect 24397 2391 24455 2397
rect 24762 2388 24768 2400
rect 24820 2388 24826 2440
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 25133 2431 25191 2437
rect 25133 2428 25145 2431
rect 24912 2400 25145 2428
rect 24912 2388 24918 2400
rect 25133 2397 25145 2400
rect 25179 2397 25191 2431
rect 25133 2391 25191 2397
rect 25682 2388 25688 2440
rect 25740 2428 25746 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 25740 2400 25881 2428
rect 25740 2388 25746 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26234 2388 26240 2440
rect 26292 2428 26298 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26292 2400 26985 2428
rect 26292 2388 26298 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 28074 2428 28080 2440
rect 28035 2400 28080 2428
rect 26973 2391 27031 2397
rect 28074 2388 28080 2400
rect 28132 2388 28138 2440
rect 28902 2388 28908 2440
rect 28960 2428 28966 2440
rect 28997 2431 29055 2437
rect 28997 2428 29009 2431
rect 28960 2400 29009 2428
rect 28960 2388 28966 2400
rect 28997 2397 29009 2400
rect 29043 2397 29055 2431
rect 29546 2428 29552 2440
rect 29507 2400 29552 2428
rect 28997 2391 29055 2397
rect 29546 2388 29552 2400
rect 29604 2388 29610 2440
rect 29730 2388 29736 2440
rect 29788 2388 29794 2440
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 30944 2437 30972 2468
rect 31386 2456 31392 2508
rect 31444 2496 31450 2508
rect 32401 2499 32459 2505
rect 32401 2496 32413 2499
rect 31444 2468 32413 2496
rect 31444 2456 31450 2468
rect 32401 2465 32413 2468
rect 32447 2465 32459 2499
rect 32401 2459 32459 2465
rect 33318 2456 33324 2508
rect 33376 2496 33382 2508
rect 34992 2505 35020 2536
rect 35158 2524 35164 2576
rect 35216 2564 35222 2576
rect 43073 2567 43131 2573
rect 43073 2564 43085 2567
rect 35216 2536 43085 2564
rect 35216 2524 35222 2536
rect 43073 2533 43085 2536
rect 43119 2533 43131 2567
rect 43073 2527 43131 2533
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 33376 2468 34713 2496
rect 33376 2456 33382 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 34701 2459 34759 2465
rect 34977 2499 35035 2505
rect 34977 2465 34989 2499
rect 35023 2465 35035 2499
rect 34977 2459 35035 2465
rect 35066 2456 35072 2508
rect 35124 2496 35130 2508
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 35124 2468 40509 2496
rect 35124 2456 35130 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 40497 2459 40555 2465
rect 54386 2456 54392 2508
rect 54444 2496 54450 2508
rect 54444 2468 57928 2496
rect 54444 2456 54450 2468
rect 30469 2431 30527 2437
rect 30469 2428 30481 2431
rect 30432 2400 30481 2428
rect 30432 2388 30438 2400
rect 30469 2397 30481 2400
rect 30515 2397 30527 2431
rect 30469 2391 30527 2397
rect 30929 2431 30987 2437
rect 30929 2397 30941 2431
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 31846 2388 31852 2440
rect 31904 2428 31910 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31904 2400 32137 2428
rect 31904 2388 31910 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 33413 2431 33471 2437
rect 33413 2397 33425 2431
rect 33459 2428 33471 2431
rect 33594 2428 33600 2440
rect 33459 2400 33600 2428
rect 33459 2397 33471 2400
rect 33413 2391 33471 2397
rect 33594 2388 33600 2400
rect 33652 2388 33658 2440
rect 33888 2400 34100 2428
rect 19426 2320 19432 2372
rect 19484 2360 19490 2372
rect 29748 2360 29776 2388
rect 19484 2332 29776 2360
rect 19484 2320 19490 2332
rect 29822 2320 29828 2372
rect 29880 2360 29886 2372
rect 33888 2360 33916 2400
rect 29880 2332 33916 2360
rect 34072 2360 34100 2400
rect 34146 2388 34152 2440
rect 34204 2428 34210 2440
rect 37366 2428 37372 2440
rect 34204 2400 37372 2428
rect 34204 2388 34210 2400
rect 37366 2388 37372 2400
rect 37424 2388 37430 2440
rect 38565 2431 38623 2437
rect 38565 2397 38577 2431
rect 38611 2428 38623 2431
rect 42426 2428 42432 2440
rect 38611 2400 42432 2428
rect 38611 2397 38623 2400
rect 38565 2391 38623 2397
rect 42426 2388 42432 2400
rect 42484 2388 42490 2440
rect 48498 2388 48504 2440
rect 48556 2428 48562 2440
rect 48777 2431 48835 2437
rect 48777 2428 48789 2431
rect 48556 2400 48789 2428
rect 48556 2388 48562 2400
rect 48777 2397 48789 2400
rect 48823 2397 48835 2431
rect 48777 2391 48835 2397
rect 52362 2388 52368 2440
rect 52420 2428 52426 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52420 2400 52745 2428
rect 52420 2388 52426 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 53834 2388 53840 2440
rect 53892 2428 53898 2440
rect 53929 2431 53987 2437
rect 53929 2428 53941 2431
rect 53892 2400 53941 2428
rect 53892 2388 53898 2400
rect 53929 2397 53941 2400
rect 53975 2397 53987 2431
rect 53929 2391 53987 2397
rect 55214 2388 55220 2440
rect 55272 2428 55278 2440
rect 55309 2431 55367 2437
rect 55309 2428 55321 2431
rect 55272 2400 55321 2428
rect 55272 2388 55278 2400
rect 55309 2397 55321 2400
rect 55355 2397 55367 2431
rect 55309 2391 55367 2397
rect 56686 2388 56692 2440
rect 56744 2428 56750 2440
rect 57900 2437 57928 2468
rect 56781 2431 56839 2437
rect 56781 2428 56793 2431
rect 56744 2400 56793 2428
rect 56744 2388 56750 2400
rect 56781 2397 56793 2400
rect 56827 2397 56839 2431
rect 56781 2391 56839 2397
rect 57885 2431 57943 2437
rect 57885 2397 57897 2431
rect 57931 2397 57943 2431
rect 57885 2391 57943 2397
rect 34072 2332 34284 2360
rect 29880 2320 29886 2332
rect 20625 2295 20683 2301
rect 20625 2292 20637 2295
rect 19352 2264 20637 2292
rect 20625 2261 20637 2264
rect 20671 2261 20683 2295
rect 20625 2255 20683 2261
rect 21634 2252 21640 2304
rect 21692 2292 21698 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21692 2264 22017 2292
rect 21692 2252 21698 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 22094 2252 22100 2304
rect 22152 2292 22158 2304
rect 22741 2295 22799 2301
rect 22741 2292 22753 2295
rect 22152 2264 22753 2292
rect 22152 2252 22158 2264
rect 22741 2261 22753 2264
rect 22787 2261 22799 2295
rect 22741 2255 22799 2261
rect 22830 2252 22836 2304
rect 22888 2292 22894 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 22888 2264 23489 2292
rect 22888 2252 22894 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24084 2264 24593 2292
rect 24084 2252 24090 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 24670 2252 24676 2304
rect 24728 2292 24734 2304
rect 25317 2295 25375 2301
rect 25317 2292 25329 2295
rect 24728 2264 25329 2292
rect 24728 2252 24734 2264
rect 25317 2261 25329 2264
rect 25363 2261 25375 2295
rect 25317 2255 25375 2261
rect 26510 2252 26516 2304
rect 26568 2292 26574 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26568 2264 27169 2292
rect 26568 2252 26574 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 27982 2252 27988 2304
rect 28040 2292 28046 2304
rect 28261 2295 28319 2301
rect 28261 2292 28273 2295
rect 28040 2264 28273 2292
rect 28040 2252 28046 2264
rect 28261 2261 28273 2264
rect 28307 2261 28319 2295
rect 28261 2255 28319 2261
rect 29454 2252 29460 2304
rect 29512 2292 29518 2304
rect 29733 2295 29791 2301
rect 29733 2292 29745 2295
rect 29512 2264 29745 2292
rect 29512 2252 29518 2264
rect 29733 2261 29745 2264
rect 29779 2261 29791 2295
rect 29733 2255 29791 2261
rect 30834 2252 30840 2304
rect 30892 2292 30898 2304
rect 31113 2295 31171 2301
rect 31113 2292 31125 2295
rect 30892 2264 31125 2292
rect 30892 2252 30898 2264
rect 31113 2261 31125 2264
rect 31159 2261 31171 2295
rect 31113 2255 31171 2261
rect 32306 2252 32312 2304
rect 32364 2292 32370 2304
rect 33597 2295 33655 2301
rect 33597 2292 33609 2295
rect 32364 2264 33609 2292
rect 32364 2252 32370 2264
rect 33597 2261 33609 2264
rect 33643 2261 33655 2295
rect 34256 2292 34284 2332
rect 36262 2320 36268 2372
rect 36320 2360 36326 2372
rect 36449 2363 36507 2369
rect 36449 2360 36461 2363
rect 36320 2332 36461 2360
rect 36320 2320 36326 2332
rect 36449 2329 36461 2332
rect 36495 2329 36507 2363
rect 36449 2323 36507 2329
rect 37734 2320 37740 2372
rect 37792 2360 37798 2372
rect 37921 2363 37979 2369
rect 37921 2360 37933 2363
rect 37792 2332 37933 2360
rect 37792 2320 37798 2332
rect 37921 2329 37933 2332
rect 37967 2329 37979 2363
rect 37921 2323 37979 2329
rect 39206 2320 39212 2372
rect 39264 2360 39270 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39264 2332 40325 2360
rect 39264 2320 39270 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 41049 2363 41107 2369
rect 41049 2360 41061 2363
rect 40644 2332 41061 2360
rect 40644 2320 40650 2332
rect 41049 2329 41061 2332
rect 41095 2329 41107 2363
rect 41049 2323 41107 2329
rect 42058 2320 42064 2372
rect 42116 2360 42122 2372
rect 42889 2363 42947 2369
rect 42889 2360 42901 2363
rect 42116 2332 42901 2360
rect 42116 2320 42122 2332
rect 42889 2329 42901 2332
rect 42935 2329 42947 2363
rect 42889 2323 42947 2329
rect 43530 2320 43536 2372
rect 43588 2360 43594 2372
rect 43717 2363 43775 2369
rect 43717 2360 43729 2363
rect 43588 2332 43729 2360
rect 43588 2320 43594 2332
rect 43717 2329 43729 2332
rect 43763 2329 43775 2363
rect 43717 2323 43775 2329
rect 45002 2320 45008 2372
rect 45060 2360 45066 2372
rect 45465 2363 45523 2369
rect 45465 2360 45477 2363
rect 45060 2332 45477 2360
rect 45060 2320 45066 2332
rect 45465 2329 45477 2332
rect 45511 2329 45523 2363
rect 45465 2323 45523 2329
rect 46474 2320 46480 2372
rect 46532 2360 46538 2372
rect 46661 2363 46719 2369
rect 46661 2360 46673 2363
rect 46532 2332 46673 2360
rect 46532 2320 46538 2332
rect 46661 2329 46673 2332
rect 46707 2329 46719 2363
rect 46661 2323 46719 2329
rect 47946 2320 47952 2372
rect 48004 2360 48010 2372
rect 48133 2363 48191 2369
rect 48133 2360 48145 2363
rect 48004 2332 48145 2360
rect 48004 2320 48010 2332
rect 48133 2329 48145 2332
rect 48179 2329 48191 2363
rect 48133 2323 48191 2329
rect 49418 2320 49424 2372
rect 49476 2360 49482 2372
rect 50617 2363 50675 2369
rect 50617 2360 50629 2363
rect 49476 2332 50629 2360
rect 49476 2320 49482 2332
rect 50617 2329 50629 2332
rect 50663 2329 50675 2363
rect 50617 2323 50675 2329
rect 50890 2320 50896 2372
rect 50948 2360 50954 2372
rect 51537 2363 51595 2369
rect 51537 2360 51549 2363
rect 50948 2332 51549 2360
rect 50948 2320 50954 2332
rect 51537 2329 51549 2332
rect 51583 2329 51595 2363
rect 53006 2360 53012 2372
rect 52967 2332 53012 2360
rect 51537 2323 51595 2329
rect 53006 2320 53012 2332
rect 53064 2320 53070 2372
rect 54202 2360 54208 2372
rect 54163 2332 54208 2360
rect 54202 2320 54208 2332
rect 54260 2320 54266 2372
rect 55582 2360 55588 2372
rect 55543 2332 55588 2360
rect 55582 2320 55588 2332
rect 55640 2320 55646 2372
rect 57054 2360 57060 2372
rect 57015 2332 57060 2360
rect 57054 2320 57060 2332
rect 57112 2320 57118 2372
rect 36541 2295 36599 2301
rect 36541 2292 36553 2295
rect 34256 2264 36553 2292
rect 33597 2255 33655 2261
rect 36541 2261 36553 2264
rect 36587 2261 36599 2295
rect 36541 2255 36599 2261
rect 40494 2252 40500 2304
rect 40552 2292 40558 2304
rect 41141 2295 41199 2301
rect 41141 2292 41153 2295
rect 40552 2264 41153 2292
rect 40552 2252 40558 2264
rect 41141 2261 41153 2264
rect 41187 2261 41199 2295
rect 43806 2292 43812 2304
rect 43767 2264 43812 2292
rect 41141 2255 41199 2261
rect 43806 2252 43812 2264
rect 43864 2252 43870 2304
rect 45554 2252 45560 2304
rect 45612 2292 45618 2304
rect 46750 2292 46756 2304
rect 45612 2264 45657 2292
rect 46711 2264 46756 2292
rect 45612 2252 45618 2264
rect 46750 2252 46756 2264
rect 46808 2252 46814 2304
rect 48222 2292 48228 2304
rect 48183 2264 48228 2292
rect 48222 2252 48228 2264
rect 48280 2252 48286 2304
rect 48406 2252 48412 2304
rect 48464 2292 48470 2304
rect 48961 2295 49019 2301
rect 48961 2292 48973 2295
rect 48464 2264 48973 2292
rect 48464 2252 48470 2264
rect 48961 2261 48973 2264
rect 49007 2261 49019 2295
rect 50706 2292 50712 2304
rect 50667 2264 50712 2292
rect 48961 2255 49019 2261
rect 50706 2252 50712 2264
rect 50764 2252 50770 2304
rect 51626 2292 51632 2304
rect 51587 2264 51632 2292
rect 51626 2252 51632 2264
rect 51684 2252 51690 2304
rect 57238 2252 57244 2304
rect 57296 2292 57302 2304
rect 58069 2295 58127 2301
rect 58069 2292 58081 2295
rect 57296 2264 58081 2292
rect 57296 2252 57302 2264
rect 58069 2261 58081 2264
rect 58115 2261 58127 2295
rect 58069 2255 58127 2261
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 10502 2048 10508 2100
rect 10560 2088 10566 2100
rect 34146 2088 34152 2100
rect 10560 2060 34152 2088
rect 10560 2048 10566 2060
rect 34146 2048 34152 2060
rect 34204 2048 34210 2100
rect 34238 2048 34244 2100
rect 34296 2088 34302 2100
rect 34296 2060 41414 2088
rect 34296 2048 34302 2060
rect 12986 1980 12992 2032
rect 13044 2020 13050 2032
rect 35802 2020 35808 2032
rect 13044 1992 35808 2020
rect 13044 1980 13050 1992
rect 35802 1980 35808 1992
rect 35860 1980 35866 2032
rect 35894 1980 35900 2032
rect 35952 2020 35958 2032
rect 40678 2020 40684 2032
rect 35952 1992 40684 2020
rect 35952 1980 35958 1992
rect 40678 1980 40684 1992
rect 40736 1980 40742 2032
rect 41386 2020 41414 2060
rect 46750 2020 46756 2032
rect 41386 1992 46756 2020
rect 46750 1980 46756 1992
rect 46808 1980 46814 2032
rect 8938 1912 8944 1964
rect 8996 1952 9002 1964
rect 16114 1952 16120 1964
rect 8996 1924 16120 1952
rect 8996 1912 9002 1924
rect 16114 1912 16120 1924
rect 16172 1912 16178 1964
rect 16850 1912 16856 1964
rect 16908 1952 16914 1964
rect 22462 1952 22468 1964
rect 16908 1924 22468 1952
rect 16908 1912 16914 1924
rect 22462 1912 22468 1924
rect 22520 1912 22526 1964
rect 33962 1912 33968 1964
rect 34020 1952 34026 1964
rect 48222 1952 48228 1964
rect 34020 1924 48228 1952
rect 34020 1912 34026 1924
rect 48222 1912 48228 1924
rect 48280 1912 48286 1964
rect 9122 1844 9128 1896
rect 9180 1884 9186 1896
rect 55582 1884 55588 1896
rect 9180 1856 55588 1884
rect 9180 1844 9186 1856
rect 55582 1844 55588 1856
rect 55640 1844 55646 1896
rect 12526 1776 12532 1828
rect 12584 1816 12590 1828
rect 51626 1816 51632 1828
rect 12584 1788 51632 1816
rect 12584 1776 12590 1788
rect 51626 1776 51632 1788
rect 51684 1776 51690 1828
rect 12894 1708 12900 1760
rect 12952 1748 12958 1760
rect 50706 1748 50712 1760
rect 12952 1720 50712 1748
rect 12952 1708 12958 1720
rect 50706 1708 50712 1720
rect 50764 1708 50770 1760
rect 10594 1640 10600 1692
rect 10652 1680 10658 1692
rect 53006 1680 53012 1692
rect 10652 1652 53012 1680
rect 10652 1640 10658 1652
rect 53006 1640 53012 1652
rect 53064 1640 53070 1692
rect 8662 1572 8668 1624
rect 8720 1612 8726 1624
rect 54202 1612 54208 1624
rect 8720 1584 54208 1612
rect 8720 1572 8726 1584
rect 54202 1572 54208 1584
rect 54260 1572 54266 1624
rect 9306 1504 9312 1556
rect 9364 1544 9370 1556
rect 57054 1544 57060 1556
rect 9364 1516 57060 1544
rect 9364 1504 9370 1516
rect 57054 1504 57060 1516
rect 57112 1504 57118 1556
rect 15746 1436 15752 1488
rect 15804 1476 15810 1488
rect 23198 1476 23204 1488
rect 15804 1448 23204 1476
rect 15804 1436 15810 1448
rect 23198 1436 23204 1448
rect 23256 1436 23262 1488
rect 23290 1436 23296 1488
rect 23348 1476 23354 1488
rect 33502 1476 33508 1488
rect 23348 1448 33508 1476
rect 23348 1436 23354 1448
rect 33502 1436 33508 1448
rect 33560 1436 33566 1488
rect 33870 1436 33876 1488
rect 33928 1476 33934 1488
rect 33928 1448 40632 1476
rect 33928 1436 33934 1448
rect 5074 1368 5080 1420
rect 5132 1408 5138 1420
rect 6638 1408 6644 1420
rect 5132 1380 6644 1408
rect 5132 1368 5138 1380
rect 6638 1368 6644 1380
rect 6696 1368 6702 1420
rect 19702 1368 19708 1420
rect 19760 1408 19766 1420
rect 20254 1408 20260 1420
rect 19760 1380 20260 1408
rect 19760 1368 19766 1380
rect 20254 1368 20260 1380
rect 20312 1368 20318 1420
rect 33226 1368 33232 1420
rect 33284 1408 33290 1420
rect 40494 1408 40500 1420
rect 33284 1380 40500 1408
rect 33284 1368 33290 1380
rect 40494 1368 40500 1380
rect 40552 1368 40558 1420
rect 40604 1408 40632 1448
rect 40678 1436 40684 1488
rect 40736 1476 40742 1488
rect 43806 1476 43812 1488
rect 40736 1448 43812 1476
rect 40736 1436 40742 1448
rect 43806 1436 43812 1448
rect 43864 1436 43870 1488
rect 45554 1408 45560 1420
rect 40604 1380 45560 1408
rect 45554 1368 45560 1380
rect 45612 1368 45618 1420
<< via1 >>
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 2780 39584 2832 39636
rect 3056 39627 3108 39636
rect 3056 39593 3065 39627
rect 3065 39593 3099 39627
rect 3099 39593 3108 39627
rect 3056 39584 3108 39593
rect 3700 39584 3752 39636
rect 26240 39584 26292 39636
rect 41420 39627 41472 39636
rect 41420 39593 41429 39627
rect 41429 39593 41463 39627
rect 41463 39593 41472 39627
rect 41420 39584 41472 39593
rect 48688 39584 48740 39636
rect 56140 39584 56192 39636
rect 1492 39380 1544 39432
rect 8852 39448 8904 39500
rect 18696 39448 18748 39500
rect 3240 39380 3292 39432
rect 26976 39423 27028 39432
rect 26976 39389 26985 39423
rect 26985 39389 27019 39423
rect 27019 39389 27028 39423
rect 26976 39380 27028 39389
rect 33692 39380 33744 39432
rect 55404 39380 55456 39432
rect 1584 39287 1636 39296
rect 1584 39253 1593 39287
rect 1593 39253 1627 39287
rect 1627 39253 1636 39287
rect 1584 39244 1636 39253
rect 4436 39287 4488 39296
rect 4436 39253 4445 39287
rect 4445 39253 4479 39287
rect 4479 39253 4488 39287
rect 4436 39244 4488 39253
rect 34244 39244 34296 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4436 39040 4488 39092
rect 26976 39040 27028 39092
rect 35808 38972 35860 39024
rect 7196 38904 7248 38956
rect 35716 38904 35768 38956
rect 1584 38743 1636 38752
rect 1584 38709 1593 38743
rect 1593 38709 1627 38743
rect 1627 38709 1636 38743
rect 1584 38700 1636 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 2872 38496 2924 38548
rect 2412 38292 2464 38344
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 1768 37816 1820 37868
rect 1584 37655 1636 37664
rect 1584 37621 1593 37655
rect 1593 37621 1627 37655
rect 1627 37621 1636 37655
rect 1584 37612 1636 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 1676 36728 1728 36780
rect 1584 36635 1636 36644
rect 1584 36601 1593 36635
rect 1593 36601 1627 36635
rect 1627 36601 1636 36635
rect 1584 36592 1636 36601
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 12808 36116 12860 36168
rect 1584 36023 1636 36032
rect 1584 35989 1593 36023
rect 1593 35989 1627 36023
rect 1627 35989 1636 36023
rect 1584 35980 1636 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1860 35003 1912 35012
rect 1860 34969 1869 35003
rect 1869 34969 1903 35003
rect 1903 34969 1912 35003
rect 1860 34960 1912 34969
rect 1952 34935 2004 34944
rect 1952 34901 1961 34935
rect 1961 34901 1995 34935
rect 1995 34901 2004 34935
rect 1952 34892 2004 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 1584 34731 1636 34740
rect 1584 34697 1593 34731
rect 1593 34697 1627 34731
rect 1627 34697 1636 34731
rect 1584 34688 1636 34697
rect 5632 34688 5684 34740
rect 2320 34595 2372 34604
rect 2320 34561 2329 34595
rect 2329 34561 2363 34595
rect 2363 34561 2372 34595
rect 2320 34552 2372 34561
rect 5724 34484 5776 34536
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 13820 33940 13872 33992
rect 1584 33847 1636 33856
rect 1584 33813 1593 33847
rect 1593 33813 1627 33847
rect 1627 33813 1636 33847
rect 1584 33804 1636 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 1860 33507 1912 33516
rect 1860 33473 1869 33507
rect 1869 33473 1903 33507
rect 1903 33473 1912 33507
rect 1860 33464 1912 33473
rect 2872 33507 2924 33516
rect 2872 33473 2881 33507
rect 2881 33473 2915 33507
rect 2915 33473 2924 33507
rect 2872 33464 2924 33473
rect 2044 33371 2096 33380
rect 2044 33337 2053 33371
rect 2053 33337 2087 33371
rect 2087 33337 2096 33371
rect 2044 33328 2096 33337
rect 5540 33260 5592 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 10876 32852 10928 32904
rect 1584 32759 1636 32768
rect 1584 32725 1593 32759
rect 1593 32725 1627 32759
rect 1627 32725 1636 32759
rect 1584 32716 1636 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 1400 32419 1452 32428
rect 1400 32385 1409 32419
rect 1409 32385 1443 32419
rect 1443 32385 1452 32419
rect 1400 32376 1452 32385
rect 2228 32172 2280 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4988 31900 5040 31952
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 1860 31331 1912 31340
rect 1860 31297 1869 31331
rect 1869 31297 1903 31331
rect 1903 31297 1912 31331
rect 1860 31288 1912 31297
rect 1676 31152 1728 31204
rect 2320 31152 2372 31204
rect 25320 31084 25372 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1584 30923 1636 30932
rect 1584 30889 1593 30923
rect 1593 30889 1627 30923
rect 1627 30889 1636 30923
rect 1584 30880 1636 30889
rect 4896 30812 4948 30864
rect 1492 30676 1544 30728
rect 2964 30719 3016 30728
rect 2964 30685 2973 30719
rect 2973 30685 3007 30719
rect 3007 30685 3016 30719
rect 2964 30676 3016 30685
rect 4804 30719 4856 30728
rect 4804 30685 4813 30719
rect 4813 30685 4847 30719
rect 4847 30685 4856 30719
rect 4804 30676 4856 30685
rect 2872 30608 2924 30660
rect 2780 30583 2832 30592
rect 2780 30549 2789 30583
rect 2789 30549 2823 30583
rect 2823 30549 2832 30583
rect 2780 30540 2832 30549
rect 4712 30540 4764 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 2780 30379 2832 30388
rect 2780 30345 2789 30379
rect 2789 30345 2823 30379
rect 2823 30345 2832 30379
rect 2780 30336 2832 30345
rect 1400 30243 1452 30252
rect 1400 30209 1409 30243
rect 1409 30209 1443 30243
rect 1443 30209 1452 30243
rect 1400 30200 1452 30209
rect 2688 30243 2740 30252
rect 2688 30209 2697 30243
rect 2697 30209 2731 30243
rect 2731 30209 2740 30243
rect 2688 30200 2740 30209
rect 4712 30243 4764 30252
rect 4712 30209 4746 30243
rect 4746 30209 4764 30243
rect 4712 30200 4764 30209
rect 2964 30175 3016 30184
rect 2964 30141 2973 30175
rect 2973 30141 3007 30175
rect 3007 30141 3016 30175
rect 2964 30132 3016 30141
rect 4068 30132 4120 30184
rect 1584 30039 1636 30048
rect 1584 30005 1593 30039
rect 1593 30005 1627 30039
rect 1627 30005 1636 30039
rect 1584 29996 1636 30005
rect 3608 29996 3660 30048
rect 4620 29996 4672 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1400 29792 1452 29844
rect 6828 29835 6880 29844
rect 4712 29724 4764 29776
rect 6828 29801 6837 29835
rect 6837 29801 6871 29835
rect 6871 29801 6880 29835
rect 6828 29792 6880 29801
rect 7472 29792 7524 29844
rect 2964 29656 3016 29708
rect 4804 29699 4856 29708
rect 4804 29665 4813 29699
rect 4813 29665 4847 29699
rect 4847 29665 4856 29699
rect 4804 29656 4856 29665
rect 15108 29656 15160 29708
rect 4160 29588 4212 29640
rect 4620 29631 4672 29640
rect 4620 29597 4629 29631
rect 4629 29597 4663 29631
rect 4663 29597 4672 29631
rect 4620 29588 4672 29597
rect 4988 29588 5040 29640
rect 3424 29520 3476 29572
rect 7012 29631 7064 29640
rect 7012 29597 7021 29631
rect 7021 29597 7055 29631
rect 7055 29597 7064 29631
rect 7932 29631 7984 29640
rect 7012 29588 7064 29597
rect 7932 29597 7941 29631
rect 7941 29597 7975 29631
rect 7975 29597 7984 29631
rect 7932 29588 7984 29597
rect 7288 29520 7340 29572
rect 2688 29452 2740 29504
rect 6828 29452 6880 29504
rect 7380 29452 7432 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 3424 29291 3476 29300
rect 1860 29223 1912 29232
rect 1860 29189 1869 29223
rect 1869 29189 1903 29223
rect 1903 29189 1912 29223
rect 1860 29180 1912 29189
rect 3424 29257 3433 29291
rect 3433 29257 3467 29291
rect 3467 29257 3476 29291
rect 3424 29248 3476 29257
rect 7288 29248 7340 29300
rect 17408 29180 17460 29232
rect 3608 29155 3660 29164
rect 3608 29121 3617 29155
rect 3617 29121 3651 29155
rect 3651 29121 3660 29155
rect 3608 29112 3660 29121
rect 4160 29112 4212 29164
rect 7380 29112 7432 29164
rect 3976 29044 4028 29096
rect 5448 29044 5500 29096
rect 2596 28976 2648 29028
rect 2872 29019 2924 29028
rect 2872 28985 2881 29019
rect 2881 28985 2915 29019
rect 2915 28985 2924 29019
rect 2872 28976 2924 28985
rect 4620 28976 4672 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4068 28704 4120 28756
rect 7932 28704 7984 28756
rect 15108 28704 15160 28756
rect 4804 28568 4856 28620
rect 5540 28568 5592 28620
rect 7564 28611 7616 28620
rect 7564 28577 7573 28611
rect 7573 28577 7607 28611
rect 7607 28577 7616 28611
rect 7564 28568 7616 28577
rect 4896 28500 4948 28552
rect 7288 28543 7340 28552
rect 7288 28509 7297 28543
rect 7297 28509 7331 28543
rect 7331 28509 7340 28543
rect 7288 28500 7340 28509
rect 10876 28543 10928 28552
rect 1860 28475 1912 28484
rect 1860 28441 1869 28475
rect 1869 28441 1903 28475
rect 1903 28441 1912 28475
rect 1860 28432 1912 28441
rect 10876 28509 10885 28543
rect 10885 28509 10919 28543
rect 10919 28509 10928 28543
rect 10876 28500 10928 28509
rect 10968 28543 11020 28552
rect 10968 28509 10977 28543
rect 10977 28509 11011 28543
rect 11011 28509 11020 28543
rect 10968 28500 11020 28509
rect 12532 28500 12584 28552
rect 13452 28432 13504 28484
rect 14648 28432 14700 28484
rect 17040 28432 17092 28484
rect 2136 28407 2188 28416
rect 2136 28373 2145 28407
rect 2145 28373 2179 28407
rect 2179 28373 2188 28407
rect 2136 28364 2188 28373
rect 7012 28364 7064 28416
rect 10508 28407 10560 28416
rect 10508 28373 10517 28407
rect 10517 28373 10551 28407
rect 10551 28373 10560 28407
rect 10508 28364 10560 28373
rect 17408 28364 17460 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 2136 28160 2188 28212
rect 13820 28203 13872 28212
rect 2412 28067 2464 28076
rect 2412 28033 2421 28067
rect 2421 28033 2455 28067
rect 2455 28033 2464 28067
rect 2412 28024 2464 28033
rect 3056 28067 3108 28076
rect 3056 28033 3065 28067
rect 3065 28033 3099 28067
rect 3099 28033 3108 28067
rect 3056 28024 3108 28033
rect 3976 28024 4028 28076
rect 4620 28092 4672 28144
rect 10508 28092 10560 28144
rect 13820 28169 13829 28203
rect 13829 28169 13863 28203
rect 13863 28169 13872 28203
rect 13820 28160 13872 28169
rect 14648 28203 14700 28212
rect 14648 28169 14657 28203
rect 14657 28169 14691 28203
rect 14691 28169 14700 28203
rect 14648 28160 14700 28169
rect 15108 28160 15160 28212
rect 17040 28203 17092 28212
rect 17040 28169 17049 28203
rect 17049 28169 17083 28203
rect 17083 28169 17092 28203
rect 17040 28160 17092 28169
rect 17408 28203 17460 28212
rect 17408 28169 17417 28203
rect 17417 28169 17451 28203
rect 17451 28169 17460 28203
rect 17408 28160 17460 28169
rect 6828 28067 6880 28076
rect 6828 28033 6837 28067
rect 6837 28033 6871 28067
rect 6871 28033 6880 28067
rect 6828 28024 6880 28033
rect 9680 28024 9732 28076
rect 12532 28024 12584 28076
rect 12716 28067 12768 28076
rect 12716 28033 12750 28067
rect 12750 28033 12768 28067
rect 12716 28024 12768 28033
rect 16948 28024 17000 28076
rect 17224 28067 17276 28076
rect 17224 28033 17233 28067
rect 17233 28033 17267 28067
rect 17267 28033 17276 28067
rect 17224 28024 17276 28033
rect 7012 27888 7064 27940
rect 7656 27888 7708 27940
rect 1584 27863 1636 27872
rect 1584 27829 1593 27863
rect 1593 27829 1627 27863
rect 1627 27829 1636 27863
rect 1584 27820 1636 27829
rect 2136 27820 2188 27872
rect 2872 27863 2924 27872
rect 2872 27829 2881 27863
rect 2881 27829 2915 27863
rect 2915 27829 2924 27863
rect 2872 27820 2924 27829
rect 6644 27863 6696 27872
rect 6644 27829 6653 27863
rect 6653 27829 6687 27863
rect 6687 27829 6696 27863
rect 6644 27820 6696 27829
rect 16764 27956 16816 28008
rect 25504 27956 25556 28008
rect 10876 27888 10928 27940
rect 17960 27820 18012 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 6828 27616 6880 27668
rect 9680 27616 9732 27668
rect 12624 27616 12676 27668
rect 12716 27616 12768 27668
rect 5632 27480 5684 27532
rect 7564 27480 7616 27532
rect 8116 27480 8168 27532
rect 9680 27523 9732 27532
rect 9680 27489 9689 27523
rect 9689 27489 9723 27523
rect 9723 27489 9732 27523
rect 9680 27480 9732 27489
rect 1860 27455 1912 27464
rect 1860 27421 1869 27455
rect 1869 27421 1903 27455
rect 1903 27421 1912 27455
rect 1860 27412 1912 27421
rect 2136 27455 2188 27464
rect 2136 27421 2170 27455
rect 2170 27421 2188 27455
rect 2136 27412 2188 27421
rect 13912 27480 13964 27532
rect 2964 27344 3016 27396
rect 4804 27344 4856 27396
rect 5724 27344 5776 27396
rect 1492 27276 1544 27328
rect 3148 27276 3200 27328
rect 3792 27276 3844 27328
rect 7012 27276 7064 27328
rect 10508 27344 10560 27396
rect 10968 27344 11020 27396
rect 12900 27344 12952 27396
rect 13820 27344 13872 27396
rect 10876 27276 10928 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 2412 27072 2464 27124
rect 2872 27072 2924 27124
rect 3148 27072 3200 27124
rect 1492 27047 1544 27056
rect 1492 27013 1501 27047
rect 1501 27013 1535 27047
rect 1535 27013 1544 27047
rect 1492 27004 1544 27013
rect 3792 27004 3844 27056
rect 6644 27047 6696 27056
rect 6644 27013 6678 27047
rect 6678 27013 6696 27047
rect 6644 27004 6696 27013
rect 7012 27072 7064 27124
rect 10508 27115 10560 27124
rect 10508 27081 10517 27115
rect 10517 27081 10551 27115
rect 10551 27081 10560 27115
rect 10508 27072 10560 27081
rect 10876 27115 10928 27124
rect 10876 27081 10885 27115
rect 10885 27081 10919 27115
rect 10919 27081 10928 27115
rect 10876 27072 10928 27081
rect 16580 27004 16632 27056
rect 3700 26979 3752 26988
rect 3700 26945 3709 26979
rect 3709 26945 3743 26979
rect 3743 26945 3752 26979
rect 3700 26936 3752 26945
rect 10692 26979 10744 26988
rect 2964 26911 3016 26920
rect 2964 26877 2973 26911
rect 2973 26877 3007 26911
rect 3007 26877 3016 26911
rect 2964 26868 3016 26877
rect 3056 26868 3108 26920
rect 5448 26868 5500 26920
rect 5908 26868 5960 26920
rect 10692 26945 10701 26979
rect 10701 26945 10735 26979
rect 10735 26945 10744 26979
rect 10692 26936 10744 26945
rect 10968 26979 11020 26988
rect 10968 26945 10977 26979
rect 10977 26945 11011 26979
rect 11011 26945 11020 26979
rect 10968 26936 11020 26945
rect 15844 26936 15896 26988
rect 16948 26936 17000 26988
rect 17776 26936 17828 26988
rect 17316 26868 17368 26920
rect 3516 26775 3568 26784
rect 3516 26741 3525 26775
rect 3525 26741 3559 26775
rect 3559 26741 3568 26775
rect 3516 26732 3568 26741
rect 24492 26800 24544 26852
rect 10692 26732 10744 26784
rect 13728 26732 13780 26784
rect 16672 26775 16724 26784
rect 16672 26741 16681 26775
rect 16681 26741 16715 26775
rect 16715 26741 16724 26775
rect 16672 26732 16724 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3424 26528 3476 26580
rect 16580 26528 16632 26580
rect 18052 26528 18104 26580
rect 3700 26460 3752 26512
rect 3056 26324 3108 26376
rect 3240 26367 3292 26376
rect 3240 26333 3249 26367
rect 3249 26333 3283 26367
rect 3283 26333 3292 26367
rect 3240 26324 3292 26333
rect 1860 26256 1912 26308
rect 1584 26231 1636 26240
rect 1584 26197 1593 26231
rect 1593 26197 1627 26231
rect 1627 26197 1636 26231
rect 1584 26188 1636 26197
rect 2320 26231 2372 26240
rect 2320 26197 2329 26231
rect 2329 26197 2363 26231
rect 2363 26197 2372 26231
rect 2320 26188 2372 26197
rect 3700 26188 3752 26240
rect 15108 26256 15160 26308
rect 16672 26324 16724 26376
rect 13636 26188 13688 26240
rect 17408 26299 17460 26308
rect 17408 26265 17442 26299
rect 17442 26265 17460 26299
rect 17408 26256 17460 26265
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 3240 25984 3292 26036
rect 3516 26027 3568 26036
rect 3516 25993 3525 26027
rect 3525 25993 3559 26027
rect 3559 25993 3568 26027
rect 3516 25984 3568 25993
rect 1676 25916 1728 25968
rect 3424 25959 3476 25968
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 2320 25891 2372 25900
rect 2320 25857 2329 25891
rect 2329 25857 2363 25891
rect 2363 25857 2372 25891
rect 2320 25848 2372 25857
rect 3424 25925 3433 25959
rect 3433 25925 3467 25959
rect 3467 25925 3476 25959
rect 3424 25916 3476 25925
rect 9312 25984 9364 26036
rect 12808 25984 12860 26036
rect 17408 25984 17460 26036
rect 17960 25984 18012 26036
rect 4804 25916 4856 25968
rect 5540 25848 5592 25900
rect 5908 25848 5960 25900
rect 9496 25848 9548 25900
rect 9680 25916 9732 25968
rect 13636 25916 13688 25968
rect 10876 25848 10928 25900
rect 12624 25848 12676 25900
rect 13084 25848 13136 25900
rect 4804 25780 4856 25832
rect 13820 25848 13872 25900
rect 17776 25891 17828 25900
rect 17776 25857 17785 25891
rect 17785 25857 17819 25891
rect 17819 25857 17828 25891
rect 17776 25848 17828 25857
rect 19248 25780 19300 25832
rect 7288 25712 7340 25764
rect 2872 25644 2924 25696
rect 10968 25687 11020 25696
rect 10968 25653 10977 25687
rect 10977 25653 11011 25687
rect 11011 25653 11020 25687
rect 10968 25644 11020 25653
rect 15752 25687 15804 25696
rect 15752 25653 15761 25687
rect 15761 25653 15795 25687
rect 15795 25653 15804 25687
rect 15752 25644 15804 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1768 25440 1820 25492
rect 7196 25372 7248 25424
rect 9496 25440 9548 25492
rect 10876 25483 10928 25492
rect 10876 25449 10885 25483
rect 10885 25449 10919 25483
rect 10919 25449 10928 25483
rect 10876 25440 10928 25449
rect 13084 25483 13136 25492
rect 13084 25449 13093 25483
rect 13093 25449 13127 25483
rect 13127 25449 13136 25483
rect 13084 25440 13136 25449
rect 1860 25347 1912 25356
rect 1860 25313 1869 25347
rect 1869 25313 1903 25347
rect 1903 25313 1912 25347
rect 1860 25304 1912 25313
rect 5908 25347 5960 25356
rect 5908 25313 5917 25347
rect 5917 25313 5951 25347
rect 5951 25313 5960 25347
rect 5908 25304 5960 25313
rect 3884 25236 3936 25288
rect 8576 25236 8628 25288
rect 9312 25279 9364 25288
rect 2320 25168 2372 25220
rect 7748 25168 7800 25220
rect 3240 25143 3292 25152
rect 3240 25109 3249 25143
rect 3249 25109 3283 25143
rect 3283 25109 3292 25143
rect 3240 25100 3292 25109
rect 5540 25100 5592 25152
rect 8668 25168 8720 25220
rect 9312 25245 9321 25279
rect 9321 25245 9355 25279
rect 9355 25245 9364 25279
rect 9312 25236 9364 25245
rect 9680 25236 9732 25288
rect 8116 25143 8168 25152
rect 8116 25109 8125 25143
rect 8125 25109 8159 25143
rect 8159 25109 8168 25143
rect 8116 25100 8168 25109
rect 9036 25100 9088 25152
rect 10416 25279 10468 25288
rect 10416 25245 10423 25279
rect 10423 25245 10468 25279
rect 10416 25236 10468 25245
rect 10968 25372 11020 25424
rect 10692 25279 10744 25288
rect 10692 25245 10706 25279
rect 10706 25245 10740 25279
rect 10740 25245 10744 25279
rect 10692 25236 10744 25245
rect 12072 25236 12124 25288
rect 12532 25279 12584 25288
rect 12532 25245 12542 25279
rect 12542 25245 12576 25279
rect 12576 25245 12584 25279
rect 12808 25279 12860 25288
rect 12532 25236 12584 25245
rect 12808 25245 12817 25279
rect 12817 25245 12851 25279
rect 12851 25245 12860 25279
rect 12808 25236 12860 25245
rect 12900 25279 12952 25288
rect 12900 25245 12914 25279
rect 12914 25245 12948 25279
rect 12948 25245 12952 25279
rect 12900 25236 12952 25245
rect 13176 25236 13228 25288
rect 17132 25279 17184 25288
rect 17132 25245 17141 25279
rect 17141 25245 17175 25279
rect 17175 25245 17184 25279
rect 17132 25236 17184 25245
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 17776 25236 17828 25288
rect 17316 25211 17368 25220
rect 17316 25177 17325 25211
rect 17325 25177 17359 25211
rect 17359 25177 17368 25211
rect 17316 25168 17368 25177
rect 12900 25100 12952 25152
rect 16948 25143 17000 25152
rect 16948 25109 16957 25143
rect 16957 25109 16991 25143
rect 16991 25109 17000 25143
rect 16948 25100 17000 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 2320 24939 2372 24948
rect 2320 24905 2329 24939
rect 2329 24905 2363 24939
rect 2363 24905 2372 24939
rect 2320 24896 2372 24905
rect 7288 24896 7340 24948
rect 21640 24896 21692 24948
rect 5632 24828 5684 24880
rect 9036 24871 9088 24880
rect 9036 24837 9045 24871
rect 9045 24837 9079 24871
rect 9079 24837 9088 24871
rect 9036 24828 9088 24837
rect 1400 24803 1452 24812
rect 1400 24769 1409 24803
rect 1409 24769 1443 24803
rect 1443 24769 1452 24803
rect 1400 24760 1452 24769
rect 2228 24760 2280 24812
rect 3148 24803 3200 24812
rect 3148 24769 3157 24803
rect 3157 24769 3191 24803
rect 3191 24769 3200 24803
rect 3148 24760 3200 24769
rect 3792 24803 3844 24812
rect 3792 24769 3801 24803
rect 3801 24769 3835 24803
rect 3835 24769 3844 24803
rect 3792 24760 3844 24769
rect 4068 24803 4120 24812
rect 4068 24769 4077 24803
rect 4077 24769 4111 24803
rect 4111 24769 4120 24803
rect 4068 24760 4120 24769
rect 8576 24760 8628 24812
rect 8852 24803 8904 24812
rect 8852 24769 8862 24803
rect 8862 24769 8896 24803
rect 8896 24769 8904 24803
rect 8852 24760 8904 24769
rect 3424 24692 3476 24744
rect 7196 24692 7248 24744
rect 9680 24760 9732 24812
rect 10692 24760 10744 24812
rect 10784 24760 10836 24812
rect 13176 24828 13228 24880
rect 16948 24871 17000 24880
rect 16948 24837 16982 24871
rect 16982 24837 17000 24871
rect 16948 24828 17000 24837
rect 12532 24692 12584 24744
rect 2412 24624 2464 24676
rect 2688 24556 2740 24608
rect 3240 24556 3292 24608
rect 6184 24556 6236 24608
rect 7748 24556 7800 24608
rect 12072 24624 12124 24676
rect 12716 24803 12768 24812
rect 12716 24769 12726 24803
rect 12726 24769 12760 24803
rect 12760 24769 12768 24803
rect 12900 24803 12952 24812
rect 12716 24760 12768 24769
rect 12900 24769 12909 24803
rect 12909 24769 12943 24803
rect 12943 24769 12952 24803
rect 12900 24760 12952 24769
rect 15752 24692 15804 24744
rect 13820 24624 13872 24676
rect 15200 24624 15252 24676
rect 17316 24556 17368 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2228 24395 2280 24404
rect 2228 24361 2237 24395
rect 2237 24361 2271 24395
rect 2271 24361 2280 24395
rect 2228 24352 2280 24361
rect 4068 24352 4120 24404
rect 2688 24259 2740 24268
rect 2688 24225 2697 24259
rect 2697 24225 2731 24259
rect 2731 24225 2740 24259
rect 2688 24216 2740 24225
rect 3056 24216 3108 24268
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 3240 24148 3292 24200
rect 5632 24148 5684 24200
rect 24584 24352 24636 24404
rect 12900 24216 12952 24268
rect 12532 24191 12584 24200
rect 12532 24157 12541 24191
rect 12541 24157 12575 24191
rect 12575 24157 12584 24191
rect 12532 24148 12584 24157
rect 15200 24148 15252 24200
rect 4160 24080 4212 24132
rect 13820 24080 13872 24132
rect 17408 24148 17460 24200
rect 15752 24123 15804 24132
rect 15752 24089 15786 24123
rect 15786 24089 15804 24123
rect 15752 24080 15804 24089
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 3884 24012 3936 24064
rect 5448 24012 5500 24064
rect 11888 24012 11940 24064
rect 16028 24012 16080 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 4068 23808 4120 23860
rect 8944 23808 8996 23860
rect 4160 23740 4212 23792
rect 10784 23783 10836 23792
rect 10784 23749 10793 23783
rect 10793 23749 10827 23783
rect 10827 23749 10836 23783
rect 10784 23740 10836 23749
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 5540 23672 5592 23724
rect 6460 23672 6512 23724
rect 9312 23715 9364 23724
rect 9312 23681 9321 23715
rect 9321 23681 9355 23715
rect 9355 23681 9364 23715
rect 9312 23672 9364 23681
rect 9404 23715 9456 23724
rect 9404 23681 9414 23715
rect 9414 23681 9448 23715
rect 9448 23681 9456 23715
rect 9588 23715 9640 23724
rect 9404 23672 9456 23681
rect 9588 23681 9597 23715
rect 9597 23681 9631 23715
rect 9631 23681 9640 23715
rect 9588 23672 9640 23681
rect 3516 23647 3568 23656
rect 3516 23613 3525 23647
rect 3525 23613 3559 23647
rect 3559 23613 3568 23647
rect 3516 23604 3568 23613
rect 3148 23536 3200 23588
rect 7104 23604 7156 23656
rect 8944 23604 8996 23656
rect 10692 23672 10744 23724
rect 12716 23808 12768 23860
rect 15752 23808 15804 23860
rect 16120 23808 16172 23860
rect 15108 23740 15160 23792
rect 16028 23783 16080 23792
rect 16028 23749 16037 23783
rect 16037 23749 16071 23783
rect 16071 23749 16080 23783
rect 16028 23740 16080 23749
rect 11796 23715 11848 23724
rect 11796 23681 11830 23715
rect 11830 23681 11848 23715
rect 11796 23672 11848 23681
rect 17408 23604 17460 23656
rect 10968 23579 11020 23588
rect 10968 23545 10977 23579
rect 10977 23545 11011 23579
rect 11011 23545 11020 23579
rect 10968 23536 11020 23545
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 3608 23468 3660 23520
rect 11704 23468 11756 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 3516 23264 3568 23316
rect 2504 23196 2556 23248
rect 9036 23264 9088 23316
rect 11796 23264 11848 23316
rect 8576 23128 8628 23180
rect 9312 23128 9364 23180
rect 1400 23060 1452 23112
rect 2228 23103 2280 23112
rect 2228 23069 2237 23103
rect 2237 23069 2271 23103
rect 2271 23069 2280 23103
rect 2228 23060 2280 23069
rect 7104 23060 7156 23112
rect 10784 23060 10836 23112
rect 10968 23128 11020 23180
rect 11244 23103 11296 23112
rect 11244 23069 11253 23103
rect 11253 23069 11287 23103
rect 11287 23069 11296 23103
rect 11244 23060 11296 23069
rect 11336 23103 11388 23112
rect 11336 23069 11346 23103
rect 11346 23069 11380 23103
rect 11380 23069 11388 23103
rect 11612 23103 11664 23112
rect 11336 23060 11388 23069
rect 11612 23069 11618 23103
rect 11618 23069 11652 23103
rect 11652 23069 11664 23103
rect 11612 23060 11664 23069
rect 12716 23128 12768 23180
rect 15200 23264 15252 23316
rect 15752 23128 15804 23180
rect 11888 23060 11940 23112
rect 17316 23103 17368 23112
rect 9312 22992 9364 23044
rect 9588 22992 9640 23044
rect 12532 22992 12584 23044
rect 13268 22992 13320 23044
rect 2964 22924 3016 22976
rect 5632 22924 5684 22976
rect 9220 22924 9272 22976
rect 11428 22924 11480 22976
rect 11796 22924 11848 22976
rect 13820 22924 13872 22976
rect 17316 23069 17325 23103
rect 17325 23069 17359 23103
rect 17359 23069 17368 23103
rect 17316 23060 17368 23069
rect 19984 23103 20036 23112
rect 14188 22992 14240 23044
rect 17500 22992 17552 23044
rect 19984 23069 19993 23103
rect 19993 23069 20027 23103
rect 20027 23069 20036 23103
rect 19984 23060 20036 23069
rect 22468 23128 22520 23180
rect 20812 22992 20864 23044
rect 14464 22924 14516 22976
rect 15936 22924 15988 22976
rect 20352 22924 20404 22976
rect 27620 23103 27672 23112
rect 27620 23069 27629 23103
rect 27629 23069 27663 23103
rect 27663 23069 27672 23103
rect 27620 23060 27672 23069
rect 29736 23060 29788 23112
rect 33508 23103 33560 23112
rect 33508 23069 33517 23103
rect 33517 23069 33551 23103
rect 33551 23069 33560 23103
rect 33508 23060 33560 23069
rect 24676 23035 24728 23044
rect 24676 23001 24710 23035
rect 24710 23001 24728 23035
rect 24676 22992 24728 23001
rect 27988 22992 28040 23044
rect 25044 22924 25096 22976
rect 29552 22924 29604 22976
rect 33048 22967 33100 22976
rect 33048 22933 33057 22967
rect 33057 22933 33091 22967
rect 33091 22933 33100 22967
rect 33048 22924 33100 22933
rect 33416 22967 33468 22976
rect 33416 22933 33425 22967
rect 33425 22933 33459 22967
rect 33459 22933 33468 22967
rect 33416 22924 33468 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 1584 22720 1636 22772
rect 4896 22720 4948 22772
rect 9312 22763 9364 22772
rect 9312 22729 9321 22763
rect 9321 22729 9355 22763
rect 9355 22729 9364 22763
rect 9312 22720 9364 22729
rect 12440 22720 12492 22772
rect 12716 22720 12768 22772
rect 14188 22720 14240 22772
rect 14464 22763 14516 22772
rect 14464 22729 14473 22763
rect 14473 22729 14507 22763
rect 14507 22729 14516 22763
rect 14464 22720 14516 22729
rect 17224 22720 17276 22772
rect 20812 22763 20864 22772
rect 20812 22729 20821 22763
rect 20821 22729 20855 22763
rect 20855 22729 20864 22763
rect 20812 22720 20864 22729
rect 24676 22763 24728 22772
rect 24676 22729 24685 22763
rect 24685 22729 24719 22763
rect 24719 22729 24728 22763
rect 24676 22720 24728 22729
rect 25044 22763 25096 22772
rect 25044 22729 25053 22763
rect 25053 22729 25087 22763
rect 25087 22729 25096 22763
rect 25044 22720 25096 22729
rect 27988 22763 28040 22772
rect 27988 22729 27997 22763
rect 27997 22729 28031 22763
rect 28031 22729 28040 22763
rect 27988 22720 28040 22729
rect 28172 22720 28224 22772
rect 33416 22720 33468 22772
rect 2780 22584 2832 22636
rect 2872 22584 2924 22636
rect 3792 22627 3844 22636
rect 3792 22593 3801 22627
rect 3801 22593 3835 22627
rect 3835 22593 3844 22627
rect 3792 22584 3844 22593
rect 3884 22584 3936 22636
rect 8576 22584 8628 22636
rect 8852 22627 8904 22636
rect 8852 22593 8859 22627
rect 8859 22593 8904 22627
rect 8852 22584 8904 22593
rect 3148 22559 3200 22568
rect 3148 22525 3157 22559
rect 3157 22525 3191 22559
rect 3191 22525 3200 22559
rect 9036 22627 9088 22636
rect 9036 22593 9045 22627
rect 9045 22593 9079 22627
rect 9079 22593 9088 22627
rect 9036 22584 9088 22593
rect 9220 22584 9272 22636
rect 3148 22516 3200 22525
rect 9588 22516 9640 22568
rect 13820 22652 13872 22704
rect 13636 22627 13688 22636
rect 13636 22593 13645 22627
rect 13645 22593 13679 22627
rect 13679 22593 13688 22627
rect 13636 22584 13688 22593
rect 16120 22584 16172 22636
rect 17592 22584 17644 22636
rect 17684 22584 17736 22636
rect 20352 22652 20404 22704
rect 21272 22627 21324 22636
rect 16028 22516 16080 22568
rect 17776 22559 17828 22568
rect 17776 22525 17785 22559
rect 17785 22525 17819 22559
rect 17819 22525 17828 22559
rect 17776 22516 17828 22525
rect 17960 22559 18012 22568
rect 17960 22525 17969 22559
rect 17969 22525 18003 22559
rect 18003 22525 18012 22559
rect 21272 22593 21281 22627
rect 21281 22593 21315 22627
rect 21315 22593 21324 22627
rect 21272 22584 21324 22593
rect 25688 22652 25740 22704
rect 25044 22584 25096 22636
rect 33048 22652 33100 22704
rect 29644 22584 29696 22636
rect 30840 22584 30892 22636
rect 17960 22516 18012 22525
rect 25780 22516 25832 22568
rect 28264 22448 28316 22500
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 3976 22380 4028 22432
rect 17224 22380 17276 22432
rect 17500 22380 17552 22432
rect 18236 22380 18288 22432
rect 27620 22380 27672 22432
rect 32036 22380 32088 22432
rect 33692 22380 33744 22432
rect 34428 22423 34480 22432
rect 34428 22389 34437 22423
rect 34437 22389 34471 22423
rect 34471 22389 34480 22423
rect 34428 22380 34480 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3884 22176 3936 22228
rect 2780 22108 2832 22160
rect 10876 22108 10928 22160
rect 16304 22108 16356 22160
rect 17316 22176 17368 22228
rect 17776 22219 17828 22228
rect 17776 22185 17785 22219
rect 17785 22185 17819 22219
rect 17819 22185 17828 22219
rect 17776 22176 17828 22185
rect 25504 22219 25556 22228
rect 15660 22040 15712 22092
rect 15844 22040 15896 22092
rect 15936 22083 15988 22092
rect 15936 22049 15945 22083
rect 15945 22049 15979 22083
rect 15979 22049 15988 22083
rect 15936 22040 15988 22049
rect 16580 22040 16632 22092
rect 17224 22083 17276 22092
rect 17224 22049 17233 22083
rect 17233 22049 17267 22083
rect 17267 22049 17276 22083
rect 17224 22040 17276 22049
rect 19984 22108 20036 22160
rect 25504 22185 25513 22219
rect 25513 22185 25547 22219
rect 25547 22185 25556 22219
rect 25504 22176 25556 22185
rect 25688 22219 25740 22228
rect 25688 22185 25697 22219
rect 25697 22185 25731 22219
rect 25731 22185 25740 22219
rect 25688 22176 25740 22185
rect 25780 22176 25832 22228
rect 26148 22176 26200 22228
rect 29736 22176 29788 22228
rect 30840 22219 30892 22228
rect 30840 22185 30849 22219
rect 30849 22185 30883 22219
rect 30883 22185 30892 22219
rect 30840 22176 30892 22185
rect 33508 22176 33560 22228
rect 20352 22040 20404 22092
rect 29644 22083 29696 22092
rect 1860 22015 1912 22024
rect 1860 21981 1869 22015
rect 1869 21981 1903 22015
rect 1903 21981 1912 22015
rect 1860 21972 1912 21981
rect 2504 21972 2556 22024
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 11520 21972 11572 22024
rect 11244 21904 11296 21956
rect 16212 22015 16264 22024
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 17040 22015 17092 22024
rect 16212 21972 16264 21981
rect 17040 21981 17049 22015
rect 17049 21981 17083 22015
rect 17083 21981 17092 22015
rect 17040 21972 17092 21981
rect 18052 22015 18104 22024
rect 15936 21904 15988 21956
rect 18052 21981 18061 22015
rect 18061 21981 18095 22015
rect 18095 21981 18104 22015
rect 18052 21972 18104 21981
rect 18236 22015 18288 22024
rect 18236 21981 18245 22015
rect 18245 21981 18279 22015
rect 18279 21981 18288 22015
rect 18236 21972 18288 21981
rect 18604 21972 18656 22024
rect 18696 21972 18748 22024
rect 22468 22015 22520 22024
rect 2688 21879 2740 21888
rect 2688 21845 2697 21879
rect 2697 21845 2731 21879
rect 2731 21845 2740 21879
rect 2688 21836 2740 21845
rect 17224 21836 17276 21888
rect 21732 21904 21784 21956
rect 22468 21981 22477 22015
rect 22477 21981 22511 22015
rect 22511 21981 22520 22015
rect 29644 22049 29653 22083
rect 29653 22049 29687 22083
rect 29687 22049 29696 22083
rect 29644 22040 29696 22049
rect 32496 22040 32548 22092
rect 22468 21972 22520 21981
rect 23112 21972 23164 22024
rect 22192 21836 22244 21888
rect 24676 21972 24728 22024
rect 25044 21972 25096 22024
rect 29736 22015 29788 22024
rect 25136 21904 25188 21956
rect 29736 21981 29745 22015
rect 29745 21981 29779 22015
rect 29779 21981 29788 22015
rect 29736 21972 29788 21981
rect 31024 22015 31076 22024
rect 31024 21981 31033 22015
rect 31033 21981 31067 22015
rect 31067 21981 31076 22015
rect 31024 21972 31076 21981
rect 31208 22015 31260 22024
rect 31208 21981 31217 22015
rect 31217 21981 31251 22015
rect 31251 21981 31260 22015
rect 31208 21972 31260 21981
rect 31300 22015 31352 22024
rect 31300 21981 31309 22015
rect 31309 21981 31343 22015
rect 31343 21981 31352 22015
rect 31300 21972 31352 21981
rect 33508 21972 33560 22024
rect 34428 21972 34480 22024
rect 25044 21836 25096 21888
rect 30104 21904 30156 21956
rect 31852 21947 31904 21956
rect 31852 21913 31861 21947
rect 31861 21913 31895 21947
rect 31895 21913 31904 21947
rect 31852 21904 31904 21913
rect 31944 21904 31996 21956
rect 25412 21836 25464 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 7656 21675 7708 21684
rect 2688 21564 2740 21616
rect 7656 21641 7665 21675
rect 7665 21641 7699 21675
rect 7699 21641 7708 21675
rect 7656 21632 7708 21641
rect 10876 21675 10928 21684
rect 10876 21641 10885 21675
rect 10885 21641 10919 21675
rect 10919 21641 10928 21675
rect 10876 21632 10928 21641
rect 16856 21632 16908 21684
rect 21732 21632 21784 21684
rect 22192 21675 22244 21684
rect 22192 21641 22201 21675
rect 22201 21641 22235 21675
rect 22235 21641 22244 21675
rect 22192 21632 22244 21641
rect 26148 21675 26200 21684
rect 4896 21607 4948 21616
rect 4896 21573 4905 21607
rect 4905 21573 4939 21607
rect 4939 21573 4948 21607
rect 4896 21564 4948 21573
rect 8300 21564 8352 21616
rect 10600 21564 10652 21616
rect 15660 21564 15712 21616
rect 18052 21564 18104 21616
rect 10140 21496 10192 21548
rect 13820 21496 13872 21548
rect 14372 21496 14424 21548
rect 15752 21496 15804 21548
rect 17224 21496 17276 21548
rect 17960 21496 18012 21548
rect 18144 21496 18196 21548
rect 18880 21564 18932 21616
rect 18512 21539 18564 21548
rect 18512 21505 18521 21539
rect 18521 21505 18555 21539
rect 18555 21505 18564 21539
rect 22100 21564 22152 21616
rect 24952 21607 25004 21616
rect 18512 21496 18564 21505
rect 8944 21428 8996 21480
rect 9496 21471 9548 21480
rect 9496 21437 9505 21471
rect 9505 21437 9539 21471
rect 9539 21437 9548 21471
rect 9496 21428 9548 21437
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 2688 21292 2740 21344
rect 3792 21292 3844 21344
rect 4068 21335 4120 21344
rect 4068 21301 4077 21335
rect 4077 21301 4111 21335
rect 4111 21301 4120 21335
rect 4068 21292 4120 21301
rect 5264 21335 5316 21344
rect 5264 21301 5273 21335
rect 5273 21301 5307 21335
rect 5307 21301 5316 21335
rect 5264 21292 5316 21301
rect 7288 21335 7340 21344
rect 7288 21301 7297 21335
rect 7297 21301 7331 21335
rect 7331 21301 7340 21335
rect 7288 21292 7340 21301
rect 11612 21292 11664 21344
rect 14188 21335 14240 21344
rect 14188 21301 14197 21335
rect 14197 21301 14231 21335
rect 14231 21301 14240 21335
rect 14188 21292 14240 21301
rect 15936 21292 15988 21344
rect 16396 21292 16448 21344
rect 16580 21292 16632 21344
rect 17592 21471 17644 21480
rect 17592 21437 17601 21471
rect 17601 21437 17635 21471
rect 17635 21437 17644 21471
rect 18328 21471 18380 21480
rect 17592 21428 17644 21437
rect 18328 21437 18337 21471
rect 18337 21437 18371 21471
rect 18371 21437 18380 21471
rect 18328 21428 18380 21437
rect 18604 21471 18656 21480
rect 18604 21437 18613 21471
rect 18613 21437 18647 21471
rect 18647 21437 18656 21471
rect 18604 21428 18656 21437
rect 21180 21428 21232 21480
rect 24676 21496 24728 21548
rect 24952 21573 24993 21607
rect 24993 21573 25004 21607
rect 24952 21564 25004 21573
rect 25412 21564 25464 21616
rect 25044 21428 25096 21480
rect 26148 21641 26157 21675
rect 26157 21641 26191 21675
rect 26191 21641 26200 21675
rect 26148 21632 26200 21641
rect 29736 21632 29788 21684
rect 31024 21632 31076 21684
rect 32496 21675 32548 21684
rect 32496 21641 32505 21675
rect 32505 21641 32539 21675
rect 32539 21641 32548 21675
rect 32496 21632 32548 21641
rect 26056 21564 26108 21616
rect 31300 21564 31352 21616
rect 31944 21564 31996 21616
rect 27896 21539 27948 21548
rect 27896 21505 27930 21539
rect 27930 21505 27948 21539
rect 29460 21539 29512 21548
rect 27896 21496 27948 21505
rect 29460 21505 29469 21539
rect 29469 21505 29503 21539
rect 29503 21505 29512 21539
rect 29460 21496 29512 21505
rect 29552 21496 29604 21548
rect 31852 21496 31904 21548
rect 27620 21471 27672 21480
rect 27620 21437 27629 21471
rect 27629 21437 27663 21471
rect 27663 21437 27672 21471
rect 27620 21428 27672 21437
rect 34796 21496 34848 21548
rect 33324 21428 33376 21480
rect 17224 21360 17276 21412
rect 23940 21360 23992 21412
rect 17868 21292 17920 21344
rect 19432 21292 19484 21344
rect 24492 21292 24544 21344
rect 25596 21360 25648 21412
rect 25136 21335 25188 21344
rect 25136 21301 25145 21335
rect 25145 21301 25179 21335
rect 25179 21301 25188 21335
rect 25136 21292 25188 21301
rect 25320 21292 25372 21344
rect 25872 21292 25924 21344
rect 29184 21292 29236 21344
rect 35440 21292 35492 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2504 21131 2556 21140
rect 2504 21097 2513 21131
rect 2513 21097 2547 21131
rect 2547 21097 2556 21131
rect 2504 21088 2556 21097
rect 7656 21131 7708 21140
rect 7656 21097 7665 21131
rect 7665 21097 7699 21131
rect 7699 21097 7708 21131
rect 7656 21088 7708 21097
rect 10140 21131 10192 21140
rect 10140 21097 10149 21131
rect 10149 21097 10183 21131
rect 10183 21097 10192 21131
rect 10140 21088 10192 21097
rect 17224 21088 17276 21140
rect 17960 21088 18012 21140
rect 18696 21088 18748 21140
rect 19248 21131 19300 21140
rect 19248 21097 19257 21131
rect 19257 21097 19291 21131
rect 19291 21097 19300 21131
rect 19248 21088 19300 21097
rect 19340 21088 19392 21140
rect 27896 21131 27948 21140
rect 13452 21020 13504 21072
rect 2964 20995 3016 21004
rect 2964 20961 2973 20995
rect 2973 20961 3007 20995
rect 3007 20961 3016 20995
rect 2964 20952 3016 20961
rect 3148 20995 3200 21004
rect 3148 20961 3157 20995
rect 3157 20961 3191 20995
rect 3191 20961 3200 20995
rect 3148 20952 3200 20961
rect 4068 20884 4120 20936
rect 1676 20859 1728 20868
rect 1676 20825 1685 20859
rect 1685 20825 1719 20859
rect 1719 20825 1728 20859
rect 1676 20816 1728 20825
rect 7288 20884 7340 20936
rect 13176 20952 13228 21004
rect 14648 20952 14700 21004
rect 16488 21020 16540 21072
rect 17132 21020 17184 21072
rect 17868 21020 17920 21072
rect 16580 20952 16632 21004
rect 17592 20952 17644 21004
rect 19432 20995 19484 21004
rect 19432 20961 19441 20995
rect 19441 20961 19475 20995
rect 19475 20961 19484 20995
rect 19432 20952 19484 20961
rect 27896 21097 27905 21131
rect 27905 21097 27939 21131
rect 27939 21097 27948 21131
rect 27896 21088 27948 21097
rect 19800 21020 19852 21072
rect 30196 21020 30248 21072
rect 33692 21020 33744 21072
rect 31944 20952 31996 21004
rect 33048 20952 33100 21004
rect 33600 20995 33652 21004
rect 33600 20961 33609 20995
rect 33609 20961 33643 20995
rect 33643 20961 33652 20995
rect 33600 20952 33652 20961
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10643 20927
rect 10643 20893 10652 20927
rect 10600 20884 10652 20893
rect 7104 20816 7156 20868
rect 10876 20816 10928 20868
rect 11520 20884 11572 20936
rect 13360 20884 13412 20936
rect 13544 20927 13596 20936
rect 13544 20893 13553 20927
rect 13553 20893 13587 20927
rect 13587 20893 13596 20927
rect 13544 20884 13596 20893
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 14372 20927 14424 20936
rect 14372 20893 14382 20927
rect 14382 20893 14416 20927
rect 14416 20893 14424 20927
rect 14372 20884 14424 20893
rect 15292 20927 15344 20936
rect 13636 20816 13688 20868
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 15568 20927 15620 20936
rect 15568 20893 15577 20927
rect 15577 20893 15611 20927
rect 15611 20893 15620 20927
rect 15568 20884 15620 20893
rect 17960 20927 18012 20936
rect 17960 20893 17969 20927
rect 17969 20893 18003 20927
rect 18003 20893 18012 20927
rect 17960 20884 18012 20893
rect 15936 20816 15988 20868
rect 18236 20927 18288 20936
rect 18236 20893 18245 20927
rect 18245 20893 18279 20927
rect 18279 20893 18288 20927
rect 18236 20884 18288 20893
rect 19340 20884 19392 20936
rect 19524 20927 19576 20936
rect 19524 20893 19533 20927
rect 19533 20893 19567 20927
rect 19567 20893 19576 20927
rect 19524 20884 19576 20893
rect 25136 20884 25188 20936
rect 28172 20884 28224 20936
rect 28540 20884 28592 20936
rect 29092 20884 29144 20936
rect 29460 20884 29512 20936
rect 33324 20927 33376 20936
rect 33324 20893 33333 20927
rect 33333 20893 33367 20927
rect 33367 20893 33376 20927
rect 33324 20884 33376 20893
rect 33508 20927 33560 20936
rect 33508 20893 33517 20927
rect 33517 20893 33551 20927
rect 33551 20893 33560 20927
rect 33508 20884 33560 20893
rect 33692 20884 33744 20936
rect 11152 20748 11204 20800
rect 12072 20748 12124 20800
rect 13084 20791 13136 20800
rect 13084 20757 13093 20791
rect 13093 20757 13127 20791
rect 13127 20757 13136 20791
rect 13084 20748 13136 20757
rect 13452 20791 13504 20800
rect 13452 20757 13461 20791
rect 13461 20757 13495 20791
rect 13495 20757 13504 20791
rect 13452 20748 13504 20757
rect 14188 20748 14240 20800
rect 14556 20748 14608 20800
rect 25688 20748 25740 20800
rect 30380 20816 30432 20868
rect 31208 20816 31260 20868
rect 31668 20816 31720 20868
rect 32772 20748 32824 20800
rect 33140 20791 33192 20800
rect 33140 20757 33149 20791
rect 33149 20757 33183 20791
rect 33183 20757 33192 20791
rect 33140 20748 33192 20757
rect 33876 20816 33928 20868
rect 35440 20927 35492 20936
rect 35440 20893 35474 20927
rect 35474 20893 35492 20927
rect 35440 20884 35492 20893
rect 35716 20884 35768 20936
rect 37648 20927 37700 20936
rect 37648 20893 37657 20927
rect 37657 20893 37691 20927
rect 37691 20893 37700 20927
rect 37648 20884 37700 20893
rect 37740 20816 37792 20868
rect 35716 20748 35768 20800
rect 37372 20748 37424 20800
rect 37464 20748 37516 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 8208 20476 8260 20528
rect 13452 20544 13504 20596
rect 14648 20544 14700 20596
rect 15292 20544 15344 20596
rect 13084 20476 13136 20528
rect 3700 20408 3752 20460
rect 3884 20451 3936 20460
rect 3884 20417 3893 20451
rect 3893 20417 3927 20451
rect 3927 20417 3936 20451
rect 3884 20408 3936 20417
rect 7840 20408 7892 20460
rect 12164 20408 12216 20460
rect 12348 20408 12400 20460
rect 14280 20408 14332 20460
rect 15292 20408 15344 20460
rect 16304 20544 16356 20596
rect 17960 20544 18012 20596
rect 18696 20544 18748 20596
rect 33692 20587 33744 20596
rect 33692 20553 33701 20587
rect 33701 20553 33735 20587
rect 33735 20553 33744 20587
rect 33692 20544 33744 20553
rect 33876 20587 33928 20596
rect 33876 20553 33885 20587
rect 33885 20553 33919 20587
rect 33919 20553 33928 20587
rect 33876 20544 33928 20553
rect 34796 20544 34848 20596
rect 23756 20476 23808 20528
rect 15936 20451 15988 20460
rect 15936 20417 15945 20451
rect 15945 20417 15979 20451
rect 15979 20417 15988 20451
rect 15936 20408 15988 20417
rect 17500 20408 17552 20460
rect 18236 20408 18288 20460
rect 3148 20383 3200 20392
rect 3148 20349 3157 20383
rect 3157 20349 3191 20383
rect 3191 20349 3200 20383
rect 3148 20340 3200 20349
rect 7104 20383 7156 20392
rect 7104 20349 7113 20383
rect 7113 20349 7147 20383
rect 7147 20349 7156 20383
rect 7104 20340 7156 20349
rect 15752 20383 15804 20392
rect 15752 20349 15761 20383
rect 15761 20349 15795 20383
rect 15795 20349 15804 20383
rect 15752 20340 15804 20349
rect 16948 20340 17000 20392
rect 18696 20340 18748 20392
rect 18880 20451 18932 20460
rect 18880 20417 18889 20451
rect 18889 20417 18923 20451
rect 18923 20417 18932 20451
rect 18880 20408 18932 20417
rect 19984 20408 20036 20460
rect 20720 20408 20772 20460
rect 23112 20408 23164 20460
rect 23296 20451 23348 20460
rect 23296 20417 23330 20451
rect 23330 20417 23348 20451
rect 23296 20408 23348 20417
rect 18972 20383 19024 20392
rect 18972 20349 18981 20383
rect 18981 20349 19015 20383
rect 19015 20349 19024 20383
rect 18972 20340 19024 20349
rect 18604 20272 18656 20324
rect 25136 20476 25188 20528
rect 26056 20476 26108 20528
rect 28448 20476 28500 20528
rect 28908 20519 28960 20528
rect 28908 20485 28933 20519
rect 28933 20485 28960 20519
rect 28908 20476 28960 20485
rect 32680 20519 32732 20528
rect 32680 20485 32689 20519
rect 32689 20485 32723 20519
rect 32723 20485 32732 20519
rect 32680 20476 32732 20485
rect 33600 20476 33652 20528
rect 37372 20476 37424 20528
rect 37740 20476 37792 20528
rect 25688 20451 25740 20460
rect 25688 20417 25697 20451
rect 25697 20417 25731 20451
rect 25731 20417 25740 20451
rect 25688 20408 25740 20417
rect 31668 20408 31720 20460
rect 31760 20408 31812 20460
rect 24492 20272 24544 20324
rect 28816 20272 28868 20324
rect 29092 20315 29144 20324
rect 29092 20281 29101 20315
rect 29101 20281 29135 20315
rect 29135 20281 29144 20315
rect 29092 20272 29144 20281
rect 32956 20408 33008 20460
rect 33048 20408 33100 20460
rect 34520 20451 34572 20460
rect 34520 20417 34529 20451
rect 34529 20417 34563 20451
rect 34563 20417 34572 20451
rect 34520 20408 34572 20417
rect 34704 20451 34756 20460
rect 34704 20417 34713 20451
rect 34713 20417 34747 20451
rect 34747 20417 34756 20451
rect 34704 20408 34756 20417
rect 33232 20340 33284 20392
rect 33600 20272 33652 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 2780 20204 2832 20256
rect 18972 20204 19024 20256
rect 21088 20204 21140 20256
rect 21916 20204 21968 20256
rect 28632 20204 28684 20256
rect 28908 20247 28960 20256
rect 28908 20213 28917 20247
rect 28917 20213 28951 20247
rect 28951 20213 28960 20247
rect 28908 20204 28960 20213
rect 29000 20204 29052 20256
rect 33416 20204 33468 20256
rect 34060 20247 34112 20256
rect 34060 20213 34069 20247
rect 34069 20213 34103 20247
rect 34103 20213 34112 20247
rect 34060 20204 34112 20213
rect 38016 20204 38068 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7840 20043 7892 20052
rect 7840 20009 7849 20043
rect 7849 20009 7883 20043
rect 7883 20009 7892 20043
rect 7840 20000 7892 20009
rect 2596 19932 2648 19984
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 2780 19839 2832 19848
rect 2780 19805 2789 19839
rect 2789 19805 2823 19839
rect 2823 19805 2832 19839
rect 5080 19839 5132 19848
rect 2780 19796 2832 19805
rect 5080 19805 5089 19839
rect 5089 19805 5123 19839
rect 5123 19805 5132 19839
rect 5080 19796 5132 19805
rect 16672 19932 16724 19984
rect 8116 19864 8168 19916
rect 11428 19864 11480 19916
rect 11520 19864 11572 19916
rect 8300 19839 8352 19848
rect 8300 19805 8309 19839
rect 8309 19805 8343 19839
rect 8343 19805 8352 19839
rect 8300 19796 8352 19805
rect 2044 19728 2096 19780
rect 11244 19796 11296 19848
rect 13544 19864 13596 19916
rect 15292 19907 15344 19916
rect 11612 19728 11664 19780
rect 14464 19796 14516 19848
rect 14832 19796 14884 19848
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 16580 19907 16632 19916
rect 16304 19839 16356 19848
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 16580 19873 16589 19907
rect 16589 19873 16623 19907
rect 16623 19873 16632 19907
rect 16580 19864 16632 19873
rect 16948 19728 17000 19780
rect 1768 19660 1820 19712
rect 2596 19703 2648 19712
rect 2596 19669 2605 19703
rect 2605 19669 2639 19703
rect 2639 19669 2648 19703
rect 2596 19660 2648 19669
rect 4896 19703 4948 19712
rect 4896 19669 4905 19703
rect 4905 19669 4939 19703
rect 4939 19669 4948 19703
rect 4896 19660 4948 19669
rect 8208 19703 8260 19712
rect 8208 19669 8217 19703
rect 8217 19669 8251 19703
rect 8251 19669 8260 19703
rect 8208 19660 8260 19669
rect 9680 19703 9732 19712
rect 9680 19669 9689 19703
rect 9689 19669 9723 19703
rect 9723 19669 9732 19703
rect 9680 19660 9732 19669
rect 9772 19660 9824 19712
rect 11244 19660 11296 19712
rect 15752 19660 15804 19712
rect 18328 20000 18380 20052
rect 18696 20000 18748 20052
rect 18880 20000 18932 20052
rect 20720 20043 20772 20052
rect 20720 20009 20729 20043
rect 20729 20009 20763 20043
rect 20763 20009 20772 20043
rect 20720 20000 20772 20009
rect 21456 20000 21508 20052
rect 22008 20043 22060 20052
rect 22008 20009 22017 20043
rect 22017 20009 22051 20043
rect 22051 20009 22060 20043
rect 22008 20000 22060 20009
rect 22100 20000 22152 20052
rect 23296 20000 23348 20052
rect 24676 20000 24728 20052
rect 17684 19932 17736 19984
rect 28540 20000 28592 20052
rect 28816 20000 28868 20052
rect 30104 20043 30156 20052
rect 29000 19932 29052 19984
rect 30104 20009 30113 20043
rect 30113 20009 30147 20043
rect 30147 20009 30156 20043
rect 30104 20000 30156 20009
rect 30196 20000 30248 20052
rect 33416 20000 33468 20052
rect 37464 20000 37516 20052
rect 37648 20000 37700 20052
rect 34704 19932 34756 19984
rect 18052 19864 18104 19916
rect 20720 19864 20772 19916
rect 17500 19796 17552 19848
rect 18604 19796 18656 19848
rect 22192 19864 22244 19916
rect 21088 19839 21140 19848
rect 21088 19805 21097 19839
rect 21097 19805 21131 19839
rect 21131 19805 21140 19839
rect 21088 19796 21140 19805
rect 21180 19839 21232 19848
rect 21180 19805 21189 19839
rect 21189 19805 21223 19839
rect 21223 19805 21232 19839
rect 23664 19864 23716 19916
rect 24492 19864 24544 19916
rect 28448 19864 28500 19916
rect 21180 19796 21232 19805
rect 23756 19839 23808 19848
rect 23756 19805 23765 19839
rect 23765 19805 23799 19839
rect 23799 19805 23808 19839
rect 23756 19796 23808 19805
rect 23848 19839 23900 19848
rect 23848 19805 23857 19839
rect 23857 19805 23891 19839
rect 23891 19805 23900 19839
rect 23848 19796 23900 19805
rect 27620 19796 27672 19848
rect 29184 19864 29236 19916
rect 29736 19864 29788 19916
rect 28816 19796 28868 19848
rect 21456 19771 21508 19780
rect 21456 19737 21465 19771
rect 21465 19737 21499 19771
rect 21499 19737 21508 19771
rect 21456 19728 21508 19737
rect 21824 19771 21876 19780
rect 21824 19737 21833 19771
rect 21833 19737 21867 19771
rect 21867 19737 21876 19771
rect 21824 19728 21876 19737
rect 22100 19728 22152 19780
rect 21732 19660 21784 19712
rect 24216 19660 24268 19712
rect 26976 19728 27028 19780
rect 31760 19839 31812 19848
rect 31760 19805 31769 19839
rect 31769 19805 31803 19839
rect 31803 19805 31812 19839
rect 31760 19796 31812 19805
rect 31944 19839 31996 19848
rect 31944 19805 31951 19839
rect 31951 19805 31996 19839
rect 31944 19796 31996 19805
rect 29552 19771 29604 19780
rect 27068 19660 27120 19712
rect 28540 19660 28592 19712
rect 29552 19737 29561 19771
rect 29561 19737 29595 19771
rect 29595 19737 29604 19771
rect 29552 19728 29604 19737
rect 29644 19728 29696 19780
rect 28908 19660 28960 19712
rect 29736 19703 29788 19712
rect 29736 19669 29745 19703
rect 29745 19669 29779 19703
rect 29779 19669 29788 19703
rect 29736 19660 29788 19669
rect 32220 19660 32272 19712
rect 32680 19864 32732 19916
rect 32864 19839 32916 19848
rect 32864 19805 32873 19839
rect 32873 19805 32907 19839
rect 32907 19805 32916 19839
rect 32864 19796 32916 19805
rect 33692 19864 33744 19916
rect 36912 19839 36964 19848
rect 33232 19771 33284 19780
rect 33232 19737 33241 19771
rect 33241 19737 33275 19771
rect 33275 19737 33284 19771
rect 33232 19728 33284 19737
rect 32680 19660 32732 19712
rect 32864 19660 32916 19712
rect 33048 19660 33100 19712
rect 36912 19805 36921 19839
rect 36921 19805 36955 19839
rect 36955 19805 36964 19839
rect 36912 19796 36964 19805
rect 37740 19839 37792 19848
rect 37740 19805 37749 19839
rect 37749 19805 37783 19839
rect 37783 19805 37792 19839
rect 37740 19796 37792 19805
rect 38292 19796 38344 19848
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 3700 19456 3752 19508
rect 7196 19456 7248 19508
rect 2596 19388 2648 19440
rect 4896 19388 4948 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 1492 19252 1544 19304
rect 2504 19252 2556 19304
rect 2688 19320 2740 19372
rect 7104 19320 7156 19372
rect 8208 19320 8260 19372
rect 9496 19320 9548 19372
rect 9864 19363 9916 19372
rect 9864 19329 9898 19363
rect 9898 19329 9916 19363
rect 11428 19456 11480 19508
rect 12072 19456 12124 19508
rect 13912 19456 13964 19508
rect 14464 19456 14516 19508
rect 9864 19320 9916 19329
rect 12808 19320 12860 19372
rect 13728 19320 13780 19372
rect 15200 19363 15252 19372
rect 13820 19252 13872 19304
rect 14188 19295 14240 19304
rect 14188 19261 14198 19295
rect 14198 19261 14232 19295
rect 14232 19261 14240 19295
rect 14188 19252 14240 19261
rect 14464 19295 14516 19304
rect 14464 19261 14473 19295
rect 14473 19261 14507 19295
rect 14507 19261 14516 19295
rect 15200 19329 15209 19363
rect 15209 19329 15243 19363
rect 15243 19329 15252 19363
rect 15200 19320 15252 19329
rect 15568 19456 15620 19508
rect 17408 19456 17460 19508
rect 15752 19320 15804 19372
rect 20628 19388 20680 19440
rect 20812 19388 20864 19440
rect 21824 19431 21876 19440
rect 21824 19397 21833 19431
rect 21833 19397 21867 19431
rect 21867 19397 21876 19431
rect 21824 19388 21876 19397
rect 22192 19499 22244 19508
rect 22192 19465 22201 19499
rect 22201 19465 22235 19499
rect 22235 19465 22244 19499
rect 22192 19456 22244 19465
rect 23848 19456 23900 19508
rect 26976 19499 27028 19508
rect 26976 19465 26985 19499
rect 26985 19465 27019 19499
rect 27019 19465 27028 19499
rect 26976 19456 27028 19465
rect 27068 19456 27120 19508
rect 21916 19320 21968 19372
rect 22100 19320 22152 19372
rect 24216 19363 24268 19372
rect 24216 19329 24225 19363
rect 24225 19329 24259 19363
rect 24259 19329 24268 19363
rect 24216 19320 24268 19329
rect 28816 19388 28868 19440
rect 29552 19388 29604 19440
rect 27988 19363 28040 19372
rect 27988 19329 27997 19363
rect 27997 19329 28031 19363
rect 28031 19329 28040 19363
rect 27988 19320 28040 19329
rect 14464 19252 14516 19261
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 16304 19252 16356 19304
rect 17592 19252 17644 19304
rect 18512 19295 18564 19304
rect 18512 19261 18522 19295
rect 18522 19261 18556 19295
rect 18556 19261 18564 19295
rect 18512 19252 18564 19261
rect 18696 19295 18748 19304
rect 18696 19261 18705 19295
rect 18705 19261 18739 19295
rect 18739 19261 18748 19295
rect 18696 19252 18748 19261
rect 18972 19252 19024 19304
rect 27160 19295 27212 19304
rect 27160 19261 27169 19295
rect 27169 19261 27203 19295
rect 27203 19261 27212 19295
rect 27160 19252 27212 19261
rect 28540 19320 28592 19372
rect 28908 19363 28960 19372
rect 28908 19329 28917 19363
rect 28917 19329 28951 19363
rect 28951 19329 28960 19363
rect 28908 19320 28960 19329
rect 32864 19388 32916 19440
rect 33140 19456 33192 19508
rect 34520 19456 34572 19508
rect 37740 19388 37792 19440
rect 20628 19184 20680 19236
rect 24216 19184 24268 19236
rect 31852 19252 31904 19304
rect 32496 19363 32548 19372
rect 32496 19329 32505 19363
rect 32505 19329 32539 19363
rect 32539 19329 32548 19363
rect 32496 19320 32548 19329
rect 32680 19320 32732 19372
rect 33048 19320 33100 19372
rect 34060 19320 34112 19372
rect 34428 19320 34480 19372
rect 44088 19363 44140 19372
rect 44088 19329 44097 19363
rect 44097 19329 44131 19363
rect 44131 19329 44140 19363
rect 44088 19320 44140 19329
rect 32956 19252 33008 19304
rect 35440 19252 35492 19304
rect 38016 19252 38068 19304
rect 38292 19252 38344 19304
rect 30380 19184 30432 19236
rect 32588 19184 32640 19236
rect 32772 19227 32824 19236
rect 32772 19193 32781 19227
rect 32781 19193 32815 19227
rect 32815 19193 32824 19227
rect 32772 19184 32824 19193
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 6000 19116 6052 19168
rect 14280 19116 14332 19168
rect 16396 19116 16448 19168
rect 19064 19116 19116 19168
rect 21640 19116 21692 19168
rect 26884 19116 26936 19168
rect 32680 19116 32732 19168
rect 33692 19159 33744 19168
rect 33692 19125 33701 19159
rect 33701 19125 33735 19159
rect 33735 19125 33744 19159
rect 33692 19116 33744 19125
rect 43904 19159 43956 19168
rect 43904 19125 43913 19159
rect 43913 19125 43947 19159
rect 43947 19125 43956 19159
rect 43904 19116 43956 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1400 18912 1452 18964
rect 2688 18912 2740 18964
rect 5080 18912 5132 18964
rect 13084 18912 13136 18964
rect 13176 18912 13228 18964
rect 15476 18912 15528 18964
rect 15660 18955 15712 18964
rect 15660 18921 15669 18955
rect 15669 18921 15703 18955
rect 15703 18921 15712 18955
rect 15660 18912 15712 18921
rect 15936 18912 15988 18964
rect 16120 18912 16172 18964
rect 20996 18912 21048 18964
rect 27160 18912 27212 18964
rect 32680 18912 32732 18964
rect 37280 18912 37332 18964
rect 9864 18887 9916 18896
rect 1492 18776 1544 18828
rect 1676 18708 1728 18760
rect 9864 18853 9873 18887
rect 9873 18853 9907 18887
rect 9907 18853 9916 18887
rect 9864 18844 9916 18853
rect 15844 18887 15896 18896
rect 15844 18853 15853 18887
rect 15853 18853 15887 18887
rect 15887 18853 15896 18887
rect 15844 18844 15896 18853
rect 6736 18776 6788 18828
rect 14924 18776 14976 18828
rect 15292 18776 15344 18828
rect 27712 18844 27764 18896
rect 27804 18844 27856 18896
rect 33692 18844 33744 18896
rect 37832 18844 37884 18896
rect 38568 18844 38620 18896
rect 3976 18751 4028 18760
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 9680 18708 9732 18760
rect 11428 18751 11480 18760
rect 11428 18717 11437 18751
rect 11437 18717 11471 18751
rect 11471 18717 11480 18751
rect 11428 18708 11480 18717
rect 12164 18708 12216 18760
rect 16120 18708 16172 18760
rect 16856 18751 16908 18760
rect 16856 18717 16865 18751
rect 16865 18717 16899 18751
rect 16899 18717 16908 18751
rect 16856 18708 16908 18717
rect 18144 18708 18196 18760
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 2320 18640 2372 18692
rect 12624 18640 12676 18692
rect 6000 18572 6052 18624
rect 6920 18615 6972 18624
rect 6920 18581 6929 18615
rect 6929 18581 6963 18615
rect 6963 18581 6972 18615
rect 6920 18572 6972 18581
rect 7564 18572 7616 18624
rect 15016 18683 15068 18692
rect 15016 18649 15025 18683
rect 15025 18649 15059 18683
rect 15059 18649 15068 18683
rect 15016 18640 15068 18649
rect 15292 18640 15344 18692
rect 12992 18572 13044 18624
rect 13268 18572 13320 18624
rect 15844 18640 15896 18692
rect 16304 18640 16356 18692
rect 16396 18640 16448 18692
rect 17500 18640 17552 18692
rect 16028 18572 16080 18624
rect 18512 18819 18564 18828
rect 18512 18785 18521 18819
rect 18521 18785 18555 18819
rect 18555 18785 18564 18819
rect 18512 18776 18564 18785
rect 18972 18776 19024 18828
rect 19064 18776 19116 18828
rect 26884 18776 26936 18828
rect 28816 18776 28868 18828
rect 18512 18640 18564 18692
rect 19984 18708 20036 18760
rect 27252 18708 27304 18760
rect 28908 18708 28960 18760
rect 29000 18708 29052 18760
rect 29644 18708 29696 18760
rect 32588 18751 32640 18760
rect 32588 18717 32597 18751
rect 32597 18717 32631 18751
rect 32631 18717 32640 18751
rect 32588 18708 32640 18717
rect 35440 18776 35492 18828
rect 33048 18751 33100 18760
rect 33048 18717 33062 18751
rect 33062 18717 33096 18751
rect 33096 18717 33100 18751
rect 36636 18751 36688 18760
rect 33048 18708 33100 18717
rect 36636 18717 36645 18751
rect 36645 18717 36679 18751
rect 36679 18717 36688 18751
rect 36636 18708 36688 18717
rect 36912 18751 36964 18760
rect 36912 18717 36921 18751
rect 36921 18717 36955 18751
rect 36955 18717 36964 18751
rect 36912 18708 36964 18717
rect 37188 18708 37240 18760
rect 43076 18751 43128 18760
rect 18972 18640 19024 18692
rect 23664 18640 23716 18692
rect 27160 18683 27212 18692
rect 27160 18649 27169 18683
rect 27169 18649 27203 18683
rect 27203 18649 27212 18683
rect 27160 18640 27212 18649
rect 27988 18640 28040 18692
rect 32864 18683 32916 18692
rect 32864 18649 32873 18683
rect 32873 18649 32907 18683
rect 32907 18649 32916 18683
rect 32864 18640 32916 18649
rect 43076 18717 43085 18751
rect 43085 18717 43119 18751
rect 43119 18717 43128 18751
rect 43076 18708 43128 18717
rect 43904 18708 43956 18760
rect 47492 18751 47544 18760
rect 47492 18717 47501 18751
rect 47501 18717 47535 18751
rect 47535 18717 47544 18751
rect 47492 18708 47544 18717
rect 30196 18572 30248 18624
rect 33048 18572 33100 18624
rect 37832 18572 37884 18624
rect 38292 18615 38344 18624
rect 38292 18581 38301 18615
rect 38301 18581 38335 18615
rect 38335 18581 38344 18615
rect 39212 18640 39264 18692
rect 38936 18615 38988 18624
rect 38292 18572 38344 18581
rect 38936 18581 38945 18615
rect 38945 18581 38979 18615
rect 38979 18581 38988 18615
rect 38936 18572 38988 18581
rect 44364 18572 44416 18624
rect 47308 18615 47360 18624
rect 47308 18581 47317 18615
rect 47317 18581 47351 18615
rect 47351 18581 47360 18615
rect 47308 18572 47360 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 1676 18368 1728 18420
rect 2320 18411 2372 18420
rect 2320 18377 2329 18411
rect 2329 18377 2363 18411
rect 2363 18377 2372 18411
rect 2320 18368 2372 18377
rect 2688 18411 2740 18420
rect 2688 18377 2697 18411
rect 2697 18377 2731 18411
rect 2731 18377 2740 18411
rect 2688 18368 2740 18377
rect 1952 18300 2004 18352
rect 7564 18368 7616 18420
rect 12624 18411 12676 18420
rect 12624 18377 12633 18411
rect 12633 18377 12667 18411
rect 12667 18377 12676 18411
rect 12624 18368 12676 18377
rect 15200 18368 15252 18420
rect 15292 18368 15344 18420
rect 15476 18368 15528 18420
rect 6920 18300 6972 18352
rect 12992 18343 13044 18352
rect 12992 18309 13001 18343
rect 13001 18309 13035 18343
rect 13035 18309 13044 18343
rect 18236 18368 18288 18420
rect 18420 18368 18472 18420
rect 19340 18368 19392 18420
rect 20996 18411 21048 18420
rect 12992 18300 13044 18309
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 2596 18232 2648 18284
rect 2780 18275 2832 18284
rect 2780 18241 2789 18275
rect 2789 18241 2823 18275
rect 2823 18241 2832 18275
rect 3424 18275 3476 18284
rect 2780 18232 2832 18241
rect 3424 18241 3433 18275
rect 3433 18241 3467 18275
rect 3467 18241 3476 18275
rect 3424 18232 3476 18241
rect 6460 18232 6512 18284
rect 6920 18164 6972 18216
rect 8208 18232 8260 18284
rect 6736 18139 6788 18148
rect 6736 18105 6745 18139
rect 6745 18105 6779 18139
rect 6779 18105 6788 18139
rect 6736 18096 6788 18105
rect 6552 18028 6604 18080
rect 6828 18028 6880 18080
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 13544 18232 13596 18284
rect 13820 18232 13872 18284
rect 14832 18232 14884 18284
rect 16856 18232 16908 18284
rect 19984 18300 20036 18352
rect 18144 18232 18196 18284
rect 15660 18164 15712 18216
rect 16028 18164 16080 18216
rect 17592 18207 17644 18216
rect 16580 18096 16632 18148
rect 17592 18173 17601 18207
rect 17601 18173 17635 18207
rect 17635 18173 17644 18207
rect 17592 18164 17644 18173
rect 17684 18207 17736 18216
rect 17684 18173 17693 18207
rect 17693 18173 17727 18207
rect 17727 18173 17736 18207
rect 18512 18207 18564 18216
rect 17684 18164 17736 18173
rect 18512 18173 18521 18207
rect 18521 18173 18555 18207
rect 18555 18173 18564 18207
rect 18512 18164 18564 18173
rect 19340 18232 19392 18284
rect 20996 18377 21005 18411
rect 21005 18377 21039 18411
rect 21039 18377 21048 18411
rect 20996 18368 21048 18377
rect 20812 18343 20864 18352
rect 20812 18309 20821 18343
rect 20821 18309 20855 18343
rect 20855 18309 20864 18343
rect 20812 18300 20864 18309
rect 33876 18368 33928 18420
rect 22192 18343 22244 18352
rect 22192 18309 22201 18343
rect 22201 18309 22235 18343
rect 22235 18309 22244 18343
rect 22192 18300 22244 18309
rect 18420 18096 18472 18148
rect 18880 18164 18932 18216
rect 19064 18096 19116 18148
rect 21916 18232 21968 18284
rect 22376 18232 22428 18284
rect 24400 18232 24452 18284
rect 25320 18232 25372 18284
rect 27804 18300 27856 18352
rect 29184 18300 29236 18352
rect 27160 18232 27212 18284
rect 29460 18275 29512 18284
rect 29460 18241 29469 18275
rect 29469 18241 29503 18275
rect 29503 18241 29512 18275
rect 29460 18232 29512 18241
rect 29644 18275 29696 18284
rect 29644 18241 29651 18275
rect 29651 18241 29696 18275
rect 29644 18232 29696 18241
rect 29736 18275 29788 18284
rect 29736 18241 29745 18275
rect 29745 18241 29779 18275
rect 29779 18241 29788 18275
rect 29736 18232 29788 18241
rect 30012 18232 30064 18284
rect 32956 18300 33008 18352
rect 34796 18368 34848 18420
rect 35440 18411 35492 18420
rect 35440 18377 35449 18411
rect 35449 18377 35483 18411
rect 35483 18377 35492 18411
rect 35440 18368 35492 18377
rect 32864 18232 32916 18284
rect 33140 18232 33192 18284
rect 34060 18343 34112 18352
rect 34060 18309 34069 18343
rect 34069 18309 34103 18343
rect 34103 18309 34112 18343
rect 34060 18300 34112 18309
rect 19708 18207 19760 18216
rect 19708 18173 19717 18207
rect 19717 18173 19751 18207
rect 19751 18173 19760 18207
rect 23204 18207 23256 18216
rect 19708 18164 19760 18173
rect 23204 18173 23213 18207
rect 23213 18173 23247 18207
rect 23247 18173 23256 18207
rect 23204 18164 23256 18173
rect 24216 18164 24268 18216
rect 15016 18028 15068 18080
rect 15108 18028 15160 18080
rect 18144 18028 18196 18080
rect 18604 18028 18656 18080
rect 19156 18028 19208 18080
rect 19708 18028 19760 18080
rect 20720 18028 20772 18080
rect 21824 18071 21876 18080
rect 21824 18037 21833 18071
rect 21833 18037 21867 18071
rect 21867 18037 21876 18071
rect 21824 18028 21876 18037
rect 24584 18071 24636 18080
rect 24584 18037 24593 18071
rect 24593 18037 24627 18071
rect 24627 18037 24636 18071
rect 24584 18028 24636 18037
rect 28172 18096 28224 18148
rect 30380 18164 30432 18216
rect 32404 18207 32456 18216
rect 32404 18173 32413 18207
rect 32413 18173 32447 18207
rect 32447 18173 32456 18207
rect 32404 18164 32456 18173
rect 33600 18096 33652 18148
rect 34152 18275 34204 18284
rect 34152 18241 34166 18275
rect 34166 18241 34200 18275
rect 34200 18241 34204 18275
rect 34152 18232 34204 18241
rect 34428 18232 34480 18284
rect 35440 18232 35492 18284
rect 36636 18300 36688 18352
rect 43168 18368 43220 18420
rect 44088 18411 44140 18420
rect 44088 18377 44097 18411
rect 44097 18377 44131 18411
rect 44131 18377 44140 18411
rect 44088 18368 44140 18377
rect 55404 18411 55456 18420
rect 42616 18300 42668 18352
rect 37188 18232 37240 18284
rect 43076 18232 43128 18284
rect 46664 18275 46716 18284
rect 46664 18241 46673 18275
rect 46673 18241 46707 18275
rect 46707 18241 46716 18275
rect 46664 18232 46716 18241
rect 47308 18300 47360 18352
rect 55404 18377 55413 18411
rect 55413 18377 55447 18411
rect 55447 18377 55456 18411
rect 55404 18368 55456 18377
rect 47584 18275 47636 18284
rect 35900 18096 35952 18148
rect 37004 18164 37056 18216
rect 37280 18207 37332 18216
rect 37280 18173 37289 18207
rect 37289 18173 37323 18207
rect 37323 18173 37332 18207
rect 37280 18164 37332 18173
rect 27528 18028 27580 18080
rect 27712 18028 27764 18080
rect 36084 18028 36136 18080
rect 36544 18028 36596 18080
rect 43904 18071 43956 18080
rect 43904 18037 43913 18071
rect 43913 18037 43947 18071
rect 43947 18037 43956 18071
rect 43904 18028 43956 18037
rect 47032 18071 47084 18080
rect 47032 18037 47041 18071
rect 47041 18037 47075 18071
rect 47075 18037 47084 18071
rect 47032 18028 47084 18037
rect 47584 18241 47593 18275
rect 47593 18241 47627 18275
rect 47627 18241 47636 18275
rect 47584 18232 47636 18241
rect 53564 18275 53616 18284
rect 53564 18241 53573 18275
rect 53573 18241 53607 18275
rect 53607 18241 53616 18275
rect 53564 18232 53616 18241
rect 53380 18164 53432 18216
rect 47860 18028 47912 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 7104 17824 7156 17876
rect 8944 17824 8996 17876
rect 16672 17824 16724 17876
rect 16856 17824 16908 17876
rect 18880 17824 18932 17876
rect 18972 17824 19024 17876
rect 39212 17824 39264 17876
rect 14280 17756 14332 17808
rect 19984 17756 20036 17808
rect 22192 17756 22244 17808
rect 24400 17799 24452 17808
rect 24400 17765 24409 17799
rect 24409 17765 24443 17799
rect 24443 17765 24452 17799
rect 24400 17756 24452 17765
rect 27160 17756 27212 17808
rect 32404 17756 32456 17808
rect 2504 17688 2556 17740
rect 6552 17688 6604 17740
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 3792 17663 3844 17672
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 2320 17527 2372 17536
rect 2320 17493 2329 17527
rect 2329 17493 2363 17527
rect 2363 17493 2372 17527
rect 2320 17484 2372 17493
rect 3792 17629 3801 17663
rect 3801 17629 3835 17663
rect 3835 17629 3844 17663
rect 3792 17620 3844 17629
rect 6736 17620 6788 17672
rect 8300 17688 8352 17740
rect 8944 17731 8996 17740
rect 8944 17697 8953 17731
rect 8953 17697 8987 17731
rect 8987 17697 8996 17731
rect 8944 17688 8996 17697
rect 11428 17620 11480 17672
rect 12532 17620 12584 17672
rect 12992 17620 13044 17672
rect 13452 17620 13504 17672
rect 3884 17552 3936 17604
rect 5632 17552 5684 17604
rect 7840 17552 7892 17604
rect 13360 17552 13412 17604
rect 15936 17620 15988 17672
rect 16396 17688 16448 17740
rect 16488 17688 16540 17740
rect 16856 17620 16908 17672
rect 16948 17620 17000 17672
rect 17684 17688 17736 17740
rect 17776 17688 17828 17740
rect 20536 17688 20588 17740
rect 18972 17620 19024 17672
rect 20168 17620 20220 17672
rect 21824 17620 21876 17672
rect 24768 17620 24820 17672
rect 24952 17620 25004 17672
rect 15016 17552 15068 17604
rect 18788 17552 18840 17604
rect 18880 17552 18932 17604
rect 20904 17552 20956 17604
rect 25412 17552 25464 17604
rect 28908 17688 28960 17740
rect 27528 17620 27580 17672
rect 29092 17620 29144 17672
rect 29460 17620 29512 17672
rect 29736 17688 29788 17740
rect 30012 17663 30064 17672
rect 30012 17629 30026 17663
rect 30026 17629 30060 17663
rect 30060 17629 30064 17663
rect 30012 17620 30064 17629
rect 25964 17552 26016 17604
rect 26516 17552 26568 17604
rect 29828 17595 29880 17604
rect 4160 17484 4212 17536
rect 5816 17527 5868 17536
rect 5816 17493 5825 17527
rect 5825 17493 5859 17527
rect 5859 17493 5868 17527
rect 5816 17484 5868 17493
rect 6368 17484 6420 17536
rect 6828 17484 6880 17536
rect 10324 17527 10376 17536
rect 10324 17493 10333 17527
rect 10333 17493 10367 17527
rect 10367 17493 10376 17527
rect 10324 17484 10376 17493
rect 15292 17484 15344 17536
rect 15844 17484 15896 17536
rect 16488 17484 16540 17536
rect 20812 17484 20864 17536
rect 24584 17484 24636 17536
rect 26148 17484 26200 17536
rect 28448 17484 28500 17536
rect 29828 17561 29837 17595
rect 29837 17561 29871 17595
rect 29871 17561 29880 17595
rect 29828 17552 29880 17561
rect 29920 17595 29972 17604
rect 29920 17561 29929 17595
rect 29929 17561 29963 17595
rect 29963 17561 29972 17595
rect 29920 17552 29972 17561
rect 30380 17552 30432 17604
rect 30196 17527 30248 17536
rect 30196 17493 30205 17527
rect 30205 17493 30239 17527
rect 30239 17493 30248 17527
rect 32588 17688 32640 17740
rect 33140 17620 33192 17672
rect 37280 17756 37332 17808
rect 36912 17688 36964 17740
rect 37832 17731 37884 17740
rect 37832 17697 37841 17731
rect 37841 17697 37875 17731
rect 37875 17697 37884 17731
rect 37832 17688 37884 17697
rect 38936 17688 38988 17740
rect 33876 17620 33928 17672
rect 34796 17620 34848 17672
rect 36728 17663 36780 17672
rect 36728 17629 36737 17663
rect 36737 17629 36771 17663
rect 36771 17629 36780 17663
rect 36728 17620 36780 17629
rect 37004 17620 37056 17672
rect 38016 17663 38068 17672
rect 38016 17629 38025 17663
rect 38025 17629 38059 17663
rect 38059 17629 38068 17663
rect 38016 17620 38068 17629
rect 38200 17620 38252 17672
rect 38568 17620 38620 17672
rect 43076 17824 43128 17876
rect 43904 17867 43956 17876
rect 43904 17833 43913 17867
rect 43913 17833 43947 17867
rect 43947 17833 43956 17867
rect 43904 17824 43956 17833
rect 47032 17867 47084 17876
rect 47032 17833 47041 17867
rect 47041 17833 47075 17867
rect 47075 17833 47084 17867
rect 47032 17824 47084 17833
rect 47492 17824 47544 17876
rect 42800 17756 42852 17808
rect 42616 17663 42668 17672
rect 42616 17629 42625 17663
rect 42625 17629 42659 17663
rect 42659 17629 42668 17663
rect 42616 17620 42668 17629
rect 32404 17552 32456 17604
rect 33508 17595 33560 17604
rect 33508 17561 33517 17595
rect 33517 17561 33551 17595
rect 33551 17561 33560 17595
rect 33508 17552 33560 17561
rect 34336 17552 34388 17604
rect 38292 17552 38344 17604
rect 30196 17484 30248 17493
rect 32128 17484 32180 17536
rect 36268 17484 36320 17536
rect 37188 17484 37240 17536
rect 37556 17484 37608 17536
rect 44456 17688 44508 17740
rect 43168 17620 43220 17672
rect 44088 17663 44140 17672
rect 44088 17629 44097 17663
rect 44097 17629 44131 17663
rect 44131 17629 44140 17663
rect 44364 17663 44416 17672
rect 44088 17620 44140 17629
rect 44364 17629 44373 17663
rect 44373 17629 44407 17663
rect 44407 17629 44416 17663
rect 44364 17620 44416 17629
rect 46664 17620 46716 17672
rect 47860 17663 47912 17672
rect 47860 17629 47869 17663
rect 47869 17629 47903 17663
rect 47903 17629 47912 17663
rect 47860 17620 47912 17629
rect 46940 17552 46992 17604
rect 42156 17527 42208 17536
rect 42156 17493 42165 17527
rect 42165 17493 42199 17527
rect 42199 17493 42208 17527
rect 42156 17484 42208 17493
rect 42524 17484 42576 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 3884 17280 3936 17332
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 7840 17323 7892 17332
rect 2780 17212 2832 17264
rect 7840 17289 7849 17323
rect 7849 17289 7883 17323
rect 7883 17289 7892 17323
rect 7840 17280 7892 17289
rect 16488 17280 16540 17332
rect 16672 17323 16724 17332
rect 16672 17289 16681 17323
rect 16681 17289 16715 17323
rect 16715 17289 16724 17323
rect 16672 17280 16724 17289
rect 1860 17187 1912 17196
rect 1860 17153 1869 17187
rect 1869 17153 1903 17187
rect 1903 17153 1912 17187
rect 1860 17144 1912 17153
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 3976 17187 4028 17196
rect 3976 17153 3985 17187
rect 3985 17153 4019 17187
rect 4019 17153 4028 17187
rect 3976 17144 4028 17153
rect 7656 17212 7708 17264
rect 10324 17212 10376 17264
rect 12808 17255 12860 17264
rect 12808 17221 12817 17255
rect 12817 17221 12851 17255
rect 12851 17221 12860 17255
rect 12808 17212 12860 17221
rect 14372 17212 14424 17264
rect 16120 17212 16172 17264
rect 5816 17144 5868 17196
rect 6736 17144 6788 17196
rect 17868 17212 17920 17264
rect 17132 17187 17184 17196
rect 17132 17153 17141 17187
rect 17141 17153 17175 17187
rect 17175 17153 17184 17187
rect 17132 17144 17184 17153
rect 17684 17144 17736 17196
rect 14280 17076 14332 17128
rect 14832 17076 14884 17128
rect 15016 17119 15068 17128
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 15936 17076 15988 17128
rect 17592 17076 17644 17128
rect 17868 17119 17920 17128
rect 17868 17085 17877 17119
rect 17877 17085 17911 17119
rect 17911 17085 17920 17119
rect 17868 17076 17920 17085
rect 18328 17280 18380 17332
rect 18788 17280 18840 17332
rect 31944 17280 31996 17332
rect 20628 17212 20680 17264
rect 23204 17212 23256 17264
rect 25412 17212 25464 17264
rect 18236 17144 18288 17196
rect 18972 17187 19024 17196
rect 18972 17153 18981 17187
rect 18981 17153 19015 17187
rect 19015 17153 19024 17187
rect 18972 17144 19024 17153
rect 18144 17119 18196 17128
rect 18144 17085 18153 17119
rect 18153 17085 18187 17119
rect 18187 17085 18196 17119
rect 18144 17076 18196 17085
rect 18604 17076 18656 17128
rect 18696 17076 18748 17128
rect 19156 17119 19208 17128
rect 19156 17085 19165 17119
rect 19165 17085 19199 17119
rect 19199 17085 19208 17119
rect 19156 17076 19208 17085
rect 20536 17144 20588 17196
rect 23020 17144 23072 17196
rect 26148 17187 26200 17196
rect 26148 17153 26157 17187
rect 26157 17153 26191 17187
rect 26191 17153 26200 17187
rect 26148 17144 26200 17153
rect 29092 17144 29144 17196
rect 29460 17187 29512 17196
rect 28448 17076 28500 17128
rect 29460 17153 29469 17187
rect 29469 17153 29503 17187
rect 29503 17153 29512 17187
rect 29460 17144 29512 17153
rect 29552 17187 29604 17196
rect 29552 17153 29561 17187
rect 29561 17153 29595 17187
rect 29595 17153 29604 17187
rect 29552 17144 29604 17153
rect 30012 17144 30064 17196
rect 32128 17187 32180 17196
rect 29828 17076 29880 17128
rect 30380 17076 30432 17128
rect 32128 17153 32137 17187
rect 32137 17153 32171 17187
rect 32171 17153 32180 17187
rect 32128 17144 32180 17153
rect 31484 17076 31536 17128
rect 33140 17144 33192 17196
rect 35900 17280 35952 17332
rect 36084 17280 36136 17332
rect 42524 17323 42576 17332
rect 42524 17289 42533 17323
rect 42533 17289 42567 17323
rect 42567 17289 42576 17323
rect 42524 17280 42576 17289
rect 43168 17280 43220 17332
rect 33508 17255 33560 17264
rect 33508 17221 33517 17255
rect 33517 17221 33551 17255
rect 33551 17221 33560 17255
rect 33508 17212 33560 17221
rect 34428 17212 34480 17264
rect 33876 17144 33928 17196
rect 36452 17212 36504 17264
rect 42984 17212 43036 17264
rect 44088 17255 44140 17264
rect 44088 17221 44097 17255
rect 44097 17221 44131 17255
rect 44131 17221 44140 17255
rect 44088 17212 44140 17221
rect 44456 17212 44508 17264
rect 45284 17212 45336 17264
rect 47860 17212 47912 17264
rect 36636 17144 36688 17196
rect 41696 17144 41748 17196
rect 42156 17144 42208 17196
rect 44364 17187 44416 17196
rect 44364 17153 44373 17187
rect 44373 17153 44407 17187
rect 44407 17153 44416 17187
rect 44364 17144 44416 17153
rect 51448 17187 51500 17196
rect 51448 17153 51457 17187
rect 51457 17153 51491 17187
rect 51491 17153 51500 17187
rect 51448 17144 51500 17153
rect 34612 17076 34664 17128
rect 7564 16940 7616 16992
rect 10692 16940 10744 16992
rect 16856 16940 16908 16992
rect 19984 17008 20036 17060
rect 25780 16940 25832 16992
rect 25964 16983 26016 16992
rect 25964 16949 25973 16983
rect 25973 16949 26007 16983
rect 26007 16949 26016 16983
rect 25964 16940 26016 16949
rect 27252 16940 27304 16992
rect 32312 16983 32364 16992
rect 32312 16949 32321 16983
rect 32321 16949 32355 16983
rect 32355 16949 32364 16983
rect 32312 16940 32364 16949
rect 33140 16940 33192 16992
rect 36544 16983 36596 16992
rect 36544 16949 36553 16983
rect 36553 16949 36587 16983
rect 36587 16949 36596 16983
rect 36544 16940 36596 16949
rect 37096 16940 37148 16992
rect 51080 16940 51132 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 7564 16736 7616 16788
rect 3976 16668 4028 16720
rect 9956 16668 10008 16720
rect 14280 16736 14332 16788
rect 16672 16736 16724 16788
rect 1492 16600 1544 16652
rect 11428 16600 11480 16652
rect 12164 16643 12216 16652
rect 12164 16609 12173 16643
rect 12173 16609 12207 16643
rect 12207 16609 12216 16643
rect 12164 16600 12216 16609
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 16856 16643 16908 16652
rect 16856 16609 16865 16643
rect 16865 16609 16899 16643
rect 16899 16609 16908 16643
rect 16856 16600 16908 16609
rect 22744 16736 22796 16788
rect 24400 16736 24452 16788
rect 24492 16736 24544 16788
rect 25688 16736 25740 16788
rect 25780 16736 25832 16788
rect 29000 16779 29052 16788
rect 27528 16668 27580 16720
rect 28448 16711 28500 16720
rect 28448 16677 28457 16711
rect 28457 16677 28491 16711
rect 28491 16677 28500 16711
rect 28448 16668 28500 16677
rect 29000 16745 29009 16779
rect 29009 16745 29043 16779
rect 29043 16745 29052 16779
rect 29000 16736 29052 16745
rect 31944 16736 31996 16788
rect 37372 16736 37424 16788
rect 38200 16736 38252 16788
rect 44088 16736 44140 16788
rect 29276 16668 29328 16720
rect 36452 16668 36504 16720
rect 17132 16643 17184 16652
rect 17132 16609 17141 16643
rect 17141 16609 17175 16643
rect 17175 16609 17184 16643
rect 17132 16600 17184 16609
rect 17500 16600 17552 16652
rect 18144 16600 18196 16652
rect 18420 16600 18472 16652
rect 20168 16600 20220 16652
rect 23020 16600 23072 16652
rect 6552 16532 6604 16584
rect 10968 16575 11020 16584
rect 10968 16541 10977 16575
rect 10977 16541 11011 16575
rect 11011 16541 11020 16575
rect 10968 16532 11020 16541
rect 17040 16575 17092 16584
rect 2320 16464 2372 16516
rect 2412 16464 2464 16516
rect 12440 16507 12492 16516
rect 12440 16473 12474 16507
rect 12474 16473 12492 16507
rect 12440 16464 12492 16473
rect 1400 16396 1452 16448
rect 2688 16396 2740 16448
rect 6828 16396 6880 16448
rect 10876 16396 10928 16448
rect 15016 16464 15068 16516
rect 15200 16507 15252 16516
rect 15200 16473 15209 16507
rect 15209 16473 15243 16507
rect 15243 16473 15252 16507
rect 15200 16464 15252 16473
rect 15384 16507 15436 16516
rect 15384 16473 15393 16507
rect 15393 16473 15427 16507
rect 15427 16473 15436 16507
rect 15384 16464 15436 16473
rect 15752 16464 15804 16516
rect 15936 16507 15988 16516
rect 15936 16473 15945 16507
rect 15945 16473 15979 16507
rect 15979 16473 15988 16507
rect 17040 16541 17049 16575
rect 17049 16541 17083 16575
rect 17083 16541 17092 16575
rect 17040 16532 17092 16541
rect 23112 16532 23164 16584
rect 15936 16464 15988 16473
rect 14372 16439 14424 16448
rect 14372 16405 14381 16439
rect 14381 16405 14415 16439
rect 14415 16405 14424 16439
rect 14372 16396 14424 16405
rect 14556 16439 14608 16448
rect 14556 16405 14565 16439
rect 14565 16405 14599 16439
rect 14599 16405 14608 16439
rect 14556 16396 14608 16405
rect 16304 16396 16356 16448
rect 16672 16439 16724 16448
rect 16672 16405 16681 16439
rect 16681 16405 16715 16439
rect 16715 16405 16724 16439
rect 16672 16396 16724 16405
rect 21824 16464 21876 16516
rect 23480 16464 23532 16516
rect 24768 16532 24820 16584
rect 28080 16532 28132 16584
rect 29000 16532 29052 16584
rect 29644 16600 29696 16652
rect 29736 16575 29788 16584
rect 29736 16541 29745 16575
rect 29745 16541 29779 16575
rect 29779 16541 29788 16575
rect 29736 16532 29788 16541
rect 35532 16600 35584 16652
rect 37556 16643 37608 16652
rect 24676 16464 24728 16516
rect 18236 16396 18288 16448
rect 20628 16396 20680 16448
rect 22192 16396 22244 16448
rect 25688 16507 25740 16516
rect 25688 16473 25697 16507
rect 25697 16473 25731 16507
rect 25731 16473 25740 16507
rect 25688 16464 25740 16473
rect 25780 16439 25832 16448
rect 25780 16405 25789 16439
rect 25789 16405 25823 16439
rect 25823 16405 25832 16439
rect 25780 16396 25832 16405
rect 28540 16464 28592 16516
rect 31300 16575 31352 16584
rect 31300 16541 31309 16575
rect 31309 16541 31343 16575
rect 31343 16541 31352 16575
rect 31484 16575 31536 16584
rect 31300 16532 31352 16541
rect 31484 16541 31498 16575
rect 31498 16541 31532 16575
rect 31532 16541 31536 16575
rect 31484 16532 31536 16541
rect 34796 16532 34848 16584
rect 36173 16575 36225 16584
rect 36173 16541 36182 16575
rect 36182 16541 36216 16575
rect 36216 16541 36225 16575
rect 36173 16532 36225 16541
rect 36268 16572 36320 16584
rect 36268 16538 36277 16572
rect 36277 16538 36311 16572
rect 36311 16538 36320 16572
rect 37556 16609 37565 16643
rect 37565 16609 37599 16643
rect 37599 16609 37608 16643
rect 37556 16600 37608 16609
rect 37096 16575 37148 16584
rect 36268 16532 36320 16538
rect 37096 16541 37105 16575
rect 37105 16541 37139 16575
rect 37139 16541 37148 16575
rect 37096 16532 37148 16541
rect 38752 16532 38804 16584
rect 31392 16507 31444 16516
rect 29460 16396 29512 16448
rect 31392 16473 31401 16507
rect 31401 16473 31435 16507
rect 31435 16473 31444 16507
rect 31392 16464 31444 16473
rect 32772 16396 32824 16448
rect 35808 16439 35860 16448
rect 35808 16405 35817 16439
rect 35817 16405 35851 16439
rect 35851 16405 35860 16439
rect 35808 16396 35860 16405
rect 37004 16396 37056 16448
rect 42892 16668 42944 16720
rect 46664 16736 46716 16788
rect 46940 16779 46992 16788
rect 46940 16745 46949 16779
rect 46949 16745 46983 16779
rect 46983 16745 46992 16779
rect 46940 16736 46992 16745
rect 42524 16643 42576 16652
rect 41696 16532 41748 16584
rect 42248 16575 42300 16584
rect 42248 16541 42257 16575
rect 42257 16541 42291 16575
rect 42291 16541 42300 16575
rect 42248 16532 42300 16541
rect 42524 16609 42533 16643
rect 42533 16609 42567 16643
rect 42567 16609 42576 16643
rect 42524 16600 42576 16609
rect 47584 16600 47636 16652
rect 53380 16736 53432 16788
rect 50804 16643 50856 16652
rect 50804 16609 50813 16643
rect 50813 16609 50847 16643
rect 50847 16609 50856 16643
rect 50804 16600 50856 16609
rect 44364 16532 44416 16584
rect 45284 16575 45336 16584
rect 45284 16541 45293 16575
rect 45293 16541 45327 16575
rect 45327 16541 45336 16575
rect 45284 16532 45336 16541
rect 45836 16575 45888 16584
rect 45836 16541 45845 16575
rect 45845 16541 45879 16575
rect 45879 16541 45888 16575
rect 45836 16532 45888 16541
rect 45928 16575 45980 16584
rect 45928 16541 45937 16575
rect 45937 16541 45971 16575
rect 45971 16541 45980 16575
rect 45928 16532 45980 16541
rect 51080 16575 51132 16584
rect 51080 16541 51114 16575
rect 51114 16541 51132 16575
rect 51080 16532 51132 16541
rect 42892 16464 42944 16516
rect 45008 16507 45060 16516
rect 45008 16473 45017 16507
rect 45017 16473 45051 16507
rect 45051 16473 45060 16507
rect 45008 16464 45060 16473
rect 47676 16464 47728 16516
rect 53196 16464 53248 16516
rect 42524 16396 42576 16448
rect 46756 16396 46808 16448
rect 47860 16396 47912 16448
rect 49240 16439 49292 16448
rect 49240 16405 49249 16439
rect 49249 16405 49283 16439
rect 49283 16405 49292 16439
rect 49240 16396 49292 16405
rect 52460 16396 52512 16448
rect 53840 16396 53892 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 2320 16235 2372 16244
rect 2320 16201 2329 16235
rect 2329 16201 2363 16235
rect 2363 16201 2372 16235
rect 2320 16192 2372 16201
rect 2688 16235 2740 16244
rect 2688 16201 2697 16235
rect 2697 16201 2731 16235
rect 2731 16201 2740 16235
rect 2688 16192 2740 16201
rect 12440 16192 12492 16244
rect 17960 16235 18012 16244
rect 17960 16201 17969 16235
rect 17969 16201 18003 16235
rect 18003 16201 18012 16235
rect 17960 16192 18012 16201
rect 21824 16235 21876 16244
rect 21824 16201 21833 16235
rect 21833 16201 21867 16235
rect 21867 16201 21876 16235
rect 21824 16192 21876 16201
rect 22192 16235 22244 16244
rect 22192 16201 22201 16235
rect 22201 16201 22235 16235
rect 22235 16201 22244 16235
rect 22192 16192 22244 16201
rect 28172 16235 28224 16244
rect 28172 16201 28181 16235
rect 28181 16201 28215 16235
rect 28215 16201 28224 16235
rect 28172 16192 28224 16201
rect 2412 16124 2464 16176
rect 2596 16124 2648 16176
rect 14464 16124 14516 16176
rect 14556 16124 14608 16176
rect 25688 16124 25740 16176
rect 1492 16099 1544 16108
rect 1492 16065 1501 16099
rect 1501 16065 1535 16099
rect 1535 16065 1544 16099
rect 1492 16056 1544 16065
rect 2504 16099 2556 16108
rect 2504 16065 2513 16099
rect 2513 16065 2547 16099
rect 2547 16065 2556 16099
rect 2504 16056 2556 16065
rect 2780 16099 2832 16108
rect 2780 16065 2789 16099
rect 2789 16065 2823 16099
rect 2823 16065 2832 16099
rect 2780 16056 2832 16065
rect 4620 16056 4672 16108
rect 6828 16056 6880 16108
rect 8944 16056 8996 16108
rect 9496 16056 9548 16108
rect 10600 16056 10652 16108
rect 10968 16056 11020 16108
rect 11888 16056 11940 16108
rect 12532 16099 12584 16108
rect 12532 16065 12541 16099
rect 12541 16065 12575 16099
rect 12575 16065 12584 16099
rect 12532 16056 12584 16065
rect 16396 16056 16448 16108
rect 17868 16056 17920 16108
rect 18236 16099 18288 16108
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 18236 16056 18288 16065
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 22192 16056 22244 16108
rect 22376 16056 22428 16108
rect 23020 16056 23072 16108
rect 23204 16099 23256 16108
rect 23204 16065 23213 16099
rect 23213 16065 23247 16099
rect 23247 16065 23256 16099
rect 23204 16056 23256 16065
rect 24400 16056 24452 16108
rect 29000 16192 29052 16244
rect 36728 16235 36780 16244
rect 36728 16201 36737 16235
rect 36737 16201 36771 16235
rect 36771 16201 36780 16235
rect 36728 16192 36780 16201
rect 42616 16192 42668 16244
rect 46756 16235 46808 16244
rect 46756 16201 46765 16235
rect 46765 16201 46799 16235
rect 46799 16201 46808 16235
rect 46756 16192 46808 16201
rect 47676 16235 47728 16244
rect 47676 16201 47685 16235
rect 47685 16201 47719 16235
rect 47719 16201 47728 16235
rect 47676 16192 47728 16201
rect 51448 16192 51500 16244
rect 28448 16124 28500 16176
rect 28540 16099 28592 16108
rect 28540 16065 28549 16099
rect 28549 16065 28583 16099
rect 28583 16065 28592 16099
rect 28540 16056 28592 16065
rect 30288 16124 30340 16176
rect 29092 16056 29144 16108
rect 29644 16099 29696 16108
rect 29644 16065 29653 16099
rect 29653 16065 29687 16099
rect 29687 16065 29696 16099
rect 29644 16056 29696 16065
rect 29828 16099 29880 16108
rect 29828 16065 29835 16099
rect 29835 16065 29880 16099
rect 29828 16056 29880 16065
rect 3792 15988 3844 16040
rect 4712 15852 4764 15904
rect 16580 15988 16632 16040
rect 6920 15852 6972 15904
rect 8116 15895 8168 15904
rect 8116 15861 8125 15895
rect 8125 15861 8159 15895
rect 8159 15861 8168 15895
rect 8116 15852 8168 15861
rect 10968 15895 11020 15904
rect 10968 15861 10977 15895
rect 10977 15861 11011 15895
rect 11011 15861 11020 15895
rect 10968 15852 11020 15861
rect 11060 15852 11112 15904
rect 16028 15895 16080 15904
rect 16028 15861 16037 15895
rect 16037 15861 16071 15895
rect 16071 15861 16080 15895
rect 16028 15852 16080 15861
rect 28172 15988 28224 16040
rect 28724 15988 28776 16040
rect 30104 16099 30156 16108
rect 32956 16124 33008 16176
rect 30104 16065 30118 16099
rect 30118 16065 30152 16099
rect 30152 16065 30156 16099
rect 30104 16056 30156 16065
rect 32864 16099 32916 16108
rect 32864 16065 32898 16099
rect 32898 16065 32916 16099
rect 35808 16124 35860 16176
rect 45836 16124 45888 16176
rect 49240 16124 49292 16176
rect 51080 16124 51132 16176
rect 52920 16124 52972 16176
rect 32864 16056 32916 16065
rect 37556 16056 37608 16108
rect 40316 16099 40368 16108
rect 40316 16065 40325 16099
rect 40325 16065 40359 16099
rect 40359 16065 40368 16099
rect 40316 16056 40368 16065
rect 40408 16099 40460 16108
rect 40408 16065 40417 16099
rect 40417 16065 40451 16099
rect 40451 16065 40460 16099
rect 43628 16099 43680 16108
rect 40408 16056 40460 16065
rect 43628 16065 43637 16099
rect 43637 16065 43671 16099
rect 43671 16065 43680 16099
rect 43628 16056 43680 16065
rect 45008 16056 45060 16108
rect 45928 16056 45980 16108
rect 47860 16099 47912 16108
rect 47860 16065 47869 16099
rect 47869 16065 47903 16099
rect 47903 16065 47912 16099
rect 47860 16056 47912 16065
rect 53288 16056 53340 16108
rect 31300 15988 31352 16040
rect 53472 16099 53524 16108
rect 53472 16065 53481 16099
rect 53481 16065 53515 16099
rect 53515 16065 53524 16099
rect 53472 16056 53524 16065
rect 55588 15988 55640 16040
rect 53196 15963 53248 15972
rect 53196 15929 53205 15963
rect 53205 15929 53239 15963
rect 53239 15929 53248 15963
rect 53196 15920 53248 15929
rect 24768 15852 24820 15904
rect 25780 15852 25832 15904
rect 25964 15852 26016 15904
rect 27528 15852 27580 15904
rect 32772 15852 32824 15904
rect 43720 15895 43772 15904
rect 43720 15861 43729 15895
rect 43729 15861 43763 15895
rect 43763 15861 43772 15895
rect 43720 15852 43772 15861
rect 51540 15895 51592 15904
rect 51540 15861 51549 15895
rect 51549 15861 51583 15895
rect 51583 15861 51592 15895
rect 51540 15852 51592 15861
rect 52552 15852 52604 15904
rect 53472 15852 53524 15904
rect 55404 15852 55456 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2228 15648 2280 15700
rect 23756 15691 23808 15700
rect 23756 15657 23765 15691
rect 23765 15657 23799 15691
rect 23799 15657 23808 15691
rect 23756 15648 23808 15657
rect 24400 15691 24452 15700
rect 24400 15657 24409 15691
rect 24409 15657 24443 15691
rect 24443 15657 24452 15691
rect 24400 15648 24452 15657
rect 24492 15648 24544 15700
rect 6552 15623 6604 15632
rect 6552 15589 6561 15623
rect 6561 15589 6595 15623
rect 6595 15589 6604 15623
rect 6552 15580 6604 15589
rect 10600 15623 10652 15632
rect 10600 15589 10609 15623
rect 10609 15589 10643 15623
rect 10643 15589 10652 15623
rect 10600 15580 10652 15589
rect 11888 15623 11940 15632
rect 11888 15589 11897 15623
rect 11897 15589 11931 15623
rect 11931 15589 11940 15623
rect 11888 15580 11940 15589
rect 14464 15580 14516 15632
rect 5908 15512 5960 15564
rect 6736 15512 6788 15564
rect 17040 15512 17092 15564
rect 17224 15512 17276 15564
rect 17776 15580 17828 15632
rect 1952 15444 2004 15496
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 3792 15444 3844 15496
rect 4712 15444 4764 15496
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 10876 15487 10928 15496
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 11060 15487 11112 15496
rect 10876 15444 10928 15453
rect 11060 15453 11069 15487
rect 11069 15453 11103 15487
rect 11103 15453 11112 15487
rect 11060 15444 11112 15453
rect 11152 15487 11204 15496
rect 11152 15453 11161 15487
rect 11161 15453 11195 15487
rect 11195 15453 11204 15487
rect 11152 15444 11204 15453
rect 11612 15376 11664 15428
rect 13268 15444 13320 15496
rect 15752 15444 15804 15496
rect 17592 15487 17644 15496
rect 17592 15453 17601 15487
rect 17601 15453 17635 15487
rect 17635 15453 17644 15487
rect 17592 15444 17644 15453
rect 17776 15487 17828 15496
rect 17776 15453 17785 15487
rect 17785 15453 17819 15487
rect 17819 15453 17828 15487
rect 17776 15444 17828 15453
rect 5448 15351 5500 15360
rect 5448 15317 5457 15351
rect 5457 15317 5491 15351
rect 5491 15317 5500 15351
rect 5448 15308 5500 15317
rect 8116 15308 8168 15360
rect 10324 15308 10376 15360
rect 17132 15376 17184 15428
rect 19432 15444 19484 15496
rect 20168 15487 20220 15496
rect 20168 15453 20177 15487
rect 20177 15453 20211 15487
rect 20211 15453 20220 15487
rect 20168 15444 20220 15453
rect 23020 15512 23072 15564
rect 24492 15444 24544 15496
rect 24676 15444 24728 15496
rect 24952 15444 25004 15496
rect 21824 15376 21876 15428
rect 23388 15419 23440 15428
rect 23388 15385 23397 15419
rect 23397 15385 23431 15419
rect 23431 15385 23440 15419
rect 23388 15376 23440 15385
rect 25412 15512 25464 15564
rect 25964 15376 26016 15428
rect 26240 15419 26292 15428
rect 26240 15385 26274 15419
rect 26274 15385 26292 15419
rect 26240 15376 26292 15385
rect 15200 15308 15252 15360
rect 21548 15351 21600 15360
rect 21548 15317 21557 15351
rect 21557 15317 21591 15351
rect 21591 15317 21600 15351
rect 21548 15308 21600 15317
rect 24768 15351 24820 15360
rect 24768 15317 24777 15351
rect 24777 15317 24811 15351
rect 24811 15317 24820 15351
rect 24768 15308 24820 15317
rect 24860 15308 24912 15360
rect 27160 15308 27212 15360
rect 29276 15444 29328 15496
rect 45928 15648 45980 15700
rect 51540 15648 51592 15700
rect 52920 15691 52972 15700
rect 52920 15657 52929 15691
rect 52929 15657 52963 15691
rect 52963 15657 52972 15691
rect 52920 15648 52972 15657
rect 41512 15580 41564 15632
rect 30932 15512 30984 15564
rect 42524 15555 42576 15564
rect 42524 15521 42533 15555
rect 42533 15521 42567 15555
rect 42567 15521 42576 15555
rect 42524 15512 42576 15521
rect 43628 15512 43680 15564
rect 32772 15487 32824 15496
rect 29092 15376 29144 15428
rect 29828 15376 29880 15428
rect 30196 15376 30248 15428
rect 32772 15453 32781 15487
rect 32781 15453 32815 15487
rect 32815 15453 32824 15487
rect 32772 15444 32824 15453
rect 43536 15444 43588 15496
rect 43720 15487 43772 15496
rect 43720 15453 43729 15487
rect 43729 15453 43763 15487
rect 43763 15453 43772 15487
rect 43720 15444 43772 15453
rect 52460 15580 52512 15632
rect 53104 15580 53156 15632
rect 53380 15580 53432 15632
rect 48044 15487 48096 15496
rect 48044 15453 48053 15487
rect 48053 15453 48087 15487
rect 48087 15453 48096 15487
rect 48044 15444 48096 15453
rect 52552 15512 52604 15564
rect 54024 15512 54076 15564
rect 52460 15487 52512 15496
rect 52460 15453 52469 15487
rect 52469 15453 52503 15487
rect 52503 15453 52512 15487
rect 52460 15444 52512 15453
rect 53288 15487 53340 15496
rect 40408 15376 40460 15428
rect 42248 15376 42300 15428
rect 44088 15419 44140 15428
rect 44088 15385 44097 15419
rect 44097 15385 44131 15419
rect 44131 15385 44140 15419
rect 44088 15376 44140 15385
rect 53288 15453 53297 15487
rect 53297 15453 53331 15487
rect 53331 15453 53340 15487
rect 53288 15444 53340 15453
rect 53380 15487 53432 15496
rect 53380 15453 53389 15487
rect 53389 15453 53423 15487
rect 53423 15453 53432 15487
rect 53380 15444 53432 15453
rect 53840 15444 53892 15496
rect 55680 15487 55732 15496
rect 55680 15453 55689 15487
rect 55689 15453 55723 15487
rect 55723 15453 55732 15487
rect 55680 15444 55732 15453
rect 29000 15308 29052 15360
rect 30012 15308 30064 15360
rect 33508 15308 33560 15360
rect 42892 15351 42944 15360
rect 42892 15317 42901 15351
rect 42901 15317 42935 15351
rect 42935 15317 42944 15351
rect 47860 15351 47912 15360
rect 42892 15308 42944 15317
rect 47860 15317 47869 15351
rect 47869 15317 47903 15351
rect 47903 15317 47912 15351
rect 47860 15308 47912 15317
rect 55220 15376 55272 15428
rect 55404 15376 55456 15428
rect 53288 15308 53340 15360
rect 55772 15351 55824 15360
rect 55772 15317 55781 15351
rect 55781 15317 55815 15351
rect 55815 15317 55824 15351
rect 55772 15308 55824 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4620 15104 4672 15156
rect 7012 15104 7064 15156
rect 2504 15036 2556 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 2780 14968 2832 15020
rect 5448 14968 5500 15020
rect 5908 14900 5960 14952
rect 6184 15036 6236 15088
rect 7472 14968 7524 15020
rect 12532 15104 12584 15156
rect 11612 15036 11664 15088
rect 16120 15104 16172 15156
rect 16396 15036 16448 15088
rect 17132 15036 17184 15088
rect 17592 15104 17644 15156
rect 21824 15147 21876 15156
rect 21824 15113 21833 15147
rect 21833 15113 21867 15147
rect 21867 15113 21876 15147
rect 21824 15104 21876 15113
rect 23480 15147 23532 15156
rect 23480 15113 23489 15147
rect 23489 15113 23523 15147
rect 23523 15113 23532 15147
rect 23480 15104 23532 15113
rect 23940 15147 23992 15156
rect 23940 15113 23949 15147
rect 23949 15113 23983 15147
rect 23983 15113 23992 15147
rect 23940 15104 23992 15113
rect 24676 15147 24728 15156
rect 24676 15113 24685 15147
rect 24685 15113 24719 15147
rect 24719 15113 24728 15147
rect 24676 15104 24728 15113
rect 26240 15104 26292 15156
rect 29276 15104 29328 15156
rect 30012 15104 30064 15156
rect 30932 15147 30984 15156
rect 17960 15036 18012 15088
rect 14096 14968 14148 15020
rect 17500 14968 17552 15020
rect 17868 14968 17920 15020
rect 23020 15079 23072 15088
rect 21548 14968 21600 15020
rect 23020 15045 23029 15079
rect 23029 15045 23063 15079
rect 23063 15045 23072 15079
rect 23020 15036 23072 15045
rect 24308 15079 24360 15088
rect 24308 15045 24317 15079
rect 24317 15045 24351 15079
rect 24351 15045 24360 15079
rect 24308 15036 24360 15045
rect 22836 15011 22888 15020
rect 8024 14900 8076 14952
rect 12072 14943 12124 14952
rect 12072 14909 12081 14943
rect 12081 14909 12115 14943
rect 12115 14909 12124 14943
rect 12072 14900 12124 14909
rect 13268 14943 13320 14952
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 17040 14943 17092 14952
rect 13268 14900 13320 14909
rect 17040 14909 17049 14943
rect 17049 14909 17083 14943
rect 17083 14909 17092 14943
rect 17040 14900 17092 14909
rect 7288 14764 7340 14816
rect 7472 14764 7524 14816
rect 8484 14832 8536 14884
rect 11888 14832 11940 14884
rect 12072 14764 12124 14816
rect 16672 14764 16724 14816
rect 17224 14943 17276 14952
rect 17224 14909 17233 14943
rect 17233 14909 17267 14943
rect 17267 14909 17276 14943
rect 17224 14900 17276 14909
rect 17776 14900 17828 14952
rect 22836 14977 22845 15011
rect 22845 14977 22879 15011
rect 22879 14977 22888 15011
rect 22836 14968 22888 14977
rect 23388 14968 23440 15020
rect 24032 14968 24084 15020
rect 26424 15036 26476 15088
rect 29828 15036 29880 15088
rect 23848 14900 23900 14952
rect 24952 14832 25004 14884
rect 23940 14764 23992 14816
rect 24492 14807 24544 14816
rect 24492 14773 24501 14807
rect 24501 14773 24535 14807
rect 24535 14773 24544 14807
rect 24492 14764 24544 14773
rect 27160 15011 27212 15020
rect 27160 14977 27169 15011
rect 27169 14977 27203 15011
rect 27203 14977 27212 15011
rect 27160 14968 27212 14977
rect 29092 14968 29144 15020
rect 29276 15011 29328 15020
rect 29276 14977 29285 15011
rect 29285 14977 29319 15011
rect 29319 14977 29328 15011
rect 29276 14968 29328 14977
rect 30472 14968 30524 15020
rect 26056 14943 26108 14952
rect 26056 14909 26065 14943
rect 26065 14909 26099 14943
rect 26099 14909 26108 14943
rect 26056 14900 26108 14909
rect 26424 14900 26476 14952
rect 26884 14900 26936 14952
rect 30380 14900 30432 14952
rect 30932 15113 30941 15147
rect 30941 15113 30975 15147
rect 30975 15113 30984 15147
rect 30932 15104 30984 15113
rect 32864 15147 32916 15156
rect 32864 15113 32873 15147
rect 32873 15113 32907 15147
rect 32907 15113 32916 15147
rect 32864 15104 32916 15113
rect 38936 15104 38988 15156
rect 41512 15104 41564 15156
rect 42892 15104 42944 15156
rect 45008 15147 45060 15156
rect 45008 15113 45017 15147
rect 45017 15113 45051 15147
rect 45051 15113 45060 15147
rect 45008 15104 45060 15113
rect 33508 15079 33560 15088
rect 33508 15045 33517 15079
rect 33517 15045 33551 15079
rect 33551 15045 33560 15079
rect 33508 15036 33560 15045
rect 37832 15036 37884 15088
rect 30932 15011 30984 15020
rect 30932 14977 30941 15011
rect 30941 14977 30975 15011
rect 30975 14977 30984 15011
rect 33140 15011 33192 15020
rect 30932 14968 30984 14977
rect 33140 14977 33149 15011
rect 33149 14977 33183 15011
rect 33183 14977 33192 15011
rect 33140 14968 33192 14977
rect 33324 14968 33376 15020
rect 38844 14968 38896 15020
rect 40316 14968 40368 15020
rect 41052 15036 41104 15088
rect 42800 15036 42852 15088
rect 43168 15036 43220 15088
rect 44088 15036 44140 15088
rect 41604 15011 41656 15020
rect 38936 14900 38988 14952
rect 41604 14977 41613 15011
rect 41613 14977 41647 15011
rect 41647 14977 41656 15011
rect 41604 14968 41656 14977
rect 53564 15104 53616 15156
rect 55036 15104 55088 15156
rect 47860 15079 47912 15088
rect 47860 15045 47894 15079
rect 47894 15045 47912 15079
rect 47860 15036 47912 15045
rect 55404 15079 55456 15088
rect 41052 14900 41104 14952
rect 33416 14832 33468 14884
rect 36452 14832 36504 14884
rect 42524 14900 42576 14952
rect 43076 14900 43128 14952
rect 46020 14900 46072 14952
rect 28540 14764 28592 14816
rect 29828 14764 29880 14816
rect 38476 14807 38528 14816
rect 38476 14773 38485 14807
rect 38485 14773 38519 14807
rect 38519 14773 38528 14807
rect 38476 14764 38528 14773
rect 38660 14764 38712 14816
rect 49056 14832 49108 14884
rect 48964 14807 49016 14816
rect 48964 14773 48973 14807
rect 48973 14773 49007 14807
rect 49007 14773 49016 14807
rect 48964 14764 49016 14773
rect 55404 15045 55413 15079
rect 55413 15045 55447 15079
rect 55447 15045 55456 15079
rect 55404 15036 55456 15045
rect 55772 15036 55824 15088
rect 52552 14968 52604 15020
rect 53288 14968 53340 15020
rect 55220 15011 55272 15020
rect 55220 14977 55229 15011
rect 55229 14977 55263 15011
rect 55263 14977 55272 15011
rect 55220 14968 55272 14977
rect 53104 14943 53156 14952
rect 53104 14909 53113 14943
rect 53113 14909 53147 14943
rect 53147 14909 53156 14943
rect 53104 14900 53156 14909
rect 53196 14943 53248 14952
rect 53196 14909 53205 14943
rect 53205 14909 53239 14943
rect 53239 14909 53248 14943
rect 53196 14900 53248 14909
rect 54024 14900 54076 14952
rect 55036 14943 55088 14952
rect 55036 14909 55045 14943
rect 55045 14909 55079 14943
rect 55079 14909 55088 14943
rect 55036 14900 55088 14909
rect 50620 14764 50672 14816
rect 50896 14807 50948 14816
rect 50896 14773 50905 14807
rect 50905 14773 50939 14807
rect 50939 14773 50948 14807
rect 50896 14764 50948 14773
rect 56324 14764 56376 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1952 14560 2004 14612
rect 2688 14560 2740 14612
rect 5448 14560 5500 14612
rect 7840 14560 7892 14612
rect 8116 14560 8168 14612
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 16028 14560 16080 14612
rect 17040 14560 17092 14612
rect 17592 14560 17644 14612
rect 17960 14560 18012 14612
rect 2596 14356 2648 14408
rect 2320 14288 2372 14340
rect 14556 14492 14608 14544
rect 23388 14560 23440 14612
rect 26056 14560 26108 14612
rect 29276 14560 29328 14612
rect 30196 14560 30248 14612
rect 36636 14560 36688 14612
rect 38660 14560 38712 14612
rect 39028 14560 39080 14612
rect 7932 14467 7984 14476
rect 7932 14433 7941 14467
rect 7941 14433 7975 14467
rect 7975 14433 7984 14467
rect 7932 14424 7984 14433
rect 7012 14356 7064 14408
rect 7380 14356 7432 14408
rect 7840 14356 7892 14408
rect 10600 14424 10652 14476
rect 17592 14467 17644 14476
rect 17592 14433 17601 14467
rect 17601 14433 17635 14467
rect 17635 14433 17644 14467
rect 17592 14424 17644 14433
rect 17776 14467 17828 14476
rect 17776 14433 17785 14467
rect 17785 14433 17819 14467
rect 17819 14433 17828 14467
rect 17776 14424 17828 14433
rect 17868 14424 17920 14476
rect 24584 14492 24636 14544
rect 21180 14424 21232 14476
rect 24308 14424 24360 14476
rect 8116 14356 8168 14408
rect 1768 14220 1820 14272
rect 7196 14288 7248 14340
rect 6644 14263 6696 14272
rect 6644 14229 6653 14263
rect 6653 14229 6687 14263
rect 6687 14229 6696 14263
rect 6644 14220 6696 14229
rect 8484 14288 8536 14340
rect 13544 14356 13596 14408
rect 14556 14399 14608 14408
rect 14556 14365 14565 14399
rect 14565 14365 14599 14399
rect 14599 14365 14608 14399
rect 16488 14399 16540 14408
rect 14556 14356 14608 14365
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 17132 14356 17184 14408
rect 17500 14399 17552 14408
rect 17500 14365 17509 14399
rect 17509 14365 17543 14399
rect 17543 14365 17552 14399
rect 17500 14356 17552 14365
rect 7748 14220 7800 14272
rect 9772 14220 9824 14272
rect 9956 14220 10008 14272
rect 17224 14288 17276 14340
rect 22836 14356 22888 14408
rect 34704 14492 34756 14544
rect 35532 14535 35584 14544
rect 35532 14501 35541 14535
rect 35541 14501 35575 14535
rect 35575 14501 35584 14535
rect 35532 14492 35584 14501
rect 37740 14492 37792 14544
rect 41696 14535 41748 14544
rect 41696 14501 41705 14535
rect 41705 14501 41739 14535
rect 41739 14501 41748 14535
rect 41696 14492 41748 14501
rect 25688 14356 25740 14408
rect 26884 14356 26936 14408
rect 28172 14399 28224 14408
rect 28172 14365 28181 14399
rect 28181 14365 28215 14399
rect 28215 14365 28224 14399
rect 28172 14356 28224 14365
rect 29460 14356 29512 14408
rect 20628 14288 20680 14340
rect 24400 14288 24452 14340
rect 27160 14288 27212 14340
rect 16764 14220 16816 14272
rect 20076 14220 20128 14272
rect 37556 14424 37608 14476
rect 29828 14399 29880 14408
rect 29828 14365 29862 14399
rect 29862 14365 29880 14399
rect 29828 14356 29880 14365
rect 33324 14356 33376 14408
rect 37832 14356 37884 14408
rect 38476 14356 38528 14408
rect 36360 14288 36412 14340
rect 36544 14331 36596 14340
rect 36544 14297 36553 14331
rect 36553 14297 36587 14331
rect 36587 14297 36596 14331
rect 36544 14288 36596 14297
rect 36728 14288 36780 14340
rect 41604 14424 41656 14476
rect 48044 14560 48096 14612
rect 51080 14560 51132 14612
rect 53196 14560 53248 14612
rect 55220 14560 55272 14612
rect 55680 14560 55732 14612
rect 50804 14467 50856 14476
rect 41512 14356 41564 14408
rect 42248 14356 42300 14408
rect 42800 14288 42852 14340
rect 50804 14433 50813 14467
rect 50813 14433 50847 14467
rect 50847 14433 50856 14467
rect 50804 14424 50856 14433
rect 55588 14467 55640 14476
rect 55588 14433 55597 14467
rect 55597 14433 55631 14467
rect 55631 14433 55640 14467
rect 55588 14424 55640 14433
rect 49056 14399 49108 14408
rect 49056 14365 49065 14399
rect 49065 14365 49099 14399
rect 49099 14365 49108 14399
rect 49056 14356 49108 14365
rect 48504 14288 48556 14340
rect 48964 14288 49016 14340
rect 50896 14356 50948 14408
rect 55036 14356 55088 14408
rect 32128 14220 32180 14272
rect 32956 14220 33008 14272
rect 37740 14220 37792 14272
rect 39028 14220 39080 14272
rect 40408 14220 40460 14272
rect 41880 14263 41932 14272
rect 41880 14229 41889 14263
rect 41889 14229 41923 14263
rect 41923 14229 41932 14263
rect 41880 14220 41932 14229
rect 47860 14220 47912 14272
rect 51908 14220 51960 14272
rect 54208 14220 54260 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 2320 14059 2372 14068
rect 2320 14025 2329 14059
rect 2329 14025 2363 14059
rect 2363 14025 2372 14059
rect 2320 14016 2372 14025
rect 2688 14059 2740 14068
rect 2688 14025 2697 14059
rect 2697 14025 2731 14059
rect 2731 14025 2740 14059
rect 2688 14016 2740 14025
rect 7288 14016 7340 14068
rect 7748 13991 7800 14000
rect 2872 13880 2924 13932
rect 3976 13880 4028 13932
rect 7748 13957 7757 13991
rect 7757 13957 7791 13991
rect 7791 13957 7800 13991
rect 7748 13948 7800 13957
rect 7932 13948 7984 14000
rect 8208 13948 8260 14000
rect 9772 13991 9824 14000
rect 9772 13957 9781 13991
rect 9781 13957 9815 13991
rect 9815 13957 9824 13991
rect 9772 13948 9824 13957
rect 12072 13948 12124 14000
rect 10048 13880 10100 13932
rect 10692 13880 10744 13932
rect 14280 13991 14332 14000
rect 14280 13957 14305 13991
rect 14305 13957 14332 13991
rect 14556 14016 14608 14068
rect 16488 14016 16540 14068
rect 20628 14016 20680 14068
rect 23664 14016 23716 14068
rect 24768 14016 24820 14068
rect 25320 14016 25372 14068
rect 26424 14016 26476 14068
rect 30472 14016 30524 14068
rect 34060 14016 34112 14068
rect 36452 14059 36504 14068
rect 36452 14025 36461 14059
rect 36461 14025 36495 14059
rect 36495 14025 36504 14059
rect 36452 14016 36504 14025
rect 37832 14059 37884 14068
rect 37832 14025 37841 14059
rect 37841 14025 37875 14059
rect 37875 14025 37884 14059
rect 37832 14016 37884 14025
rect 38568 14016 38620 14068
rect 38844 14016 38896 14068
rect 41420 14016 41472 14068
rect 41880 14016 41932 14068
rect 52184 14016 52236 14068
rect 54024 14059 54076 14068
rect 54024 14025 54033 14059
rect 54033 14025 54067 14059
rect 54067 14025 54076 14059
rect 54024 14016 54076 14025
rect 54208 14059 54260 14068
rect 54208 14025 54217 14059
rect 54217 14025 54251 14059
rect 54251 14025 54260 14059
rect 54208 14016 54260 14025
rect 14280 13948 14332 13957
rect 16764 13948 16816 14000
rect 14556 13880 14608 13932
rect 22468 13948 22520 14000
rect 23480 13948 23532 14000
rect 17224 13880 17276 13932
rect 17500 13880 17552 13932
rect 18512 13880 18564 13932
rect 19432 13923 19484 13932
rect 19432 13889 19441 13923
rect 19441 13889 19475 13923
rect 19475 13889 19484 13923
rect 19432 13880 19484 13889
rect 19984 13880 20036 13932
rect 22192 13880 22244 13932
rect 4620 13812 4672 13864
rect 6644 13812 6696 13864
rect 7288 13744 7340 13796
rect 7748 13744 7800 13796
rect 8024 13787 8076 13796
rect 8024 13753 8033 13787
rect 8033 13753 8067 13787
rect 8067 13753 8076 13787
rect 8024 13744 8076 13753
rect 9956 13787 10008 13796
rect 9956 13753 9965 13787
rect 9965 13753 9999 13787
rect 9999 13753 10008 13787
rect 9956 13744 10008 13753
rect 10600 13855 10652 13864
rect 10600 13821 10609 13855
rect 10609 13821 10643 13855
rect 10643 13821 10652 13855
rect 10600 13812 10652 13821
rect 11428 13812 11480 13864
rect 12164 13812 12216 13864
rect 16672 13855 16724 13864
rect 16672 13821 16681 13855
rect 16681 13821 16715 13855
rect 16715 13821 16724 13855
rect 16672 13812 16724 13821
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17960 13855 18012 13864
rect 17132 13812 17184 13821
rect 17960 13821 17969 13855
rect 17969 13821 18003 13855
rect 18003 13821 18012 13855
rect 17960 13812 18012 13821
rect 16764 13744 16816 13796
rect 16948 13744 17000 13796
rect 17776 13744 17828 13796
rect 18052 13744 18104 13796
rect 20996 13812 21048 13864
rect 23020 13812 23072 13864
rect 23848 13812 23900 13864
rect 24124 13812 24176 13864
rect 24676 13880 24728 13932
rect 31576 13948 31628 14000
rect 25688 13923 25740 13932
rect 25688 13889 25697 13923
rect 25697 13889 25731 13923
rect 25731 13889 25740 13923
rect 25688 13880 25740 13889
rect 32956 13880 33008 13932
rect 33324 13880 33376 13932
rect 36360 13948 36412 14000
rect 38384 13948 38436 14000
rect 38476 13948 38528 14000
rect 25688 13744 25740 13796
rect 34612 13787 34664 13796
rect 34612 13753 34621 13787
rect 34621 13753 34655 13787
rect 34655 13753 34664 13787
rect 34612 13744 34664 13753
rect 38568 13923 38620 13932
rect 38568 13889 38577 13923
rect 38577 13889 38611 13923
rect 38611 13889 38620 13923
rect 38568 13880 38620 13889
rect 38752 13923 38804 13932
rect 38752 13889 38761 13923
rect 38761 13889 38795 13923
rect 38795 13889 38804 13923
rect 40408 13923 40460 13932
rect 38752 13880 38804 13889
rect 40408 13889 40417 13923
rect 40417 13889 40451 13923
rect 40451 13889 40460 13923
rect 40408 13880 40460 13889
rect 41696 13880 41748 13932
rect 53196 13948 53248 14000
rect 53840 13991 53892 14000
rect 53840 13957 53849 13991
rect 53849 13957 53883 13991
rect 53883 13957 53892 13991
rect 53840 13948 53892 13957
rect 36176 13812 36228 13864
rect 36728 13812 36780 13864
rect 36912 13812 36964 13864
rect 40316 13812 40368 13864
rect 40776 13812 40828 13864
rect 42524 13812 42576 13864
rect 36636 13744 36688 13796
rect 47400 13880 47452 13932
rect 54116 13923 54168 13932
rect 47860 13855 47912 13864
rect 47860 13821 47869 13855
rect 47869 13821 47903 13855
rect 47903 13821 47912 13855
rect 47860 13812 47912 13821
rect 53104 13812 53156 13864
rect 54116 13889 54125 13923
rect 54125 13889 54159 13923
rect 54159 13889 54168 13923
rect 54116 13880 54168 13889
rect 54576 13812 54628 13864
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 6920 13676 6972 13728
rect 10140 13676 10192 13728
rect 14740 13676 14792 13728
rect 18144 13676 18196 13728
rect 19432 13676 19484 13728
rect 23664 13676 23716 13728
rect 24308 13676 24360 13728
rect 24584 13719 24636 13728
rect 24584 13685 24593 13719
rect 24593 13685 24627 13719
rect 24627 13685 24636 13719
rect 24584 13676 24636 13685
rect 25596 13676 25648 13728
rect 26240 13719 26292 13728
rect 26240 13685 26249 13719
rect 26249 13685 26283 13719
rect 26283 13685 26292 13719
rect 26240 13676 26292 13685
rect 30380 13676 30432 13728
rect 37924 13676 37976 13728
rect 42800 13676 42852 13728
rect 46204 13676 46256 13728
rect 53288 13719 53340 13728
rect 53288 13685 53297 13719
rect 53297 13685 53331 13719
rect 53331 13685 53340 13719
rect 53288 13676 53340 13685
rect 53932 13676 53984 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 6920 13515 6972 13524
rect 6920 13481 6929 13515
rect 6929 13481 6963 13515
rect 6963 13481 6972 13515
rect 6920 13472 6972 13481
rect 7104 13472 7156 13524
rect 7656 13472 7708 13524
rect 8024 13472 8076 13524
rect 10048 13472 10100 13524
rect 10232 13515 10284 13524
rect 10232 13481 10241 13515
rect 10241 13481 10275 13515
rect 10275 13481 10284 13515
rect 10232 13472 10284 13481
rect 19984 13515 20036 13524
rect 6644 13404 6696 13456
rect 7748 13404 7800 13456
rect 8116 13404 8168 13456
rect 9956 13404 10008 13456
rect 2596 13336 2648 13388
rect 3792 13379 3844 13388
rect 3792 13345 3801 13379
rect 3801 13345 3835 13379
rect 3835 13345 3844 13379
rect 3792 13336 3844 13345
rect 7196 13336 7248 13388
rect 10600 13404 10652 13456
rect 19984 13481 19993 13515
rect 19993 13481 20027 13515
rect 20027 13481 20036 13515
rect 19984 13472 20036 13481
rect 22100 13515 22152 13524
rect 22100 13481 22109 13515
rect 22109 13481 22143 13515
rect 22143 13481 22152 13515
rect 22100 13472 22152 13481
rect 22836 13472 22888 13524
rect 23112 13515 23164 13524
rect 23112 13481 23121 13515
rect 23121 13481 23155 13515
rect 23155 13481 23164 13515
rect 23112 13472 23164 13481
rect 30380 13472 30432 13524
rect 30472 13472 30524 13524
rect 33324 13515 33376 13524
rect 33324 13481 33333 13515
rect 33333 13481 33367 13515
rect 33367 13481 33376 13515
rect 33324 13472 33376 13481
rect 36636 13472 36688 13524
rect 38016 13472 38068 13524
rect 38476 13472 38528 13524
rect 41420 13515 41472 13524
rect 41420 13481 41429 13515
rect 41429 13481 41463 13515
rect 41463 13481 41472 13515
rect 41420 13472 41472 13481
rect 42800 13515 42852 13524
rect 42800 13481 42809 13515
rect 42809 13481 42843 13515
rect 42843 13481 42852 13515
rect 42800 13472 42852 13481
rect 50620 13472 50672 13524
rect 54576 13515 54628 13524
rect 20444 13404 20496 13456
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 2780 13268 2832 13320
rect 7564 13268 7616 13320
rect 7932 13268 7984 13320
rect 8024 13268 8076 13320
rect 11428 13379 11480 13388
rect 11428 13345 11437 13379
rect 11437 13345 11471 13379
rect 11471 13345 11480 13379
rect 11428 13336 11480 13345
rect 23296 13404 23348 13456
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 11796 13268 11848 13320
rect 12256 13268 12308 13320
rect 18144 13268 18196 13320
rect 22652 13336 22704 13388
rect 34520 13404 34572 13456
rect 25044 13336 25096 13388
rect 25412 13336 25464 13388
rect 33140 13336 33192 13388
rect 21916 13311 21968 13320
rect 4068 13243 4120 13252
rect 4068 13209 4102 13243
rect 4102 13209 4120 13243
rect 4068 13200 4120 13209
rect 8392 13200 8444 13252
rect 9772 13200 9824 13252
rect 10416 13200 10468 13252
rect 10692 13200 10744 13252
rect 14188 13200 14240 13252
rect 19432 13200 19484 13252
rect 21916 13277 21925 13311
rect 21925 13277 21959 13311
rect 21959 13277 21968 13311
rect 21916 13268 21968 13277
rect 22836 13268 22888 13320
rect 24768 13268 24820 13320
rect 25688 13268 25740 13320
rect 27896 13268 27948 13320
rect 28448 13311 28500 13320
rect 28448 13277 28457 13311
rect 28457 13277 28491 13311
rect 28491 13277 28500 13311
rect 28448 13268 28500 13277
rect 30380 13311 30432 13320
rect 30380 13277 30389 13311
rect 30389 13277 30423 13311
rect 30423 13277 30432 13311
rect 31852 13311 31904 13320
rect 30380 13268 30432 13277
rect 22100 13200 22152 13252
rect 23480 13200 23532 13252
rect 26240 13200 26292 13252
rect 31852 13277 31861 13311
rect 31861 13277 31895 13311
rect 31895 13277 31904 13311
rect 31852 13268 31904 13277
rect 33324 13268 33376 13320
rect 34060 13336 34112 13388
rect 46020 13379 46072 13388
rect 46020 13345 46029 13379
rect 46029 13345 46063 13379
rect 46063 13345 46072 13379
rect 46020 13336 46072 13345
rect 36544 13268 36596 13320
rect 38660 13268 38712 13320
rect 39028 13311 39080 13320
rect 39028 13277 39037 13311
rect 39037 13277 39071 13311
rect 39071 13277 39080 13311
rect 39028 13268 39080 13277
rect 40408 13268 40460 13320
rect 42432 13311 42484 13320
rect 42432 13277 42441 13311
rect 42441 13277 42475 13311
rect 42475 13277 42484 13311
rect 42432 13268 42484 13277
rect 42892 13268 42944 13320
rect 48504 13311 48556 13320
rect 48504 13277 48513 13311
rect 48513 13277 48547 13311
rect 48547 13277 48556 13311
rect 48504 13268 48556 13277
rect 51264 13268 51316 13320
rect 54576 13481 54585 13515
rect 54585 13481 54619 13515
rect 54619 13481 54628 13515
rect 54576 13472 54628 13481
rect 55036 13472 55088 13524
rect 54852 13404 54904 13456
rect 53288 13311 53340 13320
rect 53288 13277 53297 13311
rect 53297 13277 53331 13311
rect 53331 13277 53340 13311
rect 53288 13268 53340 13277
rect 53932 13268 53984 13320
rect 55220 13336 55272 13388
rect 56324 13311 56376 13320
rect 34612 13200 34664 13252
rect 41052 13243 41104 13252
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 2136 13175 2188 13184
rect 2136 13141 2145 13175
rect 2145 13141 2179 13175
rect 2179 13141 2188 13175
rect 2136 13132 2188 13141
rect 4620 13132 4672 13184
rect 7196 13132 7248 13184
rect 7564 13175 7616 13184
rect 7564 13141 7573 13175
rect 7573 13141 7607 13175
rect 7607 13141 7616 13175
rect 7564 13132 7616 13141
rect 7932 13132 7984 13184
rect 8484 13132 8536 13184
rect 11520 13132 11572 13184
rect 14556 13132 14608 13184
rect 20628 13132 20680 13184
rect 21732 13132 21784 13184
rect 22192 13132 22244 13184
rect 24032 13132 24084 13184
rect 26608 13175 26660 13184
rect 26608 13141 26617 13175
rect 26617 13141 26651 13175
rect 26651 13141 26660 13175
rect 26608 13132 26660 13141
rect 31668 13175 31720 13184
rect 31668 13141 31677 13175
rect 31677 13141 31711 13175
rect 31711 13141 31720 13175
rect 31668 13132 31720 13141
rect 33324 13132 33376 13184
rect 41052 13209 41061 13243
rect 41061 13209 41095 13243
rect 41095 13209 41104 13243
rect 41052 13200 41104 13209
rect 46112 13200 46164 13252
rect 48688 13200 48740 13252
rect 54116 13200 54168 13252
rect 54852 13200 54904 13252
rect 56324 13277 56333 13311
rect 56333 13277 56367 13311
rect 56367 13277 56376 13311
rect 56324 13268 56376 13277
rect 56048 13200 56100 13252
rect 38568 13175 38620 13184
rect 38568 13141 38577 13175
rect 38577 13141 38611 13175
rect 38611 13141 38620 13175
rect 38568 13132 38620 13141
rect 39120 13132 39172 13184
rect 42248 13132 42300 13184
rect 47400 13175 47452 13184
rect 47400 13141 47409 13175
rect 47409 13141 47443 13175
rect 47443 13141 47452 13175
rect 47400 13132 47452 13141
rect 48596 13175 48648 13184
rect 48596 13141 48605 13175
rect 48605 13141 48639 13175
rect 48639 13141 48648 13175
rect 48596 13132 48648 13141
rect 51172 13175 51224 13184
rect 51172 13141 51181 13175
rect 51181 13141 51215 13175
rect 51215 13141 51224 13175
rect 51172 13132 51224 13141
rect 51816 13175 51868 13184
rect 51816 13141 51825 13175
rect 51825 13141 51859 13175
rect 51859 13141 51868 13175
rect 51816 13132 51868 13141
rect 52000 13132 52052 13184
rect 56232 13132 56284 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4068 12971 4120 12980
rect 4068 12937 4077 12971
rect 4077 12937 4111 12971
rect 4111 12937 4120 12971
rect 4068 12928 4120 12937
rect 4620 12928 4672 12980
rect 7104 12928 7156 12980
rect 7380 12928 7432 12980
rect 7748 12928 7800 12980
rect 10416 12928 10468 12980
rect 14188 12971 14240 12980
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 3608 12835 3660 12844
rect 3608 12801 3617 12835
rect 3617 12801 3651 12835
rect 3651 12801 3660 12835
rect 3608 12792 3660 12801
rect 2872 12631 2924 12640
rect 2872 12597 2881 12631
rect 2881 12597 2915 12631
rect 2915 12597 2924 12631
rect 2872 12588 2924 12597
rect 3424 12631 3476 12640
rect 3424 12597 3433 12631
rect 3433 12597 3467 12631
rect 3467 12597 3476 12631
rect 3424 12588 3476 12597
rect 4344 12792 4396 12844
rect 5264 12792 5316 12844
rect 6644 12792 6696 12844
rect 7380 12792 7432 12844
rect 7564 12792 7616 12844
rect 8484 12792 8536 12844
rect 10784 12860 10836 12912
rect 14188 12937 14197 12971
rect 14197 12937 14231 12971
rect 14231 12937 14240 12971
rect 14188 12928 14240 12937
rect 14556 12971 14608 12980
rect 14556 12937 14565 12971
rect 14565 12937 14599 12971
rect 14599 12937 14608 12971
rect 14556 12928 14608 12937
rect 24032 12928 24084 12980
rect 24492 12928 24544 12980
rect 24676 12928 24728 12980
rect 24768 12928 24820 12980
rect 7748 12724 7800 12776
rect 8116 12724 8168 12776
rect 11244 12792 11296 12844
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 13820 12792 13872 12844
rect 10876 12724 10928 12776
rect 15108 12792 15160 12844
rect 18144 12860 18196 12912
rect 18512 12860 18564 12912
rect 19432 12835 19484 12844
rect 19432 12801 19441 12835
rect 19441 12801 19475 12835
rect 19475 12801 19484 12835
rect 19432 12792 19484 12801
rect 7012 12656 7064 12708
rect 9588 12656 9640 12708
rect 9772 12656 9824 12708
rect 16028 12656 16080 12708
rect 5448 12588 5500 12640
rect 7840 12588 7892 12640
rect 8576 12631 8628 12640
rect 8576 12597 8585 12631
rect 8585 12597 8619 12631
rect 8619 12597 8628 12631
rect 8576 12588 8628 12597
rect 10600 12631 10652 12640
rect 10600 12597 10609 12631
rect 10609 12597 10643 12631
rect 10643 12597 10652 12631
rect 10600 12588 10652 12597
rect 11060 12588 11112 12640
rect 11244 12588 11296 12640
rect 12808 12588 12860 12640
rect 19340 12724 19392 12776
rect 18512 12699 18564 12708
rect 18512 12665 18521 12699
rect 18521 12665 18555 12699
rect 18555 12665 18564 12699
rect 18512 12656 18564 12665
rect 30564 12860 30616 12912
rect 31484 12928 31536 12980
rect 21916 12835 21968 12844
rect 21916 12801 21925 12835
rect 21925 12801 21959 12835
rect 21959 12801 21968 12835
rect 21916 12792 21968 12801
rect 22192 12724 22244 12776
rect 22652 12767 22704 12776
rect 22652 12733 22661 12767
rect 22661 12733 22695 12767
rect 22695 12733 22704 12767
rect 22652 12724 22704 12733
rect 22836 12724 22888 12776
rect 25412 12724 25464 12776
rect 31668 12860 31720 12912
rect 35440 12860 35492 12912
rect 38568 12860 38620 12912
rect 39028 12860 39080 12912
rect 32128 12835 32180 12844
rect 32128 12801 32137 12835
rect 32137 12801 32171 12835
rect 32171 12801 32180 12835
rect 32128 12792 32180 12801
rect 32680 12792 32732 12844
rect 35992 12792 36044 12844
rect 37556 12792 37608 12844
rect 35900 12724 35952 12776
rect 21456 12656 21508 12708
rect 30380 12656 30432 12708
rect 30564 12656 30616 12708
rect 41052 12860 41104 12912
rect 42432 12860 42484 12912
rect 46112 12928 46164 12980
rect 49056 12928 49108 12980
rect 52184 12971 52236 12980
rect 52184 12937 52193 12971
rect 52193 12937 52227 12971
rect 52227 12937 52236 12971
rect 52184 12928 52236 12937
rect 55036 12971 55088 12980
rect 55036 12937 55045 12971
rect 55045 12937 55079 12971
rect 55079 12937 55088 12971
rect 55036 12928 55088 12937
rect 56048 12971 56100 12980
rect 56048 12937 56057 12971
rect 56057 12937 56091 12971
rect 56091 12937 56100 12971
rect 56048 12928 56100 12937
rect 48044 12860 48096 12912
rect 51816 12860 51868 12912
rect 54576 12860 54628 12912
rect 55128 12860 55180 12912
rect 40776 12835 40828 12844
rect 40776 12801 40785 12835
rect 40785 12801 40819 12835
rect 40819 12801 40828 12835
rect 40776 12792 40828 12801
rect 42616 12835 42668 12844
rect 41052 12724 41104 12776
rect 42616 12801 42625 12835
rect 42625 12801 42659 12835
rect 42659 12801 42668 12835
rect 42616 12792 42668 12801
rect 44456 12792 44508 12844
rect 46204 12835 46256 12844
rect 46204 12801 46213 12835
rect 46213 12801 46247 12835
rect 46247 12801 46256 12835
rect 46204 12792 46256 12801
rect 48688 12835 48740 12844
rect 48688 12801 48697 12835
rect 48697 12801 48731 12835
rect 48731 12801 48740 12835
rect 48688 12792 48740 12801
rect 48872 12835 48924 12844
rect 48872 12801 48881 12835
rect 48881 12801 48915 12835
rect 48915 12801 48924 12835
rect 48872 12792 48924 12801
rect 50804 12835 50856 12844
rect 50804 12801 50813 12835
rect 50813 12801 50847 12835
rect 50847 12801 50856 12835
rect 50804 12792 50856 12801
rect 54852 12792 54904 12844
rect 56232 12835 56284 12844
rect 56232 12801 56241 12835
rect 56241 12801 56275 12835
rect 56275 12801 56284 12835
rect 56232 12792 56284 12801
rect 42892 12724 42944 12776
rect 43536 12767 43588 12776
rect 43536 12733 43545 12767
rect 43545 12733 43579 12767
rect 43579 12733 43588 12767
rect 43536 12724 43588 12733
rect 43720 12767 43772 12776
rect 43720 12733 43729 12767
rect 43729 12733 43763 12767
rect 43763 12733 43772 12767
rect 43720 12724 43772 12733
rect 55404 12724 55456 12776
rect 22928 12588 22980 12640
rect 23112 12588 23164 12640
rect 24860 12631 24912 12640
rect 24860 12597 24869 12631
rect 24869 12597 24903 12631
rect 24903 12597 24912 12631
rect 24860 12588 24912 12597
rect 25688 12588 25740 12640
rect 30840 12631 30892 12640
rect 30840 12597 30849 12631
rect 30849 12597 30883 12631
rect 30883 12597 30892 12631
rect 30840 12588 30892 12597
rect 33508 12631 33560 12640
rect 33508 12597 33517 12631
rect 33517 12597 33551 12631
rect 33551 12597 33560 12631
rect 33508 12588 33560 12597
rect 38844 12588 38896 12640
rect 39120 12588 39172 12640
rect 43996 12656 44048 12708
rect 43536 12588 43588 12640
rect 43628 12631 43680 12640
rect 43628 12597 43637 12631
rect 43637 12597 43671 12631
rect 43671 12597 43680 12631
rect 43628 12588 43680 12597
rect 51080 12588 51132 12640
rect 54668 12588 54720 12640
rect 56324 12588 56376 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 6644 12427 6696 12436
rect 6644 12393 6653 12427
rect 6653 12393 6687 12427
rect 6687 12393 6696 12427
rect 6644 12384 6696 12393
rect 15844 12384 15896 12436
rect 16396 12427 16448 12436
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 20812 12427 20864 12436
rect 20812 12393 20821 12427
rect 20821 12393 20855 12427
rect 20855 12393 20864 12427
rect 20812 12384 20864 12393
rect 21364 12384 21416 12436
rect 21916 12427 21968 12436
rect 21916 12393 21925 12427
rect 21925 12393 21959 12427
rect 21959 12393 21968 12427
rect 21916 12384 21968 12393
rect 3240 12359 3292 12368
rect 3240 12325 3249 12359
rect 3249 12325 3283 12359
rect 3283 12325 3292 12359
rect 3240 12316 3292 12325
rect 7196 12316 7248 12368
rect 6000 12248 6052 12300
rect 3424 12180 3476 12232
rect 8300 12248 8352 12300
rect 8576 12248 8628 12300
rect 10784 12316 10836 12368
rect 15200 12316 15252 12368
rect 19340 12316 19392 12368
rect 22284 12384 22336 12436
rect 23112 12427 23164 12436
rect 23112 12393 23121 12427
rect 23121 12393 23155 12427
rect 23155 12393 23164 12427
rect 23112 12384 23164 12393
rect 24032 12384 24084 12436
rect 24676 12384 24728 12436
rect 25596 12427 25648 12436
rect 25596 12393 25605 12427
rect 25605 12393 25639 12427
rect 25639 12393 25648 12427
rect 25596 12384 25648 12393
rect 9588 12248 9640 12300
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 7472 12180 7524 12232
rect 10232 12223 10284 12232
rect 2596 12112 2648 12164
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 16028 12248 16080 12300
rect 16396 12248 16448 12300
rect 17408 12248 17460 12300
rect 18052 12248 18104 12300
rect 18972 12248 19024 12300
rect 21548 12248 21600 12300
rect 23112 12248 23164 12300
rect 27436 12384 27488 12436
rect 29460 12384 29512 12436
rect 29828 12384 29880 12436
rect 31852 12427 31904 12436
rect 31852 12393 31861 12427
rect 31861 12393 31895 12427
rect 31895 12393 31904 12427
rect 31852 12384 31904 12393
rect 38752 12384 38804 12436
rect 39948 12384 40000 12436
rect 37280 12316 37332 12368
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 12440 12180 12492 12232
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 14740 12180 14792 12189
rect 15936 12180 15988 12232
rect 16304 12180 16356 12232
rect 13728 12112 13780 12164
rect 15568 12112 15620 12164
rect 21824 12180 21876 12232
rect 21088 12155 21140 12164
rect 21088 12121 21097 12155
rect 21097 12121 21131 12155
rect 21131 12121 21140 12155
rect 21088 12112 21140 12121
rect 21732 12112 21784 12164
rect 22376 12180 22428 12232
rect 22836 12180 22888 12232
rect 29460 12248 29512 12300
rect 28540 12180 28592 12232
rect 28908 12180 28960 12232
rect 36636 12248 36688 12300
rect 38016 12248 38068 12300
rect 42340 12316 42392 12368
rect 42524 12384 42576 12436
rect 43076 12384 43128 12436
rect 43260 12316 43312 12368
rect 31484 12223 31536 12232
rect 31484 12189 31493 12223
rect 31493 12189 31527 12223
rect 31527 12189 31536 12223
rect 31484 12180 31536 12189
rect 23480 12112 23532 12164
rect 24860 12112 24912 12164
rect 25596 12112 25648 12164
rect 26608 12112 26660 12164
rect 7472 12044 7524 12096
rect 7932 12044 7984 12096
rect 12624 12044 12676 12096
rect 13084 12044 13136 12096
rect 13636 12044 13688 12096
rect 16580 12044 16632 12096
rect 22744 12044 22796 12096
rect 25228 12044 25280 12096
rect 34520 12180 34572 12232
rect 35992 12180 36044 12232
rect 36728 12180 36780 12232
rect 38568 12223 38620 12232
rect 38568 12189 38601 12223
rect 38601 12189 38620 12223
rect 38568 12180 38620 12189
rect 38752 12223 38804 12232
rect 38752 12189 38761 12223
rect 38761 12189 38795 12223
rect 38795 12189 38804 12223
rect 38752 12180 38804 12189
rect 38844 12223 38896 12232
rect 38844 12189 38853 12223
rect 38853 12189 38887 12223
rect 38887 12189 38896 12223
rect 38844 12180 38896 12189
rect 39120 12180 39172 12232
rect 40776 12180 40828 12232
rect 42524 12180 42576 12232
rect 43260 12223 43312 12232
rect 43260 12189 43269 12223
rect 43269 12189 43303 12223
rect 43303 12189 43312 12223
rect 43720 12384 43772 12436
rect 48596 12384 48648 12436
rect 51172 12384 51224 12436
rect 51448 12384 51500 12436
rect 51908 12384 51960 12436
rect 48688 12316 48740 12368
rect 51264 12316 51316 12368
rect 52000 12359 52052 12368
rect 52000 12325 52009 12359
rect 52009 12325 52043 12359
rect 52043 12325 52052 12359
rect 52000 12316 52052 12325
rect 43260 12180 43312 12189
rect 43996 12223 44048 12232
rect 43996 12189 44005 12223
rect 44005 12189 44039 12223
rect 44039 12189 44048 12223
rect 43996 12180 44048 12189
rect 47400 12248 47452 12300
rect 47676 12180 47728 12232
rect 48320 12180 48372 12232
rect 51448 12248 51500 12300
rect 55588 12291 55640 12300
rect 55588 12257 55597 12291
rect 55597 12257 55631 12291
rect 55631 12257 55640 12291
rect 55588 12248 55640 12257
rect 48688 12180 48740 12232
rect 48780 12180 48832 12232
rect 28816 12044 28868 12096
rect 36452 12112 36504 12164
rect 36912 12112 36964 12164
rect 34796 12044 34848 12096
rect 35624 12044 35676 12096
rect 36544 12044 36596 12096
rect 38384 12087 38436 12096
rect 38384 12053 38393 12087
rect 38393 12053 38427 12087
rect 38427 12053 38436 12087
rect 38384 12044 38436 12053
rect 38476 12044 38528 12096
rect 41696 12112 41748 12164
rect 41880 12155 41932 12164
rect 41880 12121 41889 12155
rect 41889 12121 41923 12155
rect 41923 12121 41932 12155
rect 41880 12112 41932 12121
rect 55128 12180 55180 12232
rect 55404 12223 55456 12232
rect 55404 12189 55413 12223
rect 55413 12189 55447 12223
rect 55447 12189 55456 12223
rect 55404 12180 55456 12189
rect 52184 12112 52236 12164
rect 42708 12044 42760 12096
rect 43996 12044 44048 12096
rect 47860 12087 47912 12096
rect 47860 12053 47869 12087
rect 47869 12053 47903 12087
rect 47903 12053 47912 12087
rect 47860 12044 47912 12053
rect 51540 12044 51592 12096
rect 53932 12044 53984 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 2136 11840 2188 11892
rect 11428 11840 11480 11892
rect 11520 11840 11572 11892
rect 26884 11840 26936 11892
rect 26976 11840 27028 11892
rect 33508 11840 33560 11892
rect 33600 11840 33652 11892
rect 37096 11840 37148 11892
rect 41696 11840 41748 11892
rect 46572 11883 46624 11892
rect 5632 11815 5684 11824
rect 3240 11704 3292 11756
rect 3516 11747 3568 11756
rect 3516 11713 3525 11747
rect 3525 11713 3559 11747
rect 3559 11713 3568 11747
rect 3516 11704 3568 11713
rect 5632 11781 5641 11815
rect 5641 11781 5675 11815
rect 5675 11781 5684 11815
rect 5632 11772 5684 11781
rect 7472 11815 7524 11824
rect 7472 11781 7481 11815
rect 7481 11781 7515 11815
rect 7515 11781 7524 11815
rect 7472 11772 7524 11781
rect 12440 11772 12492 11824
rect 12624 11772 12676 11824
rect 15568 11815 15620 11824
rect 5908 11704 5960 11756
rect 8484 11704 8536 11756
rect 10048 11704 10100 11756
rect 10876 11704 10928 11756
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 9404 11636 9456 11688
rect 3608 11568 3660 11620
rect 8300 11568 8352 11620
rect 12256 11704 12308 11756
rect 13176 11747 13228 11756
rect 13176 11713 13185 11747
rect 13185 11713 13219 11747
rect 13219 11713 13228 11747
rect 13176 11704 13228 11713
rect 15568 11781 15577 11815
rect 15577 11781 15611 11815
rect 15611 11781 15620 11815
rect 15568 11772 15620 11781
rect 16028 11772 16080 11824
rect 22192 11772 22244 11824
rect 24124 11815 24176 11824
rect 24124 11781 24133 11815
rect 24133 11781 24167 11815
rect 24167 11781 24176 11815
rect 24124 11772 24176 11781
rect 24492 11772 24544 11824
rect 28632 11772 28684 11824
rect 41880 11772 41932 11824
rect 42892 11815 42944 11824
rect 42892 11781 42901 11815
rect 42901 11781 42935 11815
rect 42935 11781 42944 11815
rect 42892 11772 42944 11781
rect 43076 11772 43128 11824
rect 15936 11704 15988 11756
rect 16764 11704 16816 11756
rect 17132 11747 17184 11756
rect 17132 11713 17141 11747
rect 17141 11713 17175 11747
rect 17175 11713 17184 11747
rect 17132 11704 17184 11713
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 19156 11747 19208 11756
rect 19156 11713 19165 11747
rect 19165 11713 19199 11747
rect 19199 11713 19208 11747
rect 19156 11704 19208 11713
rect 19432 11704 19484 11756
rect 19984 11704 20036 11756
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22284 11747 22336 11756
rect 22100 11704 22152 11713
rect 22284 11713 22293 11747
rect 22293 11713 22327 11747
rect 22327 11713 22336 11747
rect 22284 11704 22336 11713
rect 23572 11704 23624 11756
rect 13360 11636 13412 11688
rect 15660 11679 15712 11688
rect 15660 11645 15669 11679
rect 15669 11645 15703 11679
rect 15703 11645 15712 11679
rect 15660 11636 15712 11645
rect 16672 11636 16724 11688
rect 16948 11636 17000 11688
rect 17040 11636 17092 11688
rect 21272 11636 21324 11688
rect 21548 11636 21600 11688
rect 26424 11704 26476 11756
rect 26516 11704 26568 11756
rect 24216 11636 24268 11688
rect 28816 11636 28868 11688
rect 13084 11611 13136 11620
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 9956 11500 10008 11552
rect 13084 11577 13093 11611
rect 13093 11577 13127 11611
rect 13127 11577 13136 11611
rect 13084 11568 13136 11577
rect 12532 11500 12584 11552
rect 13728 11500 13780 11552
rect 14280 11500 14332 11552
rect 17040 11500 17092 11552
rect 18788 11543 18840 11552
rect 18788 11509 18797 11543
rect 18797 11509 18831 11543
rect 18831 11509 18840 11543
rect 18788 11500 18840 11509
rect 21824 11543 21876 11552
rect 21824 11509 21833 11543
rect 21833 11509 21867 11543
rect 21867 11509 21876 11543
rect 21824 11500 21876 11509
rect 24216 11500 24268 11552
rect 24952 11500 25004 11552
rect 29920 11704 29972 11756
rect 31116 11704 31168 11756
rect 31484 11704 31536 11756
rect 32680 11704 32732 11756
rect 36176 11704 36228 11756
rect 36360 11747 36412 11756
rect 36360 11713 36369 11747
rect 36369 11713 36403 11747
rect 36403 11713 36412 11747
rect 36360 11704 36412 11713
rect 36544 11704 36596 11756
rect 42616 11704 42668 11756
rect 29276 11679 29328 11688
rect 29276 11645 29285 11679
rect 29285 11645 29319 11679
rect 29319 11645 29328 11679
rect 29460 11679 29512 11688
rect 29276 11636 29328 11645
rect 29460 11645 29469 11679
rect 29469 11645 29503 11679
rect 29503 11645 29512 11679
rect 29460 11636 29512 11645
rect 29828 11636 29880 11688
rect 30104 11568 30156 11620
rect 33600 11568 33652 11620
rect 35900 11611 35952 11620
rect 35900 11577 35909 11611
rect 35909 11577 35943 11611
rect 35943 11577 35952 11611
rect 35900 11568 35952 11577
rect 35992 11568 36044 11620
rect 42524 11568 42576 11620
rect 28632 11543 28684 11552
rect 28632 11509 28641 11543
rect 28641 11509 28675 11543
rect 28675 11509 28684 11543
rect 28632 11500 28684 11509
rect 29552 11500 29604 11552
rect 30840 11500 30892 11552
rect 36544 11543 36596 11552
rect 36544 11509 36553 11543
rect 36553 11509 36587 11543
rect 36587 11509 36596 11543
rect 36544 11500 36596 11509
rect 40316 11500 40368 11552
rect 41052 11500 41104 11552
rect 43260 11704 43312 11756
rect 43996 11772 44048 11824
rect 46572 11849 46581 11883
rect 46581 11849 46615 11883
rect 46615 11849 46624 11883
rect 46572 11840 46624 11849
rect 48412 11840 48464 11892
rect 48688 11840 48740 11892
rect 53932 11815 53984 11824
rect 46020 11704 46072 11756
rect 46572 11704 46624 11756
rect 48780 11704 48832 11756
rect 51448 11747 51500 11756
rect 48596 11636 48648 11688
rect 51448 11713 51457 11747
rect 51457 11713 51491 11747
rect 51491 11713 51500 11747
rect 51448 11704 51500 11713
rect 51540 11679 51592 11688
rect 51540 11645 51549 11679
rect 51549 11645 51583 11679
rect 51583 11645 51592 11679
rect 51540 11636 51592 11645
rect 53932 11781 53941 11815
rect 53941 11781 53975 11815
rect 53975 11781 53984 11815
rect 53932 11772 53984 11781
rect 52000 11704 52052 11756
rect 55404 11840 55456 11892
rect 55128 11772 55180 11824
rect 51356 11568 51408 11620
rect 48688 11543 48740 11552
rect 48688 11509 48697 11543
rect 48697 11509 48731 11543
rect 48731 11509 48740 11543
rect 48688 11500 48740 11509
rect 48872 11500 48924 11552
rect 54668 11679 54720 11688
rect 54668 11645 54677 11679
rect 54677 11645 54711 11679
rect 54711 11645 54720 11679
rect 54668 11636 54720 11645
rect 55588 11500 55640 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 8024 11296 8076 11348
rect 12440 11296 12492 11348
rect 14372 11296 14424 11348
rect 16856 11296 16908 11348
rect 21548 11339 21600 11348
rect 21548 11305 21557 11339
rect 21557 11305 21591 11339
rect 21591 11305 21600 11339
rect 21548 11296 21600 11305
rect 23572 11339 23624 11348
rect 12624 11228 12676 11280
rect 2044 11160 2096 11212
rect 2596 11160 2648 11212
rect 10876 11160 10928 11212
rect 13176 11228 13228 11280
rect 15660 11228 15712 11280
rect 15936 11228 15988 11280
rect 22928 11228 22980 11280
rect 23112 11228 23164 11280
rect 23572 11305 23581 11339
rect 23581 11305 23615 11339
rect 23615 11305 23624 11339
rect 23572 11296 23624 11305
rect 34796 11339 34848 11348
rect 34796 11305 34805 11339
rect 34805 11305 34839 11339
rect 34839 11305 34848 11339
rect 34796 11296 34848 11305
rect 24492 11228 24544 11280
rect 26884 11228 26936 11280
rect 35072 11228 35124 11280
rect 2136 11092 2188 11144
rect 9956 11092 10008 11144
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 11520 11092 11572 11144
rect 12256 11092 12308 11144
rect 12624 11092 12676 11144
rect 13452 11160 13504 11212
rect 13728 11092 13780 11144
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 16396 11160 16448 11212
rect 17132 11160 17184 11212
rect 18052 11203 18104 11212
rect 18052 11169 18061 11203
rect 18061 11169 18095 11203
rect 18095 11169 18104 11203
rect 18052 11160 18104 11169
rect 16856 11092 16908 11144
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 2596 11024 2648 11076
rect 4896 11024 4948 11076
rect 6920 11024 6972 11076
rect 7932 11024 7984 11076
rect 9404 11067 9456 11076
rect 9404 11033 9413 11067
rect 9413 11033 9447 11067
rect 9447 11033 9456 11067
rect 9404 11024 9456 11033
rect 2504 10999 2556 11008
rect 2504 10965 2513 10999
rect 2513 10965 2547 10999
rect 2547 10965 2556 10999
rect 2504 10956 2556 10965
rect 7012 10956 7064 11008
rect 10140 10999 10192 11008
rect 10140 10965 10149 10999
rect 10149 10965 10183 10999
rect 10183 10965 10192 10999
rect 10140 10956 10192 10965
rect 11796 11024 11848 11076
rect 12900 11067 12952 11076
rect 12900 11033 12909 11067
rect 12909 11033 12943 11067
rect 12943 11033 12952 11067
rect 12900 11024 12952 11033
rect 16488 11024 16540 11076
rect 19432 11092 19484 11144
rect 22560 11160 22612 11212
rect 26056 11160 26108 11212
rect 29552 11160 29604 11212
rect 22284 11092 22336 11144
rect 21180 11067 21232 11076
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 27436 11092 27488 11144
rect 28632 11092 28684 11144
rect 29920 11160 29972 11212
rect 35440 11296 35492 11348
rect 36176 11339 36228 11348
rect 36176 11305 36185 11339
rect 36185 11305 36219 11339
rect 36219 11305 36228 11339
rect 36176 11296 36228 11305
rect 36820 11296 36872 11348
rect 43076 11296 43128 11348
rect 43260 11339 43312 11348
rect 43260 11305 43269 11339
rect 43269 11305 43303 11339
rect 43303 11305 43312 11339
rect 43260 11296 43312 11305
rect 44456 11296 44508 11348
rect 15568 10956 15620 11008
rect 21732 10956 21784 11008
rect 24860 11024 24912 11076
rect 25228 11024 25280 11076
rect 28540 11067 28592 11076
rect 28540 11033 28549 11067
rect 28549 11033 28583 11067
rect 28583 11033 28592 11067
rect 28540 11024 28592 11033
rect 29460 11024 29512 11076
rect 29828 11135 29880 11144
rect 29828 11101 29837 11135
rect 29837 11101 29871 11135
rect 29871 11101 29880 11135
rect 30104 11135 30156 11144
rect 29828 11092 29880 11101
rect 30104 11101 30113 11135
rect 30113 11101 30147 11135
rect 30147 11101 30156 11135
rect 30104 11092 30156 11101
rect 33784 11092 33836 11144
rect 39948 11228 40000 11280
rect 40592 11228 40644 11280
rect 29920 11067 29972 11076
rect 29920 11033 29929 11067
rect 29929 11033 29963 11067
rect 29963 11033 29972 11067
rect 29920 11024 29972 11033
rect 34152 10956 34204 11008
rect 35440 10956 35492 11008
rect 36544 11160 36596 11212
rect 36176 11135 36228 11144
rect 36176 11101 36185 11135
rect 36185 11101 36219 11135
rect 36219 11101 36228 11135
rect 36176 11092 36228 11101
rect 36820 11092 36872 11144
rect 38384 11160 38436 11212
rect 36084 11024 36136 11076
rect 36360 11024 36412 11076
rect 38936 11092 38988 11144
rect 40868 11092 40920 11144
rect 41052 11135 41104 11144
rect 41052 11101 41061 11135
rect 41061 11101 41095 11135
rect 41095 11101 41104 11135
rect 41052 11092 41104 11101
rect 42708 11135 42760 11144
rect 37096 11024 37148 11076
rect 40776 11067 40828 11076
rect 35716 10956 35768 11008
rect 36176 10956 36228 11008
rect 36544 10956 36596 11008
rect 40776 11033 40785 11067
rect 40785 11033 40819 11067
rect 40819 11033 40828 11067
rect 40776 11024 40828 11033
rect 42708 11101 42717 11135
rect 42717 11101 42751 11135
rect 42751 11101 42760 11135
rect 42708 11092 42760 11101
rect 43628 11160 43680 11212
rect 43076 11135 43128 11144
rect 43076 11101 43085 11135
rect 43085 11101 43119 11135
rect 43119 11101 43128 11135
rect 43076 11092 43128 11101
rect 43720 11092 43772 11144
rect 47676 11135 47728 11144
rect 47676 11101 47685 11135
rect 47685 11101 47719 11135
rect 47719 11101 47728 11135
rect 47676 11092 47728 11101
rect 43168 11024 43220 11076
rect 48596 11271 48648 11280
rect 48596 11237 48605 11271
rect 48605 11237 48639 11271
rect 48639 11237 48648 11271
rect 48596 11228 48648 11237
rect 51632 11228 51684 11280
rect 48412 11135 48464 11144
rect 48412 11101 48421 11135
rect 48421 11101 48455 11135
rect 48455 11101 48464 11135
rect 48412 11092 48464 11101
rect 51356 11135 51408 11144
rect 51356 11101 51365 11135
rect 51365 11101 51399 11135
rect 51399 11101 51408 11135
rect 51356 11092 51408 11101
rect 51540 11092 51592 11144
rect 51448 10956 51500 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4896 10795 4948 10804
rect 4896 10761 4905 10795
rect 4905 10761 4939 10795
rect 4939 10761 4948 10795
rect 4896 10752 4948 10761
rect 5448 10752 5500 10804
rect 2504 10684 2556 10736
rect 2596 10684 2648 10736
rect 12808 10752 12860 10804
rect 13268 10752 13320 10804
rect 15568 10795 15620 10804
rect 15568 10761 15577 10795
rect 15577 10761 15611 10795
rect 15611 10761 15620 10795
rect 15568 10752 15620 10761
rect 10140 10684 10192 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 5080 10659 5132 10668
rect 5080 10625 5089 10659
rect 5089 10625 5123 10659
rect 5123 10625 5132 10659
rect 5080 10616 5132 10625
rect 5724 10616 5776 10668
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 7288 10616 7340 10668
rect 8024 10616 8076 10668
rect 11796 10616 11848 10668
rect 12164 10616 12216 10668
rect 11520 10591 11572 10600
rect 7472 10480 7524 10532
rect 1400 10455 1452 10464
rect 1400 10421 1409 10455
rect 1409 10421 1443 10455
rect 1443 10421 1452 10455
rect 1400 10412 1452 10421
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 10600 10523 10652 10532
rect 10600 10489 10609 10523
rect 10609 10489 10643 10523
rect 10643 10489 10652 10523
rect 12256 10548 12308 10600
rect 10600 10480 10652 10489
rect 12348 10480 12400 10532
rect 12900 10616 12952 10668
rect 13452 10616 13504 10668
rect 14740 10684 14792 10736
rect 17868 10684 17920 10736
rect 18788 10684 18840 10736
rect 16764 10616 16816 10668
rect 16856 10659 16908 10668
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 19156 10616 19208 10668
rect 22100 10752 22152 10804
rect 23112 10752 23164 10804
rect 24860 10752 24912 10804
rect 40316 10795 40368 10804
rect 40316 10761 40325 10795
rect 40325 10761 40359 10795
rect 40359 10761 40368 10795
rect 40316 10752 40368 10761
rect 40868 10752 40920 10804
rect 48320 10752 48372 10804
rect 21180 10684 21232 10736
rect 22192 10684 22244 10736
rect 22284 10727 22336 10736
rect 22284 10693 22293 10727
rect 22293 10693 22327 10727
rect 22327 10693 22336 10727
rect 38660 10727 38712 10736
rect 22284 10684 22336 10693
rect 38660 10693 38669 10727
rect 38669 10693 38703 10727
rect 38703 10693 38712 10727
rect 38660 10684 38712 10693
rect 21732 10616 21784 10668
rect 22560 10616 22612 10668
rect 24952 10616 25004 10668
rect 27896 10659 27948 10668
rect 27896 10625 27905 10659
rect 27905 10625 27939 10659
rect 27939 10625 27948 10659
rect 27896 10616 27948 10625
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 15752 10591 15804 10600
rect 13268 10548 13320 10557
rect 15752 10557 15761 10591
rect 15761 10557 15795 10591
rect 15795 10557 15804 10591
rect 15752 10548 15804 10557
rect 15936 10591 15988 10600
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 16488 10548 16540 10600
rect 17132 10591 17184 10600
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 17408 10548 17460 10600
rect 18144 10591 18196 10600
rect 18144 10557 18153 10591
rect 18153 10557 18187 10591
rect 18187 10557 18196 10591
rect 18144 10548 18196 10557
rect 9496 10412 9548 10464
rect 10968 10412 11020 10464
rect 12808 10412 12860 10464
rect 13728 10412 13780 10464
rect 16672 10455 16724 10464
rect 16672 10421 16681 10455
rect 16681 10421 16715 10455
rect 16715 10421 16724 10455
rect 16672 10412 16724 10421
rect 27620 10548 27672 10600
rect 29920 10616 29972 10668
rect 30748 10616 30800 10668
rect 38476 10659 38528 10668
rect 38476 10625 38485 10659
rect 38485 10625 38519 10659
rect 38519 10625 38528 10659
rect 39120 10659 39172 10668
rect 38476 10616 38528 10625
rect 39120 10625 39129 10659
rect 39129 10625 39163 10659
rect 39163 10625 39172 10659
rect 39120 10616 39172 10625
rect 39580 10616 39632 10668
rect 47584 10616 47636 10668
rect 24952 10480 25004 10532
rect 25596 10480 25648 10532
rect 47124 10548 47176 10600
rect 31208 10480 31260 10532
rect 21732 10412 21784 10464
rect 27988 10455 28040 10464
rect 27988 10421 27997 10455
rect 27997 10421 28031 10455
rect 28031 10421 28040 10455
rect 27988 10412 28040 10421
rect 31484 10455 31536 10464
rect 31484 10421 31493 10455
rect 31493 10421 31527 10455
rect 31527 10421 31536 10455
rect 31484 10412 31536 10421
rect 38568 10412 38620 10464
rect 38844 10412 38896 10464
rect 40776 10480 40828 10532
rect 39580 10455 39632 10464
rect 39580 10421 39589 10455
rect 39589 10421 39623 10455
rect 39623 10421 39632 10455
rect 39580 10412 39632 10421
rect 40592 10455 40644 10464
rect 40592 10421 40601 10455
rect 40601 10421 40635 10455
rect 40635 10421 40644 10455
rect 40592 10412 40644 10421
rect 41328 10412 41380 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2136 10251 2188 10260
rect 2136 10217 2145 10251
rect 2145 10217 2179 10251
rect 2179 10217 2188 10251
rect 2136 10208 2188 10217
rect 3424 10208 3476 10260
rect 7288 10251 7340 10260
rect 7288 10217 7297 10251
rect 7297 10217 7331 10251
rect 7331 10217 7340 10251
rect 7288 10208 7340 10217
rect 10048 10208 10100 10260
rect 10232 10208 10284 10260
rect 11520 10208 11572 10260
rect 13268 10208 13320 10260
rect 15752 10208 15804 10260
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 6368 10072 6420 10124
rect 6828 10072 6880 10124
rect 3332 10004 3384 10056
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 6736 10004 6788 10056
rect 8484 10140 8536 10192
rect 38016 10208 38068 10260
rect 38476 10208 38528 10260
rect 39120 10251 39172 10260
rect 39120 10217 39129 10251
rect 39129 10217 39163 10251
rect 39163 10217 39172 10251
rect 39120 10208 39172 10217
rect 40776 10208 40828 10260
rect 47584 10251 47636 10260
rect 47584 10217 47593 10251
rect 47593 10217 47627 10251
rect 47627 10217 47636 10251
rect 47584 10208 47636 10217
rect 47860 10208 47912 10260
rect 51448 10208 51500 10260
rect 7196 10072 7248 10124
rect 7656 10004 7708 10056
rect 9772 10004 9824 10056
rect 22468 10140 22520 10192
rect 42248 10140 42300 10192
rect 48688 10140 48740 10192
rect 13728 10072 13780 10124
rect 16856 10072 16908 10124
rect 18052 10072 18104 10124
rect 26332 10072 26384 10124
rect 27436 10115 27488 10124
rect 27436 10081 27445 10115
rect 27445 10081 27479 10115
rect 27479 10081 27488 10115
rect 27436 10072 27488 10081
rect 31668 10072 31720 10124
rect 42432 10072 42484 10124
rect 48044 10115 48096 10124
rect 48044 10081 48053 10115
rect 48053 10081 48087 10115
rect 48087 10081 48096 10115
rect 48044 10072 48096 10081
rect 51080 10072 51132 10124
rect 51540 10115 51592 10124
rect 51540 10081 51549 10115
rect 51549 10081 51583 10115
rect 51583 10081 51592 10115
rect 51540 10072 51592 10081
rect 7472 9936 7524 9988
rect 8484 9936 8536 9988
rect 13360 10004 13412 10056
rect 14096 10004 14148 10056
rect 15844 10004 15896 10056
rect 16488 10004 16540 10056
rect 20076 10004 20128 10056
rect 21916 10004 21968 10056
rect 11060 9868 11112 9920
rect 12164 9868 12216 9920
rect 13452 9868 13504 9920
rect 16304 9868 16356 9920
rect 21732 9936 21784 9988
rect 22468 10047 22520 10056
rect 22468 10013 22482 10047
rect 22482 10013 22516 10047
rect 22516 10013 22520 10047
rect 22468 10004 22520 10013
rect 24584 10004 24636 10056
rect 24952 10047 25004 10056
rect 24952 10013 24959 10047
rect 24959 10013 25004 10047
rect 24952 10004 25004 10013
rect 25044 10047 25096 10056
rect 25044 10013 25053 10047
rect 25053 10013 25087 10047
rect 25087 10013 25096 10047
rect 25044 10004 25096 10013
rect 25228 10047 25280 10056
rect 25228 10013 25242 10047
rect 25242 10013 25276 10047
rect 25276 10013 25280 10047
rect 30932 10047 30984 10056
rect 25228 10004 25280 10013
rect 30932 10013 30941 10047
rect 30941 10013 30975 10047
rect 30975 10013 30984 10047
rect 30932 10004 30984 10013
rect 23664 9936 23716 9988
rect 22744 9868 22796 9920
rect 23388 9868 23440 9920
rect 28080 9936 28132 9988
rect 36452 10004 36504 10056
rect 37648 10047 37700 10056
rect 37648 10013 37657 10047
rect 37657 10013 37691 10047
rect 37691 10013 37700 10047
rect 37648 10004 37700 10013
rect 38844 10047 38896 10056
rect 36544 9936 36596 9988
rect 37188 9979 37240 9988
rect 37188 9945 37197 9979
rect 37197 9945 37231 9979
rect 37231 9945 37240 9979
rect 37188 9936 37240 9945
rect 37280 9936 37332 9988
rect 38844 10013 38853 10047
rect 38853 10013 38887 10047
rect 38887 10013 38896 10047
rect 38844 10004 38896 10013
rect 41236 10047 41288 10056
rect 41236 10013 41245 10047
rect 41245 10013 41279 10047
rect 41279 10013 41288 10047
rect 41236 10004 41288 10013
rect 41328 10004 41380 10056
rect 37924 9936 37976 9988
rect 44640 9936 44692 9988
rect 46572 10004 46624 10056
rect 46480 9936 46532 9988
rect 51632 10004 51684 10056
rect 48780 9936 48832 9988
rect 28172 9868 28224 9920
rect 28816 9911 28868 9920
rect 28816 9877 28825 9911
rect 28825 9877 28859 9911
rect 28859 9877 28868 9911
rect 28816 9868 28868 9877
rect 30748 9868 30800 9920
rect 36452 9868 36504 9920
rect 37464 9868 37516 9920
rect 38936 9868 38988 9920
rect 45928 9911 45980 9920
rect 45928 9877 45937 9911
rect 45937 9877 45971 9911
rect 45971 9877 45980 9911
rect 45928 9868 45980 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 1400 9664 1452 9716
rect 5080 9664 5132 9716
rect 3332 9596 3384 9648
rect 10600 9596 10652 9648
rect 12532 9596 12584 9648
rect 8208 9528 8260 9580
rect 9956 9528 10008 9580
rect 12440 9571 12492 9580
rect 12440 9537 12449 9571
rect 12449 9537 12483 9571
rect 12483 9537 12492 9571
rect 12440 9528 12492 9537
rect 13360 9528 13412 9580
rect 14924 9596 14976 9648
rect 16672 9664 16724 9716
rect 17224 9596 17276 9648
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 4896 9460 4948 9512
rect 7196 9460 7248 9512
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 11060 9460 11112 9512
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 6000 9392 6052 9444
rect 7288 9435 7340 9444
rect 7288 9401 7297 9435
rect 7297 9401 7331 9435
rect 7331 9401 7340 9435
rect 7288 9392 7340 9401
rect 8300 9392 8352 9444
rect 8484 9435 8536 9444
rect 8484 9401 8493 9435
rect 8493 9401 8527 9435
rect 8527 9401 8536 9435
rect 8484 9392 8536 9401
rect 14096 9392 14148 9444
rect 14924 9392 14976 9444
rect 15844 9503 15896 9512
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 15844 9460 15896 9469
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 2412 9324 2464 9376
rect 9864 9324 9916 9376
rect 15568 9324 15620 9376
rect 21824 9596 21876 9648
rect 22284 9664 22336 9716
rect 23112 9664 23164 9716
rect 28080 9707 28132 9716
rect 28080 9673 28089 9707
rect 28089 9673 28123 9707
rect 28123 9673 28132 9707
rect 28080 9664 28132 9673
rect 30932 9707 30984 9716
rect 23204 9596 23256 9648
rect 23388 9596 23440 9648
rect 18144 9528 18196 9580
rect 19156 9528 19208 9580
rect 19340 9528 19392 9580
rect 28816 9634 28868 9686
rect 28908 9634 28960 9686
rect 30932 9673 30941 9707
rect 30941 9673 30975 9707
rect 30975 9673 30984 9707
rect 30932 9664 30984 9673
rect 31208 9664 31260 9716
rect 42248 9664 42300 9716
rect 42432 9707 42484 9716
rect 42432 9673 42441 9707
rect 42441 9673 42475 9707
rect 42475 9673 42484 9707
rect 42432 9664 42484 9673
rect 31484 9639 31536 9648
rect 24676 9503 24728 9512
rect 19432 9392 19484 9444
rect 18144 9324 18196 9376
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 25228 9460 25280 9512
rect 25688 9460 25740 9512
rect 27988 9528 28040 9580
rect 28632 9460 28684 9512
rect 28908 9460 28960 9512
rect 31484 9605 31493 9639
rect 31493 9605 31527 9639
rect 31527 9605 31536 9639
rect 31484 9596 31536 9605
rect 33140 9596 33192 9648
rect 33324 9596 33376 9648
rect 34060 9596 34112 9648
rect 36820 9596 36872 9648
rect 37648 9596 37700 9648
rect 42800 9639 42852 9648
rect 42800 9605 42809 9639
rect 42809 9605 42843 9639
rect 42843 9605 42852 9639
rect 45928 9639 45980 9648
rect 42800 9596 42852 9605
rect 45928 9605 45962 9639
rect 45962 9605 45980 9639
rect 45928 9596 45980 9605
rect 33600 9571 33652 9580
rect 33600 9537 33623 9571
rect 33623 9537 33652 9571
rect 33600 9528 33652 9537
rect 36544 9571 36596 9580
rect 36544 9537 36556 9571
rect 36556 9537 36590 9571
rect 36590 9537 36596 9571
rect 37280 9571 37332 9580
rect 36544 9528 36596 9537
rect 37280 9537 37289 9571
rect 37289 9537 37323 9571
rect 37323 9537 37332 9571
rect 37280 9528 37332 9537
rect 38936 9571 38988 9580
rect 38936 9537 38945 9571
rect 38945 9537 38979 9571
rect 38979 9537 38988 9571
rect 38936 9528 38988 9537
rect 39580 9571 39632 9580
rect 39580 9537 39589 9571
rect 39589 9537 39623 9571
rect 39623 9537 39632 9571
rect 39580 9528 39632 9537
rect 39764 9571 39816 9580
rect 39764 9537 39773 9571
rect 39773 9537 39807 9571
rect 39807 9537 39816 9571
rect 39764 9528 39816 9537
rect 42616 9571 42668 9580
rect 42616 9537 42625 9571
rect 42625 9537 42659 9571
rect 42659 9537 42668 9571
rect 42616 9528 42668 9537
rect 42708 9571 42760 9580
rect 42708 9537 42717 9571
rect 42717 9537 42751 9571
rect 42751 9537 42760 9571
rect 42708 9528 42760 9537
rect 42892 9571 42944 9580
rect 42892 9537 42927 9571
rect 42927 9537 42944 9571
rect 42892 9528 42944 9537
rect 31852 9460 31904 9512
rect 32680 9460 32732 9512
rect 22468 9324 22520 9376
rect 23204 9367 23256 9376
rect 23204 9333 23213 9367
rect 23213 9333 23247 9367
rect 23247 9333 23256 9367
rect 23204 9324 23256 9333
rect 23388 9324 23440 9376
rect 26148 9367 26200 9376
rect 26148 9333 26157 9367
rect 26157 9333 26191 9367
rect 26191 9333 26200 9367
rect 26148 9324 26200 9333
rect 33140 9392 33192 9444
rect 42800 9460 42852 9512
rect 47124 9528 47176 9580
rect 49700 9596 49752 9648
rect 30196 9324 30248 9376
rect 30840 9324 30892 9376
rect 35348 9324 35400 9376
rect 35808 9367 35860 9376
rect 35808 9333 35817 9367
rect 35817 9333 35851 9367
rect 35851 9333 35860 9367
rect 35808 9324 35860 9333
rect 36176 9324 36228 9376
rect 36728 9367 36780 9376
rect 36728 9333 36737 9367
rect 36737 9333 36771 9367
rect 36771 9333 36780 9367
rect 36728 9324 36780 9333
rect 36820 9324 36872 9376
rect 39764 9392 39816 9444
rect 39856 9392 39908 9444
rect 49516 9460 49568 9512
rect 43168 9392 43220 9444
rect 45376 9392 45428 9444
rect 38476 9324 38528 9376
rect 41696 9324 41748 9376
rect 46296 9324 46348 9376
rect 47032 9367 47084 9376
rect 47032 9333 47041 9367
rect 47041 9333 47075 9367
rect 47075 9333 47084 9367
rect 47032 9324 47084 9333
rect 48504 9324 48556 9376
rect 49424 9367 49476 9376
rect 49424 9333 49433 9367
rect 49433 9333 49467 9367
rect 49467 9333 49476 9367
rect 49424 9324 49476 9333
rect 49608 9367 49660 9376
rect 49608 9333 49617 9367
rect 49617 9333 49651 9367
rect 49651 9333 49660 9367
rect 49608 9324 49660 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 5908 9163 5960 9172
rect 5908 9129 5917 9163
rect 5917 9129 5951 9163
rect 5951 9129 5960 9163
rect 5908 9120 5960 9129
rect 8208 9163 8260 9172
rect 8208 9129 8217 9163
rect 8217 9129 8251 9163
rect 8251 9129 8260 9163
rect 8208 9120 8260 9129
rect 9404 9120 9456 9172
rect 10048 9163 10100 9172
rect 10048 9129 10057 9163
rect 10057 9129 10091 9163
rect 10091 9129 10100 9163
rect 10048 9120 10100 9129
rect 10324 9163 10376 9172
rect 10324 9129 10333 9163
rect 10333 9129 10367 9163
rect 10367 9129 10376 9163
rect 10324 9120 10376 9129
rect 13544 9163 13596 9172
rect 13544 9129 13553 9163
rect 13553 9129 13587 9163
rect 13587 9129 13596 9163
rect 13544 9120 13596 9129
rect 13728 9120 13780 9172
rect 19156 9120 19208 9172
rect 1860 8984 1912 9036
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 4620 8916 4672 8968
rect 5172 8848 5224 8900
rect 8852 8916 8904 8968
rect 9864 8959 9916 8968
rect 9864 8925 9873 8959
rect 9873 8925 9907 8959
rect 9907 8925 9916 8959
rect 9864 8916 9916 8925
rect 13084 9052 13136 9104
rect 13084 8959 13136 8968
rect 13084 8925 13091 8959
rect 13091 8925 13136 8959
rect 13084 8916 13136 8925
rect 13452 9052 13504 9104
rect 13268 8984 13320 9036
rect 13544 8916 13596 8968
rect 10048 8848 10100 8900
rect 13268 8891 13320 8900
rect 13268 8857 13277 8891
rect 13277 8857 13311 8891
rect 13311 8857 13320 8891
rect 14096 8891 14148 8900
rect 13268 8848 13320 8857
rect 14096 8857 14105 8891
rect 14105 8857 14139 8891
rect 14139 8857 14148 8891
rect 14096 8848 14148 8857
rect 2044 8780 2096 8832
rect 2228 8823 2280 8832
rect 2228 8789 2237 8823
rect 2237 8789 2271 8823
rect 2271 8789 2280 8823
rect 2228 8780 2280 8789
rect 5816 8780 5868 8832
rect 19340 8984 19392 9036
rect 14832 8780 14884 8832
rect 15016 8823 15068 8832
rect 15016 8789 15025 8823
rect 15025 8789 15059 8823
rect 15059 8789 15068 8823
rect 15016 8780 15068 8789
rect 15752 8916 15804 8968
rect 15936 8916 15988 8968
rect 15844 8848 15896 8900
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 17408 8916 17460 8968
rect 20168 9052 20220 9104
rect 21732 9052 21784 9104
rect 22560 9120 22612 9172
rect 23204 9120 23256 9172
rect 25136 9120 25188 9172
rect 33600 9120 33652 9172
rect 33876 9120 33928 9172
rect 37372 9120 37424 9172
rect 37556 9120 37608 9172
rect 39856 9120 39908 9172
rect 41788 9120 41840 9172
rect 42248 9120 42300 9172
rect 46204 9120 46256 9172
rect 46296 9163 46348 9172
rect 46296 9129 46305 9163
rect 46305 9129 46339 9163
rect 46339 9129 46348 9163
rect 46296 9120 46348 9129
rect 23020 9052 23072 9104
rect 24768 9052 24820 9104
rect 19984 8916 20036 8968
rect 16856 8848 16908 8900
rect 17040 8848 17092 8900
rect 24676 8984 24728 9036
rect 28908 9052 28960 9104
rect 44548 9052 44600 9104
rect 44732 9052 44784 9104
rect 33600 8984 33652 9036
rect 22560 8916 22612 8968
rect 22652 8916 22704 8968
rect 21916 8848 21968 8900
rect 24584 8916 24636 8968
rect 25044 8959 25096 8968
rect 23204 8848 23256 8900
rect 25044 8925 25053 8959
rect 25053 8925 25087 8959
rect 25087 8925 25096 8959
rect 25044 8916 25096 8925
rect 25228 8959 25280 8968
rect 25228 8925 25242 8959
rect 25242 8925 25276 8959
rect 25276 8925 25280 8959
rect 25228 8916 25280 8925
rect 27804 8916 27856 8968
rect 28816 8916 28868 8968
rect 28908 8916 28960 8968
rect 33508 8959 33560 8968
rect 33508 8925 33517 8959
rect 33517 8925 33551 8959
rect 33551 8925 33560 8959
rect 33508 8916 33560 8925
rect 33876 8916 33928 8968
rect 34060 8916 34112 8968
rect 34244 8916 34296 8968
rect 36268 8916 36320 8968
rect 37464 9027 37516 9036
rect 36636 8959 36688 8968
rect 26056 8848 26108 8900
rect 27712 8848 27764 8900
rect 16580 8780 16632 8832
rect 19432 8780 19484 8832
rect 22100 8780 22152 8832
rect 22744 8780 22796 8832
rect 27896 8780 27948 8832
rect 28540 8848 28592 8900
rect 28908 8780 28960 8832
rect 33692 8891 33744 8900
rect 33692 8857 33701 8891
rect 33701 8857 33735 8891
rect 33735 8857 33744 8891
rect 33692 8848 33744 8857
rect 35532 8848 35584 8900
rect 36636 8925 36645 8959
rect 36645 8925 36679 8959
rect 36679 8925 36688 8959
rect 36636 8916 36688 8925
rect 37188 8916 37240 8968
rect 37464 8993 37473 9027
rect 37473 8993 37507 9027
rect 37507 8993 37516 9027
rect 37464 8984 37516 8993
rect 37648 8916 37700 8968
rect 37740 8959 37792 8968
rect 37740 8925 37749 8959
rect 37749 8925 37783 8959
rect 37783 8925 37792 8959
rect 41512 8984 41564 9036
rect 37740 8916 37792 8925
rect 39120 8916 39172 8968
rect 37004 8848 37056 8900
rect 41880 8848 41932 8900
rect 42432 8916 42484 8968
rect 45008 8984 45060 9036
rect 43168 8916 43220 8968
rect 44916 8916 44968 8968
rect 45376 8984 45428 9036
rect 46664 8984 46716 9036
rect 51540 9027 51592 9036
rect 51540 8993 51549 9027
rect 51549 8993 51583 9027
rect 51583 8993 51592 9027
rect 51540 8984 51592 8993
rect 34796 8780 34848 8832
rect 36360 8780 36412 8832
rect 36912 8780 36964 8832
rect 38752 8780 38804 8832
rect 42248 8848 42300 8900
rect 44180 8848 44232 8900
rect 45468 8891 45520 8900
rect 47032 8916 47084 8968
rect 47124 8916 47176 8968
rect 45468 8857 45503 8891
rect 45503 8857 45520 8891
rect 45468 8848 45520 8857
rect 46296 8891 46348 8900
rect 46296 8857 46337 8891
rect 46337 8857 46348 8891
rect 49700 8916 49752 8968
rect 46296 8848 46348 8857
rect 48596 8848 48648 8900
rect 51080 8959 51132 8968
rect 51080 8925 51089 8959
rect 51089 8925 51123 8959
rect 51123 8925 51132 8959
rect 51080 8916 51132 8925
rect 42340 8823 42392 8832
rect 42340 8789 42349 8823
rect 42349 8789 42383 8823
rect 42383 8789 42392 8823
rect 42340 8780 42392 8789
rect 46204 8780 46256 8832
rect 46572 8780 46624 8832
rect 46664 8780 46716 8832
rect 49516 8780 49568 8832
rect 52736 8780 52788 8832
rect 52920 8823 52972 8832
rect 52920 8789 52929 8823
rect 52929 8789 52963 8823
rect 52963 8789 52972 8823
rect 52920 8780 52972 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 5816 8576 5868 8628
rect 13728 8576 13780 8628
rect 2228 8551 2280 8560
rect 2228 8517 2262 8551
rect 2262 8517 2280 8551
rect 2228 8508 2280 8517
rect 5908 8508 5960 8560
rect 13544 8508 13596 8560
rect 17040 8576 17092 8628
rect 17868 8576 17920 8628
rect 15568 8508 15620 8560
rect 20076 8576 20128 8628
rect 1860 8440 1912 8492
rect 5724 8440 5776 8492
rect 16856 8440 16908 8492
rect 18144 8440 18196 8492
rect 19248 8440 19300 8492
rect 21180 8508 21232 8560
rect 24400 8508 24452 8560
rect 25044 8576 25096 8628
rect 25964 8576 26016 8628
rect 28632 8576 28684 8628
rect 30472 8576 30524 8628
rect 21272 8440 21324 8492
rect 21732 8440 21784 8492
rect 15016 8372 15068 8424
rect 15292 8415 15344 8424
rect 15292 8381 15301 8415
rect 15301 8381 15335 8415
rect 15335 8381 15344 8415
rect 15292 8372 15344 8381
rect 15752 8372 15804 8424
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 3332 8347 3384 8356
rect 3332 8313 3341 8347
rect 3341 8313 3375 8347
rect 3375 8313 3384 8347
rect 3332 8304 3384 8313
rect 6736 8304 6788 8356
rect 16948 8304 17000 8356
rect 21824 8304 21876 8356
rect 22100 8483 22152 8492
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 22468 8440 22520 8492
rect 24584 8440 24636 8492
rect 24768 8483 24820 8492
rect 24768 8449 24778 8483
rect 24778 8449 24812 8483
rect 24812 8449 24820 8483
rect 24768 8440 24820 8449
rect 25228 8440 25280 8492
rect 27712 8508 27764 8560
rect 28724 8551 28776 8560
rect 28724 8517 28733 8551
rect 28733 8517 28767 8551
rect 28767 8517 28776 8551
rect 28724 8508 28776 8517
rect 28816 8508 28868 8560
rect 33324 8551 33376 8560
rect 30196 8483 30248 8492
rect 22468 8304 22520 8356
rect 26148 8304 26200 8356
rect 30196 8449 30205 8483
rect 30205 8449 30239 8483
rect 30239 8449 30248 8483
rect 30196 8440 30248 8449
rect 30932 8440 30984 8492
rect 33324 8517 33333 8551
rect 33333 8517 33367 8551
rect 33367 8517 33376 8551
rect 33324 8508 33376 8517
rect 33508 8576 33560 8628
rect 33876 8576 33928 8628
rect 39580 8576 39632 8628
rect 41604 8576 41656 8628
rect 41788 8576 41840 8628
rect 41880 8576 41932 8628
rect 42892 8551 42944 8560
rect 42892 8517 42927 8551
rect 42927 8517 42944 8551
rect 44732 8551 44784 8560
rect 42892 8508 42944 8517
rect 44732 8517 44741 8551
rect 44741 8517 44775 8551
rect 44775 8517 44784 8551
rect 44732 8508 44784 8517
rect 45008 8551 45060 8560
rect 45008 8517 45017 8551
rect 45017 8517 45051 8551
rect 45051 8517 45060 8551
rect 45008 8508 45060 8517
rect 45468 8576 45520 8628
rect 48596 8619 48648 8628
rect 48596 8585 48605 8619
rect 48605 8585 48639 8619
rect 48639 8585 48648 8619
rect 48596 8576 48648 8585
rect 49700 8576 49752 8628
rect 51080 8576 51132 8628
rect 46204 8508 46256 8560
rect 32956 8440 33008 8492
rect 33876 8372 33928 8424
rect 35348 8372 35400 8424
rect 36544 8440 36596 8492
rect 38752 8483 38804 8492
rect 38752 8449 38761 8483
rect 38761 8449 38795 8483
rect 38795 8449 38804 8483
rect 38752 8440 38804 8449
rect 36820 8372 36872 8424
rect 37004 8372 37056 8424
rect 39764 8440 39816 8492
rect 41512 8440 41564 8492
rect 42340 8440 42392 8492
rect 42616 8483 42668 8492
rect 42616 8449 42625 8483
rect 42625 8449 42659 8483
rect 42659 8449 42668 8483
rect 42616 8440 42668 8449
rect 42708 8483 42760 8492
rect 42708 8449 42717 8483
rect 42717 8449 42751 8483
rect 42751 8449 42760 8483
rect 44916 8483 44968 8492
rect 42708 8440 42760 8449
rect 28540 8304 28592 8356
rect 30380 8304 30432 8356
rect 32312 8347 32364 8356
rect 32312 8313 32321 8347
rect 32321 8313 32355 8347
rect 32355 8313 32364 8347
rect 36360 8347 36412 8356
rect 32312 8304 32364 8313
rect 8944 8236 8996 8288
rect 9404 8236 9456 8288
rect 21364 8236 21416 8288
rect 27620 8236 27672 8288
rect 27896 8236 27948 8288
rect 28724 8236 28776 8288
rect 29000 8236 29052 8288
rect 33140 8236 33192 8288
rect 36360 8313 36369 8347
rect 36369 8313 36403 8347
rect 36403 8313 36412 8347
rect 36360 8304 36412 8313
rect 37924 8347 37976 8356
rect 37924 8313 37933 8347
rect 37933 8313 37967 8347
rect 37967 8313 37976 8347
rect 37924 8304 37976 8313
rect 38568 8304 38620 8356
rect 39120 8372 39172 8424
rect 44916 8449 44925 8483
rect 44925 8449 44959 8483
rect 44959 8449 44968 8483
rect 44916 8440 44968 8449
rect 48780 8483 48832 8492
rect 41696 8304 41748 8356
rect 44548 8372 44600 8424
rect 48228 8372 48280 8424
rect 48780 8449 48789 8483
rect 48789 8449 48823 8483
rect 48823 8449 48832 8483
rect 48780 8440 48832 8449
rect 49608 8440 49660 8492
rect 52460 8440 52512 8492
rect 52920 8440 52972 8492
rect 49700 8372 49752 8424
rect 54852 8372 54904 8424
rect 33692 8236 33744 8288
rect 35440 8279 35492 8288
rect 35440 8245 35449 8279
rect 35449 8245 35483 8279
rect 35483 8245 35492 8279
rect 35440 8236 35492 8245
rect 35808 8236 35860 8288
rect 37004 8236 37056 8288
rect 37188 8236 37240 8288
rect 41512 8236 41564 8288
rect 49424 8236 49476 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 6000 8075 6052 8084
rect 2688 7964 2740 8016
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 6000 8041 6009 8075
rect 6009 8041 6043 8075
rect 6043 8041 6052 8075
rect 6000 8032 6052 8041
rect 10048 8032 10100 8084
rect 13084 8075 13136 8084
rect 13084 8041 13093 8075
rect 13093 8041 13127 8075
rect 13127 8041 13136 8075
rect 13084 8032 13136 8041
rect 14188 8032 14240 8084
rect 17500 8032 17552 8084
rect 19248 8075 19300 8084
rect 19248 8041 19257 8075
rect 19257 8041 19291 8075
rect 19291 8041 19300 8075
rect 19248 8032 19300 8041
rect 23112 8032 23164 8084
rect 24676 8075 24728 8084
rect 24676 8041 24685 8075
rect 24685 8041 24719 8075
rect 24719 8041 24728 8075
rect 24676 8032 24728 8041
rect 4620 7939 4672 7948
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 6276 7828 6328 7880
rect 2872 7735 2924 7744
rect 2872 7701 2881 7735
rect 2881 7701 2915 7735
rect 2915 7701 2924 7735
rect 2872 7692 2924 7701
rect 5264 7760 5316 7812
rect 7748 7896 7800 7948
rect 8484 7896 8536 7948
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 8852 7828 8904 7880
rect 13912 7964 13964 8016
rect 17592 7964 17644 8016
rect 24308 7964 24360 8016
rect 10968 7896 11020 7948
rect 15936 7896 15988 7948
rect 19248 7896 19300 7948
rect 21088 7896 21140 7948
rect 25136 7896 25188 7948
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 12256 7828 12308 7880
rect 15292 7828 15344 7880
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 15568 7871 15620 7880
rect 15568 7837 15577 7871
rect 15577 7837 15611 7871
rect 15611 7837 15620 7871
rect 15568 7828 15620 7837
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 19432 7871 19484 7880
rect 15752 7828 15804 7837
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 19984 7828 20036 7880
rect 25228 7828 25280 7880
rect 27620 8032 27672 8084
rect 25596 7896 25648 7948
rect 27896 8032 27948 8084
rect 32588 8032 32640 8084
rect 46480 8075 46532 8084
rect 33324 7964 33376 8016
rect 34796 7964 34848 8016
rect 35532 7964 35584 8016
rect 38384 7964 38436 8016
rect 38752 8007 38804 8016
rect 38752 7973 38761 8007
rect 38761 7973 38795 8007
rect 38795 7973 38804 8007
rect 38752 7964 38804 7973
rect 42432 7964 42484 8016
rect 46480 8041 46489 8075
rect 46489 8041 46523 8075
rect 46523 8041 46532 8075
rect 46480 8032 46532 8041
rect 49700 8032 49752 8084
rect 49424 7964 49476 8016
rect 9680 7760 9732 7812
rect 12624 7760 12676 7812
rect 14096 7803 14148 7812
rect 14096 7769 14105 7803
rect 14105 7769 14139 7803
rect 14139 7769 14148 7803
rect 14096 7760 14148 7769
rect 14280 7803 14332 7812
rect 14280 7769 14305 7803
rect 14305 7769 14332 7803
rect 14280 7760 14332 7769
rect 20076 7760 20128 7812
rect 24492 7803 24544 7812
rect 24492 7769 24501 7803
rect 24501 7769 24535 7803
rect 24535 7769 24544 7803
rect 24492 7760 24544 7769
rect 5540 7692 5592 7744
rect 8208 7735 8260 7744
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 8300 7692 8352 7744
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 10232 7692 10284 7744
rect 12440 7692 12492 7744
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 14464 7692 14516 7701
rect 14556 7692 14608 7744
rect 16212 7692 16264 7744
rect 19340 7692 19392 7744
rect 20536 7692 20588 7744
rect 21640 7692 21692 7744
rect 24124 7692 24176 7744
rect 24860 7735 24912 7744
rect 24860 7701 24869 7735
rect 24869 7701 24903 7735
rect 24903 7701 24912 7735
rect 24860 7692 24912 7701
rect 25412 7692 25464 7744
rect 26240 7803 26292 7812
rect 26240 7769 26249 7803
rect 26249 7769 26283 7803
rect 26283 7769 26292 7803
rect 26240 7760 26292 7769
rect 27436 7760 27488 7812
rect 27896 7828 27948 7880
rect 28172 7871 28224 7880
rect 28172 7837 28181 7871
rect 28181 7837 28215 7871
rect 28215 7837 28224 7871
rect 28172 7828 28224 7837
rect 27712 7760 27764 7812
rect 25688 7735 25740 7744
rect 25688 7701 25697 7735
rect 25697 7701 25731 7735
rect 25731 7701 25740 7735
rect 25688 7692 25740 7701
rect 26332 7735 26384 7744
rect 26332 7701 26341 7735
rect 26341 7701 26375 7735
rect 26375 7701 26384 7735
rect 26332 7692 26384 7701
rect 27988 7692 28040 7744
rect 28264 7692 28316 7744
rect 28908 7692 28960 7744
rect 30104 7692 30156 7744
rect 32680 7828 32732 7880
rect 37740 7896 37792 7948
rect 35072 7828 35124 7880
rect 35440 7828 35492 7880
rect 39120 7896 39172 7948
rect 40040 7896 40092 7948
rect 41236 7939 41288 7948
rect 41236 7905 41245 7939
rect 41245 7905 41279 7939
rect 41279 7905 41288 7939
rect 41236 7896 41288 7905
rect 42892 7896 42944 7948
rect 45468 7896 45520 7948
rect 38016 7871 38068 7880
rect 38016 7837 38025 7871
rect 38025 7837 38059 7871
rect 38059 7837 38068 7871
rect 38016 7828 38068 7837
rect 38568 7871 38620 7880
rect 38568 7837 38577 7871
rect 38577 7837 38611 7871
rect 38611 7837 38620 7871
rect 38568 7828 38620 7837
rect 41512 7871 41564 7880
rect 41512 7837 41546 7871
rect 41546 7837 41564 7871
rect 41512 7828 41564 7837
rect 42340 7828 42392 7880
rect 44180 7828 44232 7880
rect 44272 7828 44324 7880
rect 52736 7871 52788 7880
rect 52736 7837 52745 7871
rect 52745 7837 52779 7871
rect 52779 7837 52788 7871
rect 52736 7828 52788 7837
rect 53012 7871 53064 7880
rect 53012 7837 53021 7871
rect 53021 7837 53055 7871
rect 53055 7837 53064 7871
rect 53012 7828 53064 7837
rect 32128 7760 32180 7812
rect 31852 7692 31904 7744
rect 32956 7760 33008 7812
rect 34796 7760 34848 7812
rect 32588 7692 32640 7744
rect 35256 7692 35308 7744
rect 35532 7692 35584 7744
rect 37188 7692 37240 7744
rect 37280 7692 37332 7744
rect 38108 7760 38160 7812
rect 45928 7760 45980 7812
rect 46020 7760 46072 7812
rect 42524 7692 42576 7744
rect 52552 7735 52604 7744
rect 52552 7701 52561 7735
rect 52561 7701 52595 7735
rect 52595 7701 52604 7735
rect 52552 7692 52604 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 2044 7488 2096 7540
rect 5264 7531 5316 7540
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 12624 7531 12676 7540
rect 4896 7420 4948 7472
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 6000 7420 6052 7472
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 7748 7395 7800 7404
rect 5724 7352 5776 7361
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 8208 7420 8260 7472
rect 12256 7420 12308 7472
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 13084 7488 13136 7540
rect 14096 7488 14148 7540
rect 14556 7420 14608 7472
rect 15476 7488 15528 7540
rect 22836 7488 22888 7540
rect 19248 7463 19300 7472
rect 19248 7429 19257 7463
rect 19257 7429 19291 7463
rect 19291 7429 19300 7463
rect 19248 7420 19300 7429
rect 2688 7327 2740 7336
rect 2688 7293 2697 7327
rect 2697 7293 2731 7327
rect 2731 7293 2740 7327
rect 2688 7284 2740 7293
rect 5540 7284 5592 7336
rect 6460 7284 6512 7336
rect 9220 7284 9272 7336
rect 9496 7284 9548 7336
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 10416 7352 10468 7404
rect 12440 7284 12492 7336
rect 9588 7216 9640 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 2872 7148 2924 7200
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 13636 7352 13688 7404
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 19156 7352 19208 7404
rect 14464 7284 14516 7336
rect 15200 7284 15252 7336
rect 16672 7284 16724 7336
rect 16304 7216 16356 7268
rect 17408 7284 17460 7336
rect 17040 7216 17092 7268
rect 22376 7352 22428 7404
rect 24860 7488 24912 7540
rect 25136 7531 25188 7540
rect 25136 7497 25145 7531
rect 25145 7497 25179 7531
rect 25179 7497 25188 7531
rect 25136 7488 25188 7497
rect 25228 7488 25280 7540
rect 26240 7488 26292 7540
rect 28172 7488 28224 7540
rect 28816 7488 28868 7540
rect 30196 7488 30248 7540
rect 32128 7531 32180 7540
rect 32128 7497 32137 7531
rect 32137 7497 32171 7531
rect 32171 7497 32180 7531
rect 32128 7488 32180 7497
rect 33876 7488 33928 7540
rect 34336 7488 34388 7540
rect 23388 7420 23440 7472
rect 24124 7463 24176 7472
rect 24124 7429 24133 7463
rect 24133 7429 24167 7463
rect 24167 7429 24176 7463
rect 24124 7420 24176 7429
rect 25412 7420 25464 7472
rect 25504 7420 25556 7472
rect 26516 7420 26568 7472
rect 27988 7463 28040 7472
rect 23204 7395 23256 7404
rect 23204 7361 23213 7395
rect 23213 7361 23247 7395
rect 23247 7361 23256 7395
rect 23204 7352 23256 7361
rect 25228 7352 25280 7404
rect 25596 7352 25648 7404
rect 27988 7429 27997 7463
rect 27997 7429 28031 7463
rect 28031 7429 28040 7463
rect 27988 7420 28040 7429
rect 28448 7420 28500 7472
rect 28908 7463 28960 7472
rect 28908 7429 28933 7463
rect 28933 7429 28960 7463
rect 30932 7463 30984 7472
rect 28908 7420 28960 7429
rect 19432 7284 19484 7336
rect 20536 7284 20588 7336
rect 29920 7352 29972 7404
rect 30932 7429 30941 7463
rect 30941 7429 30975 7463
rect 30975 7429 30984 7463
rect 30932 7420 30984 7429
rect 30472 7352 30524 7404
rect 31116 7395 31168 7404
rect 31116 7361 31125 7395
rect 31125 7361 31159 7395
rect 31159 7361 31168 7395
rect 31116 7352 31168 7361
rect 19984 7216 20036 7268
rect 20168 7216 20220 7268
rect 21272 7216 21324 7268
rect 19340 7148 19392 7200
rect 20260 7148 20312 7200
rect 22468 7148 22520 7200
rect 22744 7191 22796 7200
rect 22744 7157 22753 7191
rect 22753 7157 22787 7191
rect 22787 7157 22796 7191
rect 22744 7148 22796 7157
rect 24400 7216 24452 7268
rect 27712 7284 27764 7336
rect 27804 7284 27856 7336
rect 34888 7395 34940 7404
rect 34888 7361 34897 7395
rect 34897 7361 34931 7395
rect 34931 7361 34940 7395
rect 34888 7352 34940 7361
rect 35072 7395 35124 7404
rect 35072 7361 35081 7395
rect 35081 7361 35115 7395
rect 35115 7361 35124 7395
rect 35072 7352 35124 7361
rect 36912 7420 36964 7472
rect 37096 7488 37148 7540
rect 42340 7488 42392 7540
rect 41972 7420 42024 7472
rect 35256 7395 35308 7404
rect 35256 7361 35265 7395
rect 35265 7361 35299 7395
rect 35299 7361 35308 7395
rect 35256 7352 35308 7361
rect 36176 7352 36228 7404
rect 37464 7352 37516 7404
rect 38384 7352 38436 7404
rect 42524 7420 42576 7472
rect 42616 7395 42668 7404
rect 42616 7361 42625 7395
rect 42625 7361 42659 7395
rect 42659 7361 42668 7395
rect 42616 7352 42668 7361
rect 42708 7395 42760 7404
rect 42708 7361 42717 7395
rect 42717 7361 42751 7395
rect 42751 7361 42760 7395
rect 42708 7352 42760 7361
rect 42892 7395 42944 7404
rect 42892 7361 42927 7395
rect 42927 7361 42944 7395
rect 45928 7488 45980 7540
rect 54852 7531 54904 7540
rect 46204 7463 46256 7472
rect 46204 7429 46213 7463
rect 46213 7429 46247 7463
rect 46247 7429 46256 7463
rect 46204 7420 46256 7429
rect 42892 7352 42944 7361
rect 44548 7395 44600 7404
rect 32588 7327 32640 7336
rect 32588 7293 32597 7327
rect 32597 7293 32631 7327
rect 32631 7293 32640 7327
rect 32588 7284 32640 7293
rect 33140 7284 33192 7336
rect 37740 7327 37792 7336
rect 24492 7191 24544 7200
rect 24492 7157 24501 7191
rect 24501 7157 24535 7191
rect 24535 7157 24544 7191
rect 24492 7148 24544 7157
rect 24676 7148 24728 7200
rect 26240 7216 26292 7268
rect 29920 7216 29972 7268
rect 30380 7216 30432 7268
rect 25412 7148 25464 7200
rect 27804 7148 27856 7200
rect 27896 7148 27948 7200
rect 28172 7191 28224 7200
rect 28172 7157 28181 7191
rect 28181 7157 28215 7191
rect 28215 7157 28224 7191
rect 28172 7148 28224 7157
rect 28724 7148 28776 7200
rect 29092 7191 29144 7200
rect 29092 7157 29101 7191
rect 29101 7157 29135 7191
rect 29135 7157 29144 7191
rect 29092 7148 29144 7157
rect 29184 7148 29236 7200
rect 37096 7216 37148 7268
rect 35624 7191 35676 7200
rect 35624 7157 35633 7191
rect 35633 7157 35667 7191
rect 35667 7157 35676 7191
rect 35624 7148 35676 7157
rect 37740 7293 37749 7327
rect 37749 7293 37783 7327
rect 37783 7293 37792 7327
rect 37740 7284 37792 7293
rect 42432 7284 42484 7336
rect 44548 7361 44557 7395
rect 44557 7361 44591 7395
rect 44591 7361 44600 7395
rect 44548 7352 44600 7361
rect 44640 7395 44692 7404
rect 44640 7361 44649 7395
rect 44649 7361 44683 7395
rect 44683 7361 44692 7395
rect 44640 7352 44692 7361
rect 45928 7352 45980 7404
rect 46020 7395 46072 7404
rect 46020 7361 46029 7395
rect 46029 7361 46063 7395
rect 46063 7361 46072 7395
rect 54852 7497 54861 7531
rect 54861 7497 54895 7531
rect 54895 7497 54904 7531
rect 54852 7488 54904 7497
rect 52552 7420 52604 7472
rect 46020 7352 46072 7361
rect 48780 7352 48832 7404
rect 49332 7395 49384 7404
rect 49332 7361 49341 7395
rect 49341 7361 49375 7395
rect 49375 7361 49384 7395
rect 49332 7352 49384 7361
rect 49424 7352 49476 7404
rect 49608 7327 49660 7336
rect 49608 7293 49617 7327
rect 49617 7293 49651 7327
rect 49651 7293 49660 7327
rect 49608 7284 49660 7293
rect 49884 7284 49936 7336
rect 51540 7352 51592 7404
rect 53104 7352 53156 7404
rect 39120 7191 39172 7200
rect 39120 7157 39129 7191
rect 39129 7157 39163 7191
rect 39163 7157 39172 7191
rect 39120 7148 39172 7157
rect 43076 7148 43128 7200
rect 45284 7148 45336 7200
rect 47216 7148 47268 7200
rect 51540 7148 51592 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6944 1636 6996
rect 14188 6944 14240 6996
rect 17132 6944 17184 6996
rect 5724 6808 5776 6860
rect 15200 6876 15252 6928
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 2872 6783 2924 6792
rect 2872 6749 2881 6783
rect 2881 6749 2915 6783
rect 2915 6749 2924 6783
rect 2872 6740 2924 6749
rect 6276 6783 6328 6792
rect 3516 6672 3568 6724
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 11888 6808 11940 6860
rect 8116 6740 8168 6792
rect 9588 6740 9640 6792
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 14464 6740 14516 6792
rect 15108 6808 15160 6860
rect 15660 6851 15712 6860
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 19708 6944 19760 6996
rect 23388 6944 23440 6996
rect 23756 6944 23808 6996
rect 27804 6944 27856 6996
rect 27896 6944 27948 6996
rect 19432 6876 19484 6928
rect 21732 6876 21784 6928
rect 23204 6876 23256 6928
rect 34520 6944 34572 6996
rect 34796 6944 34848 6996
rect 35808 6944 35860 6996
rect 37464 6987 37516 6996
rect 37464 6953 37473 6987
rect 37473 6953 37507 6987
rect 37507 6953 37516 6987
rect 37464 6944 37516 6953
rect 37740 6944 37792 6996
rect 40040 6944 40092 6996
rect 30656 6919 30708 6928
rect 17408 6851 17460 6860
rect 17408 6817 17417 6851
rect 17417 6817 17451 6851
rect 17451 6817 17460 6851
rect 17408 6808 17460 6817
rect 17500 6808 17552 6860
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 17316 6783 17368 6792
rect 17316 6749 17325 6783
rect 17325 6749 17359 6783
rect 17359 6749 17368 6783
rect 19432 6783 19484 6792
rect 17316 6740 17368 6749
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 19708 6783 19760 6792
rect 19708 6749 19717 6783
rect 19717 6749 19751 6783
rect 19751 6749 19760 6783
rect 19708 6740 19760 6749
rect 2596 6604 2648 6656
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 9128 6672 9180 6724
rect 19156 6672 19208 6724
rect 7472 6604 7524 6656
rect 10232 6604 10284 6656
rect 11152 6604 11204 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 14464 6647 14516 6656
rect 14464 6613 14473 6647
rect 14473 6613 14507 6647
rect 14507 6613 14516 6647
rect 14464 6604 14516 6613
rect 15384 6604 15436 6656
rect 19248 6647 19300 6656
rect 19248 6613 19257 6647
rect 19257 6613 19291 6647
rect 19291 6613 19300 6647
rect 19248 6604 19300 6613
rect 19340 6604 19392 6656
rect 25228 6808 25280 6860
rect 26148 6808 26200 6860
rect 26332 6808 26384 6860
rect 30656 6885 30665 6919
rect 30665 6885 30699 6919
rect 30699 6885 30708 6919
rect 30656 6876 30708 6885
rect 31116 6876 31168 6928
rect 30196 6808 30248 6860
rect 20628 6740 20680 6792
rect 22744 6740 22796 6792
rect 32496 6808 32548 6860
rect 33416 6808 33468 6860
rect 37188 6808 37240 6860
rect 25596 6672 25648 6724
rect 32312 6783 32364 6792
rect 32312 6749 32321 6783
rect 32321 6749 32355 6783
rect 32355 6749 32364 6783
rect 32312 6740 32364 6749
rect 22836 6604 22888 6656
rect 26424 6604 26476 6656
rect 27528 6604 27580 6656
rect 27988 6647 28040 6656
rect 27988 6613 28013 6647
rect 28013 6613 28040 6647
rect 27988 6604 28040 6613
rect 30840 6672 30892 6724
rect 33324 6740 33376 6792
rect 34704 6740 34756 6792
rect 35624 6740 35676 6792
rect 36544 6740 36596 6792
rect 36912 6783 36964 6792
rect 36912 6749 36921 6783
rect 36921 6749 36955 6783
rect 36955 6749 36964 6783
rect 36912 6740 36964 6749
rect 37372 6808 37424 6860
rect 37464 6808 37516 6860
rect 44180 6808 44232 6860
rect 45376 6944 45428 6996
rect 51540 6808 51592 6860
rect 32496 6715 32548 6724
rect 32496 6681 32505 6715
rect 32505 6681 32539 6715
rect 32539 6681 32548 6715
rect 32496 6672 32548 6681
rect 32864 6647 32916 6656
rect 32864 6613 32873 6647
rect 32873 6613 32907 6647
rect 32907 6613 32916 6647
rect 32864 6604 32916 6613
rect 36176 6647 36228 6656
rect 36176 6613 36185 6647
rect 36185 6613 36219 6647
rect 36219 6613 36228 6647
rect 36176 6604 36228 6613
rect 36820 6672 36872 6724
rect 46940 6740 46992 6792
rect 47124 6783 47176 6792
rect 47124 6749 47133 6783
rect 47133 6749 47167 6783
rect 47167 6749 47176 6783
rect 47124 6740 47176 6749
rect 47216 6740 47268 6792
rect 48228 6740 48280 6792
rect 48872 6740 48924 6792
rect 49332 6783 49384 6792
rect 49332 6749 49341 6783
rect 49341 6749 49375 6783
rect 49375 6749 49384 6783
rect 49332 6740 49384 6749
rect 40684 6672 40736 6724
rect 45284 6715 45336 6724
rect 45284 6681 45318 6715
rect 45318 6681 45336 6715
rect 45284 6672 45336 6681
rect 45376 6672 45428 6724
rect 50160 6740 50212 6792
rect 52736 6808 52788 6860
rect 50068 6672 50120 6724
rect 52920 6783 52972 6792
rect 52920 6749 52929 6783
rect 52929 6749 52963 6783
rect 52963 6749 52972 6783
rect 52920 6740 52972 6749
rect 37372 6604 37424 6656
rect 39120 6604 39172 6656
rect 41420 6647 41472 6656
rect 41420 6613 41429 6647
rect 41429 6613 41463 6647
rect 41463 6613 41472 6647
rect 41420 6604 41472 6613
rect 45928 6604 45980 6656
rect 48412 6604 48464 6656
rect 49700 6604 49752 6656
rect 53288 6604 53340 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 3332 6400 3384 6452
rect 3516 6332 3568 6384
rect 15660 6400 15712 6452
rect 17316 6400 17368 6452
rect 23388 6400 23440 6452
rect 24584 6400 24636 6452
rect 32680 6400 32732 6452
rect 33600 6400 33652 6452
rect 36820 6400 36872 6452
rect 38292 6400 38344 6452
rect 44548 6443 44600 6452
rect 5908 6332 5960 6384
rect 14096 6332 14148 6384
rect 2688 6239 2740 6248
rect 2688 6205 2697 6239
rect 2697 6205 2731 6239
rect 2731 6205 2740 6239
rect 2688 6196 2740 6205
rect 5724 6264 5776 6316
rect 10416 6264 10468 6316
rect 10968 6264 11020 6316
rect 13820 6264 13872 6316
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 15752 6264 15804 6316
rect 15936 6264 15988 6316
rect 19248 6332 19300 6384
rect 22100 6332 22152 6384
rect 22560 6332 22612 6384
rect 28356 6332 28408 6384
rect 29460 6375 29512 6384
rect 29460 6341 29469 6375
rect 29469 6341 29503 6375
rect 29503 6341 29512 6375
rect 29460 6332 29512 6341
rect 31300 6332 31352 6384
rect 32864 6332 32916 6384
rect 44548 6409 44557 6443
rect 44557 6409 44591 6443
rect 44591 6409 44600 6443
rect 44548 6400 44600 6409
rect 46204 6400 46256 6452
rect 46848 6400 46900 6452
rect 44180 6375 44232 6384
rect 18144 6264 18196 6316
rect 20628 6264 20680 6316
rect 21364 6264 21416 6316
rect 22284 6307 22336 6316
rect 22284 6273 22293 6307
rect 22293 6273 22327 6307
rect 22327 6273 22336 6307
rect 22284 6264 22336 6273
rect 25688 6264 25740 6316
rect 36268 6307 36320 6316
rect 36268 6273 36277 6307
rect 36277 6273 36311 6307
rect 36311 6273 36320 6307
rect 36268 6264 36320 6273
rect 5356 6196 5408 6248
rect 15568 6239 15620 6248
rect 15568 6205 15577 6239
rect 15577 6205 15611 6239
rect 15611 6205 15620 6239
rect 15568 6196 15620 6205
rect 16856 6239 16908 6248
rect 16856 6205 16865 6239
rect 16865 6205 16899 6239
rect 16899 6205 16908 6239
rect 16856 6196 16908 6205
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 5448 6128 5500 6180
rect 8852 6128 8904 6180
rect 9220 6128 9272 6180
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 3608 6060 3660 6112
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 6276 6060 6328 6112
rect 8944 6060 8996 6112
rect 9128 6060 9180 6112
rect 14464 6103 14516 6112
rect 14464 6069 14473 6103
rect 14473 6069 14507 6103
rect 14507 6069 14516 6103
rect 14464 6060 14516 6069
rect 19156 6060 19208 6112
rect 23848 6128 23900 6180
rect 30840 6196 30892 6248
rect 31852 6196 31904 6248
rect 36360 6196 36412 6248
rect 40040 6264 40092 6316
rect 41420 6264 41472 6316
rect 43076 6307 43128 6316
rect 43076 6273 43085 6307
rect 43085 6273 43119 6307
rect 43119 6273 43128 6307
rect 43076 6264 43128 6273
rect 36636 6196 36688 6248
rect 28172 6128 28224 6180
rect 22284 6060 22336 6112
rect 24952 6060 25004 6112
rect 25780 6060 25832 6112
rect 28724 6060 28776 6112
rect 28908 6060 28960 6112
rect 29828 6103 29880 6112
rect 29828 6069 29837 6103
rect 29837 6069 29871 6103
rect 29871 6069 29880 6103
rect 29828 6060 29880 6069
rect 39672 6128 39724 6180
rect 40592 6196 40644 6248
rect 43168 6239 43220 6248
rect 43168 6205 43177 6239
rect 43177 6205 43211 6239
rect 43211 6205 43220 6239
rect 43168 6196 43220 6205
rect 44180 6341 44189 6375
rect 44189 6341 44223 6375
rect 44223 6341 44232 6375
rect 44180 6332 44232 6341
rect 45928 6332 45980 6384
rect 43996 6307 44048 6316
rect 43996 6273 44005 6307
rect 44005 6273 44039 6307
rect 44039 6273 44048 6307
rect 43996 6264 44048 6273
rect 44364 6307 44416 6316
rect 44364 6273 44373 6307
rect 44373 6273 44407 6307
rect 44407 6273 44416 6307
rect 44364 6264 44416 6273
rect 48872 6375 48924 6384
rect 46296 6264 46348 6316
rect 48872 6341 48881 6375
rect 48881 6341 48915 6375
rect 48915 6341 48924 6375
rect 48872 6332 48924 6341
rect 49608 6400 49660 6452
rect 50160 6443 50212 6452
rect 50160 6409 50169 6443
rect 50169 6409 50203 6443
rect 50203 6409 50212 6443
rect 50160 6400 50212 6409
rect 53012 6400 53064 6452
rect 50988 6332 51040 6384
rect 52184 6332 52236 6384
rect 48412 6264 48464 6316
rect 48780 6307 48832 6316
rect 48780 6273 48789 6307
rect 48789 6273 48823 6307
rect 48823 6273 48832 6307
rect 48780 6264 48832 6273
rect 49424 6264 49476 6316
rect 49608 6307 49660 6316
rect 49608 6273 49617 6307
rect 49617 6273 49651 6307
rect 49651 6273 49660 6307
rect 49608 6264 49660 6273
rect 49792 6264 49844 6316
rect 52736 6307 52788 6316
rect 41880 6128 41932 6180
rect 42616 6128 42668 6180
rect 42892 6128 42944 6180
rect 46480 6196 46532 6248
rect 48596 6128 48648 6180
rect 49516 6128 49568 6180
rect 52736 6273 52745 6307
rect 52745 6273 52779 6307
rect 52779 6273 52788 6307
rect 52736 6264 52788 6273
rect 54852 6332 54904 6384
rect 52368 6128 52420 6180
rect 33140 6060 33192 6112
rect 37004 6060 37056 6112
rect 39948 6060 40000 6112
rect 43812 6060 43864 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 5448 5899 5500 5908
rect 5448 5865 5457 5899
rect 5457 5865 5491 5899
rect 5491 5865 5500 5899
rect 5448 5856 5500 5865
rect 8668 5856 8720 5908
rect 9128 5856 9180 5908
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 5540 5720 5592 5772
rect 11980 5856 12032 5908
rect 12348 5856 12400 5908
rect 16856 5856 16908 5908
rect 21272 5856 21324 5908
rect 27436 5856 27488 5908
rect 27988 5856 28040 5908
rect 28540 5856 28592 5908
rect 28908 5856 28960 5908
rect 31576 5856 31628 5908
rect 15108 5788 15160 5840
rect 19340 5788 19392 5840
rect 22192 5788 22244 5840
rect 14464 5720 14516 5772
rect 17408 5720 17460 5772
rect 22008 5720 22060 5772
rect 2596 5652 2648 5704
rect 2044 5584 2096 5636
rect 4160 5652 4212 5704
rect 4804 5652 4856 5704
rect 8944 5695 8996 5704
rect 8944 5661 8953 5695
rect 8953 5661 8987 5695
rect 8987 5661 8996 5695
rect 8944 5652 8996 5661
rect 9772 5652 9824 5704
rect 10968 5652 11020 5704
rect 11888 5652 11940 5704
rect 15200 5652 15252 5704
rect 3332 5584 3384 5636
rect 8116 5584 8168 5636
rect 11152 5627 11204 5636
rect 11152 5593 11186 5627
rect 11186 5593 11204 5627
rect 11152 5584 11204 5593
rect 4896 5516 4948 5568
rect 8576 5516 8628 5568
rect 9680 5559 9732 5568
rect 9680 5525 9689 5559
rect 9689 5525 9723 5559
rect 9723 5525 9732 5559
rect 9680 5516 9732 5525
rect 17132 5652 17184 5704
rect 22100 5695 22152 5704
rect 22100 5661 22109 5695
rect 22109 5661 22143 5695
rect 22143 5661 22152 5695
rect 22100 5652 22152 5661
rect 23296 5652 23348 5704
rect 26332 5788 26384 5840
rect 26976 5788 27028 5840
rect 38752 5856 38804 5908
rect 25872 5720 25924 5772
rect 26792 5763 26844 5772
rect 26792 5729 26801 5763
rect 26801 5729 26835 5763
rect 26835 5729 26844 5763
rect 26792 5720 26844 5729
rect 26884 5720 26936 5772
rect 25688 5695 25740 5704
rect 25688 5661 25697 5695
rect 25697 5661 25731 5695
rect 25731 5661 25740 5695
rect 26332 5695 26384 5704
rect 25688 5652 25740 5661
rect 26332 5661 26341 5695
rect 26341 5661 26375 5695
rect 26375 5661 26384 5695
rect 26332 5652 26384 5661
rect 27436 5695 27488 5704
rect 21456 5627 21508 5636
rect 21456 5593 21465 5627
rect 21465 5593 21499 5627
rect 21499 5593 21508 5627
rect 21456 5584 21508 5593
rect 25320 5627 25372 5636
rect 25320 5593 25329 5627
rect 25329 5593 25363 5627
rect 25363 5593 25372 5627
rect 25320 5584 25372 5593
rect 26424 5630 26476 5682
rect 27436 5661 27445 5695
rect 27445 5661 27479 5695
rect 27479 5661 27488 5695
rect 27436 5652 27488 5661
rect 33048 5788 33100 5840
rect 38292 5831 38344 5840
rect 38292 5797 38301 5831
rect 38301 5797 38335 5831
rect 38335 5797 38344 5831
rect 38292 5788 38344 5797
rect 27896 5695 27948 5704
rect 27896 5661 27905 5695
rect 27905 5661 27939 5695
rect 27939 5661 27948 5695
rect 27896 5652 27948 5661
rect 28540 5695 28592 5704
rect 28540 5661 28549 5695
rect 28549 5661 28583 5695
rect 28583 5661 28592 5695
rect 28540 5652 28592 5661
rect 28724 5695 28776 5704
rect 28724 5661 28733 5695
rect 28733 5661 28767 5695
rect 28767 5661 28776 5695
rect 28724 5652 28776 5661
rect 33416 5720 33468 5772
rect 35808 5720 35860 5772
rect 37464 5720 37516 5772
rect 39856 5763 39908 5772
rect 39856 5729 39865 5763
rect 39865 5729 39899 5763
rect 39899 5729 39908 5763
rect 39856 5720 39908 5729
rect 41328 5720 41380 5772
rect 52920 5856 52972 5908
rect 42524 5788 42576 5840
rect 50068 5788 50120 5840
rect 25044 5559 25096 5568
rect 25044 5525 25053 5559
rect 25053 5525 25087 5559
rect 25087 5525 25096 5559
rect 25044 5516 25096 5525
rect 26148 5559 26200 5568
rect 26148 5525 26157 5559
rect 26157 5525 26191 5559
rect 26191 5525 26200 5559
rect 26148 5516 26200 5525
rect 26516 5627 26568 5636
rect 26516 5593 26525 5627
rect 26525 5593 26559 5627
rect 26559 5593 26568 5627
rect 26516 5584 26568 5593
rect 26976 5584 27028 5636
rect 27528 5627 27580 5636
rect 27528 5593 27537 5627
rect 27537 5593 27571 5627
rect 27571 5593 27580 5627
rect 27528 5584 27580 5593
rect 29460 5652 29512 5704
rect 29552 5627 29604 5636
rect 29552 5593 29561 5627
rect 29561 5593 29595 5627
rect 29595 5593 29604 5627
rect 29552 5584 29604 5593
rect 31300 5584 31352 5636
rect 27988 5516 28040 5568
rect 29000 5516 29052 5568
rect 29920 5559 29972 5568
rect 29920 5525 29929 5559
rect 29929 5525 29963 5559
rect 29963 5525 29972 5559
rect 29920 5516 29972 5525
rect 32404 5652 32456 5704
rect 32496 5627 32548 5636
rect 32496 5593 32505 5627
rect 32505 5593 32539 5627
rect 32539 5593 32548 5627
rect 32496 5584 32548 5593
rect 33600 5652 33652 5704
rect 36268 5652 36320 5704
rect 36452 5695 36504 5704
rect 36452 5661 36461 5695
rect 36461 5661 36495 5695
rect 36495 5661 36504 5695
rect 36452 5652 36504 5661
rect 38568 5652 38620 5704
rect 39948 5652 40000 5704
rect 41880 5695 41932 5704
rect 41880 5661 41889 5695
rect 41889 5661 41923 5695
rect 41923 5661 41932 5695
rect 41880 5652 41932 5661
rect 41972 5695 42024 5704
rect 41972 5661 41981 5695
rect 41981 5661 42015 5695
rect 42015 5661 42024 5695
rect 41972 5652 42024 5661
rect 42892 5652 42944 5704
rect 46020 5652 46072 5704
rect 52460 5720 52512 5772
rect 52184 5695 52236 5704
rect 52184 5661 52193 5695
rect 52193 5661 52227 5695
rect 52227 5661 52236 5695
rect 52184 5652 52236 5661
rect 52368 5695 52420 5704
rect 52368 5661 52377 5695
rect 52377 5661 52411 5695
rect 52411 5661 52420 5695
rect 52368 5652 52420 5661
rect 53104 5652 53156 5704
rect 53288 5695 53340 5704
rect 53288 5661 53322 5695
rect 53322 5661 53340 5695
rect 53288 5652 53340 5661
rect 32680 5516 32732 5568
rect 33324 5516 33376 5568
rect 35716 5516 35768 5568
rect 35900 5559 35952 5568
rect 35900 5525 35909 5559
rect 35909 5525 35943 5559
rect 35943 5525 35952 5559
rect 35900 5516 35952 5525
rect 39856 5516 39908 5568
rect 40316 5516 40368 5568
rect 40408 5516 40460 5568
rect 41328 5516 41380 5568
rect 41696 5559 41748 5568
rect 41696 5525 41705 5559
rect 41705 5525 41739 5559
rect 41739 5525 41748 5559
rect 41696 5516 41748 5525
rect 41972 5516 42024 5568
rect 42708 5584 42760 5636
rect 42800 5559 42852 5568
rect 42800 5525 42809 5559
rect 42809 5525 42843 5559
rect 42843 5525 42852 5559
rect 42800 5516 42852 5525
rect 42984 5516 43036 5568
rect 45376 5584 45428 5636
rect 46388 5627 46440 5636
rect 46388 5593 46397 5627
rect 46397 5593 46431 5627
rect 46431 5593 46440 5627
rect 46388 5584 46440 5593
rect 49516 5584 49568 5636
rect 52736 5516 52788 5568
rect 54392 5559 54444 5568
rect 54392 5525 54401 5559
rect 54401 5525 54435 5559
rect 54435 5525 54444 5559
rect 54392 5516 54444 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 1860 5287 1912 5296
rect 1860 5253 1869 5287
rect 1869 5253 1903 5287
rect 1903 5253 1912 5287
rect 1860 5244 1912 5253
rect 5540 5312 5592 5364
rect 8852 5312 8904 5364
rect 11152 5312 11204 5364
rect 14832 5312 14884 5364
rect 19432 5312 19484 5364
rect 22100 5312 22152 5364
rect 25688 5312 25740 5364
rect 32312 5312 32364 5364
rect 32680 5312 32732 5364
rect 32956 5312 33008 5364
rect 33140 5312 33192 5364
rect 35992 5312 36044 5364
rect 38752 5355 38804 5364
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 4160 5176 4212 5228
rect 4804 5176 4856 5228
rect 3792 5108 3844 5160
rect 7288 5176 7340 5228
rect 8484 5244 8536 5296
rect 9680 5176 9732 5228
rect 14832 5219 14884 5228
rect 14832 5185 14841 5219
rect 14841 5185 14875 5219
rect 14875 5185 14884 5219
rect 14832 5176 14884 5185
rect 15016 5219 15068 5228
rect 15016 5185 15025 5219
rect 15025 5185 15059 5219
rect 15059 5185 15068 5219
rect 15016 5176 15068 5185
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 2872 5015 2924 5024
rect 2872 4981 2881 5015
rect 2881 4981 2915 5015
rect 2915 4981 2924 5015
rect 2872 4972 2924 4981
rect 3424 5015 3476 5024
rect 3424 4981 3433 5015
rect 3433 4981 3467 5015
rect 3467 4981 3476 5015
rect 3424 4972 3476 4981
rect 3516 4972 3568 5024
rect 4804 4972 4856 5024
rect 5264 4972 5316 5024
rect 10876 5108 10928 5160
rect 13636 5108 13688 5160
rect 18328 5176 18380 5228
rect 20076 5176 20128 5228
rect 20260 5108 20312 5160
rect 21824 5151 21876 5160
rect 21824 5117 21833 5151
rect 21833 5117 21867 5151
rect 21867 5117 21876 5151
rect 21824 5108 21876 5117
rect 21640 5040 21692 5092
rect 8944 4972 8996 5024
rect 14648 5015 14700 5024
rect 14648 4981 14657 5015
rect 14657 4981 14691 5015
rect 14691 4981 14700 5015
rect 14648 4972 14700 4981
rect 18512 5015 18564 5024
rect 18512 4981 18521 5015
rect 18521 4981 18555 5015
rect 18555 4981 18564 5015
rect 18512 4972 18564 4981
rect 19432 5015 19484 5024
rect 19432 4981 19441 5015
rect 19441 4981 19475 5015
rect 19475 4981 19484 5015
rect 19432 4972 19484 4981
rect 20076 4972 20128 5024
rect 22192 5219 22244 5228
rect 22192 5185 22201 5219
rect 22201 5185 22235 5219
rect 22235 5185 22244 5219
rect 22192 5176 22244 5185
rect 25228 5176 25280 5228
rect 25504 5176 25556 5228
rect 26148 5176 26200 5228
rect 27988 5219 28040 5228
rect 27528 5108 27580 5160
rect 27988 5185 27997 5219
rect 27997 5185 28031 5219
rect 28031 5185 28040 5219
rect 27988 5176 28040 5185
rect 29920 5244 29972 5296
rect 29000 5219 29052 5228
rect 29000 5185 29009 5219
rect 29009 5185 29043 5219
rect 29043 5185 29052 5219
rect 29000 5176 29052 5185
rect 29828 5176 29880 5228
rect 30472 5244 30524 5296
rect 31116 5244 31168 5296
rect 31300 5287 31352 5296
rect 31300 5253 31309 5287
rect 31309 5253 31343 5287
rect 31343 5253 31352 5287
rect 31300 5244 31352 5253
rect 32128 5244 32180 5296
rect 30104 5176 30156 5228
rect 34152 5244 34204 5296
rect 38752 5321 38761 5355
rect 38761 5321 38795 5355
rect 38795 5321 38804 5355
rect 38752 5312 38804 5321
rect 40592 5312 40644 5364
rect 40960 5312 41012 5364
rect 38292 5244 38344 5296
rect 40224 5244 40276 5296
rect 42708 5287 42760 5296
rect 42708 5253 42717 5287
rect 42717 5253 42751 5287
rect 42751 5253 42760 5287
rect 42708 5244 42760 5253
rect 42892 5287 42944 5296
rect 42892 5253 42917 5287
rect 42917 5253 42944 5287
rect 43168 5312 43220 5364
rect 42892 5244 42944 5253
rect 44364 5244 44416 5296
rect 45376 5287 45428 5296
rect 45376 5253 45385 5287
rect 45385 5253 45419 5287
rect 45419 5253 45428 5287
rect 45376 5244 45428 5253
rect 32496 5219 32548 5228
rect 32496 5185 32505 5219
rect 32505 5185 32539 5219
rect 32539 5185 32548 5219
rect 32496 5176 32548 5185
rect 32956 5176 33008 5228
rect 26332 4972 26384 5024
rect 27620 5015 27672 5024
rect 27620 4981 27629 5015
rect 27629 4981 27663 5015
rect 27663 4981 27672 5015
rect 27620 4972 27672 4981
rect 28632 5015 28684 5024
rect 28632 4981 28641 5015
rect 28641 4981 28675 5015
rect 28675 4981 28684 5015
rect 28632 4972 28684 4981
rect 31208 4972 31260 5024
rect 31300 4972 31352 5024
rect 34520 4972 34572 5024
rect 34704 5151 34756 5160
rect 34704 5117 34713 5151
rect 34713 5117 34747 5151
rect 34747 5117 34756 5151
rect 35900 5176 35952 5228
rect 38568 5176 38620 5228
rect 40132 5219 40184 5228
rect 40132 5185 40141 5219
rect 40141 5185 40175 5219
rect 40175 5185 40184 5219
rect 40132 5176 40184 5185
rect 40408 5219 40460 5228
rect 40408 5185 40417 5219
rect 40417 5185 40451 5219
rect 40451 5185 40460 5219
rect 40408 5176 40460 5185
rect 40500 5219 40552 5228
rect 40500 5185 40533 5219
rect 40533 5185 40552 5219
rect 40500 5176 40552 5185
rect 47124 5176 47176 5228
rect 34704 5108 34756 5117
rect 36176 5108 36228 5160
rect 36452 5108 36504 5160
rect 37556 5151 37608 5160
rect 37556 5117 37565 5151
rect 37565 5117 37599 5151
rect 37599 5117 37608 5151
rect 37556 5108 37608 5117
rect 46480 5151 46532 5160
rect 36176 4972 36228 5024
rect 40500 5040 40552 5092
rect 46480 5117 46489 5151
rect 46489 5117 46523 5151
rect 46523 5117 46532 5151
rect 46480 5108 46532 5117
rect 48228 5108 48280 5160
rect 49884 5312 49936 5364
rect 50988 5355 51040 5364
rect 50988 5321 50997 5355
rect 50997 5321 51031 5355
rect 51031 5321 51040 5355
rect 50988 5312 51040 5321
rect 49700 5176 49752 5228
rect 40132 4972 40184 5024
rect 41420 4972 41472 5024
rect 41604 4972 41656 5024
rect 42616 4972 42668 5024
rect 45468 5015 45520 5024
rect 45468 4981 45477 5015
rect 45477 4981 45511 5015
rect 45511 4981 45520 5015
rect 45468 4972 45520 4981
rect 46756 4972 46808 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 7288 4811 7340 4820
rect 1584 4700 1636 4752
rect 3976 4700 4028 4752
rect 7288 4777 7297 4811
rect 7297 4777 7331 4811
rect 7331 4777 7340 4811
rect 7288 4768 7340 4777
rect 10048 4768 10100 4820
rect 15016 4768 15068 4820
rect 20260 4768 20312 4820
rect 21272 4811 21324 4820
rect 8484 4700 8536 4752
rect 21272 4777 21281 4811
rect 21281 4777 21315 4811
rect 21315 4777 21324 4811
rect 21272 4768 21324 4777
rect 22192 4768 22244 4820
rect 24492 4768 24544 4820
rect 25044 4768 25096 4820
rect 2688 4564 2740 4616
rect 2964 4564 3016 4616
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 3148 4496 3200 4548
rect 5356 4496 5408 4548
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 8576 4632 8628 4684
rect 10692 4632 10744 4684
rect 13820 4632 13872 4684
rect 16120 4632 16172 4684
rect 19432 4675 19484 4684
rect 19432 4641 19441 4675
rect 19441 4641 19475 4675
rect 19475 4641 19484 4675
rect 19432 4632 19484 4641
rect 21640 4675 21692 4684
rect 7748 4564 7800 4616
rect 7840 4564 7892 4616
rect 8944 4607 8996 4616
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 11888 4564 11940 4616
rect 14648 4564 14700 4616
rect 16488 4564 16540 4616
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 1124 4428 1176 4480
rect 2780 4428 2832 4480
rect 4620 4471 4672 4480
rect 4620 4437 4629 4471
rect 4629 4437 4663 4471
rect 4663 4437 4672 4471
rect 4620 4428 4672 4437
rect 4712 4428 4764 4480
rect 7472 4471 7524 4480
rect 7472 4437 7481 4471
rect 7481 4437 7515 4471
rect 7515 4437 7524 4471
rect 7472 4428 7524 4437
rect 18236 4496 18288 4548
rect 21640 4641 21649 4675
rect 21649 4641 21683 4675
rect 21683 4641 21692 4675
rect 21640 4632 21692 4641
rect 10600 4428 10652 4480
rect 12808 4428 12860 4480
rect 18696 4471 18748 4480
rect 18696 4437 18705 4471
rect 18705 4437 18739 4471
rect 18739 4437 18748 4471
rect 18696 4428 18748 4437
rect 19248 4471 19300 4480
rect 19248 4437 19257 4471
rect 19257 4437 19291 4471
rect 19291 4437 19300 4471
rect 19248 4428 19300 4437
rect 19432 4428 19484 4480
rect 19984 4564 20036 4616
rect 20260 4607 20312 4616
rect 20260 4573 20269 4607
rect 20269 4573 20303 4607
rect 20303 4573 20312 4607
rect 20260 4564 20312 4573
rect 20076 4496 20128 4548
rect 21824 4564 21876 4616
rect 23204 4564 23256 4616
rect 24860 4607 24912 4616
rect 24860 4573 24869 4607
rect 24869 4573 24903 4607
rect 24903 4573 24912 4607
rect 24860 4564 24912 4573
rect 25504 4607 25556 4616
rect 25504 4573 25513 4607
rect 25513 4573 25547 4607
rect 25547 4573 25556 4607
rect 25504 4564 25556 4573
rect 20352 4428 20404 4480
rect 20536 4428 20588 4480
rect 23112 4428 23164 4480
rect 24400 4471 24452 4480
rect 24400 4437 24409 4471
rect 24409 4437 24443 4471
rect 24443 4437 24452 4471
rect 24400 4428 24452 4437
rect 24952 4428 25004 4480
rect 26240 4496 26292 4548
rect 26792 4564 26844 4616
rect 27528 4811 27580 4820
rect 27528 4777 27537 4811
rect 27537 4777 27571 4811
rect 27571 4777 27580 4811
rect 27528 4768 27580 4777
rect 28908 4700 28960 4752
rect 41604 4768 41656 4820
rect 41696 4768 41748 4820
rect 42800 4768 42852 4820
rect 46480 4811 46532 4820
rect 46480 4777 46489 4811
rect 46489 4777 46523 4811
rect 46523 4777 46532 4811
rect 46480 4768 46532 4777
rect 29092 4632 29144 4684
rect 34520 4632 34572 4684
rect 40592 4632 40644 4684
rect 32128 4564 32180 4616
rect 32312 4607 32364 4616
rect 32312 4573 32321 4607
rect 32321 4573 32355 4607
rect 32355 4573 32364 4607
rect 32312 4564 32364 4573
rect 32956 4564 33008 4616
rect 35624 4607 35676 4616
rect 35624 4573 35633 4607
rect 35633 4573 35667 4607
rect 35667 4573 35676 4607
rect 35624 4564 35676 4573
rect 35992 4607 36044 4616
rect 27988 4496 28040 4548
rect 32496 4496 32548 4548
rect 35440 4496 35492 4548
rect 35992 4573 36001 4607
rect 36001 4573 36035 4607
rect 36035 4573 36044 4607
rect 35992 4564 36044 4573
rect 36176 4564 36228 4616
rect 36728 4564 36780 4616
rect 37004 4607 37056 4616
rect 37004 4573 37013 4607
rect 37013 4573 37047 4607
rect 37047 4573 37056 4607
rect 37004 4564 37056 4573
rect 37556 4564 37608 4616
rect 38568 4564 38620 4616
rect 40040 4564 40092 4616
rect 42984 4564 43036 4616
rect 43536 4607 43588 4616
rect 43536 4573 43545 4607
rect 43545 4573 43579 4607
rect 43579 4573 43588 4607
rect 43536 4564 43588 4573
rect 44916 4564 44968 4616
rect 46112 4607 46164 4616
rect 31300 4428 31352 4480
rect 32588 4471 32640 4480
rect 32588 4437 32597 4471
rect 32597 4437 32631 4471
rect 32631 4437 32640 4471
rect 32588 4428 32640 4437
rect 36452 4496 36504 4548
rect 39028 4496 39080 4548
rect 40132 4496 40184 4548
rect 40684 4539 40736 4548
rect 40684 4505 40693 4539
rect 40693 4505 40727 4539
rect 40727 4505 40736 4539
rect 40684 4496 40736 4505
rect 46112 4573 46121 4607
rect 46121 4573 46155 4607
rect 46155 4573 46164 4607
rect 46112 4564 46164 4573
rect 46388 4564 46440 4616
rect 47124 4607 47176 4616
rect 47124 4573 47133 4607
rect 47133 4573 47167 4607
rect 47167 4573 47176 4607
rect 47124 4564 47176 4573
rect 47400 4607 47452 4616
rect 47400 4573 47409 4607
rect 47409 4573 47443 4607
rect 47443 4573 47452 4607
rect 48228 4607 48280 4616
rect 47400 4564 47452 4573
rect 48228 4573 48237 4607
rect 48237 4573 48271 4607
rect 48271 4573 48280 4607
rect 48228 4564 48280 4573
rect 46204 4539 46256 4548
rect 36268 4471 36320 4480
rect 36268 4437 36277 4471
rect 36277 4437 36311 4471
rect 36311 4437 36320 4471
rect 36268 4428 36320 4437
rect 38292 4471 38344 4480
rect 38292 4437 38301 4471
rect 38301 4437 38335 4471
rect 38335 4437 38344 4471
rect 38292 4428 38344 4437
rect 40224 4428 40276 4480
rect 46204 4505 46213 4539
rect 46213 4505 46247 4539
rect 46247 4505 46256 4539
rect 46204 4496 46256 4505
rect 42248 4428 42300 4480
rect 45376 4428 45428 4480
rect 46848 4428 46900 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 2136 4224 2188 4276
rect 20536 4224 20588 4276
rect 24860 4224 24912 4276
rect 32588 4224 32640 4276
rect 35808 4224 35860 4276
rect 8668 4156 8720 4208
rect 9956 4156 10008 4208
rect 204 3884 256 3936
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 3424 4088 3476 4140
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 4712 4088 4764 4140
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 5080 4088 5132 4140
rect 4068 4020 4120 4072
rect 7472 4088 7524 4140
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 8484 4131 8536 4140
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 9404 4088 9456 4140
rect 9864 4020 9916 4072
rect 10416 4088 10468 4140
rect 11888 4088 11940 4140
rect 16396 4088 16448 4140
rect 19340 4156 19392 4208
rect 28632 4156 28684 4208
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 18512 4088 18564 4140
rect 18696 4088 18748 4140
rect 11796 4063 11848 4072
rect 11796 4029 11805 4063
rect 11805 4029 11839 4063
rect 11839 4029 11848 4063
rect 11796 4020 11848 4029
rect 13452 4020 13504 4072
rect 15200 4020 15252 4072
rect 16028 4020 16080 4072
rect 19432 4088 19484 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 20168 4020 20220 4072
rect 20260 4020 20312 4072
rect 33140 4088 33192 4140
rect 33508 4088 33560 4140
rect 34520 4131 34572 4140
rect 34520 4097 34529 4131
rect 34529 4097 34563 4131
rect 34563 4097 34572 4131
rect 34520 4088 34572 4097
rect 34704 4131 34756 4140
rect 34704 4097 34713 4131
rect 34713 4097 34747 4131
rect 34747 4097 34756 4131
rect 34704 4088 34756 4097
rect 35532 4156 35584 4208
rect 28264 4063 28316 4072
rect 28264 4029 28273 4063
rect 28273 4029 28307 4063
rect 28307 4029 28316 4063
rect 28264 4020 28316 4029
rect 33692 4020 33744 4072
rect 35624 4088 35676 4140
rect 37556 4224 37608 4276
rect 39028 4224 39080 4276
rect 40960 4224 41012 4276
rect 41052 4224 41104 4276
rect 42800 4267 42852 4276
rect 42800 4233 42825 4267
rect 42825 4233 42852 4267
rect 42984 4267 43036 4276
rect 42800 4224 42852 4233
rect 42984 4233 42993 4267
rect 42993 4233 43027 4267
rect 43027 4233 43036 4267
rect 42984 4224 43036 4233
rect 43536 4224 43588 4276
rect 36544 4156 36596 4208
rect 4620 3952 4672 4004
rect 3608 3884 3660 3936
rect 6276 3952 6328 4004
rect 7472 3952 7524 4004
rect 7564 3952 7616 4004
rect 27252 3952 27304 4004
rect 6552 3884 6604 3936
rect 6644 3884 6696 3936
rect 9220 3884 9272 3936
rect 13452 3884 13504 3936
rect 14004 3884 14056 3936
rect 18788 3884 18840 3936
rect 19432 3884 19484 3936
rect 19524 3884 19576 3936
rect 21548 3884 21600 3936
rect 22652 3884 22704 3936
rect 23480 3884 23532 3936
rect 28172 3884 28224 3936
rect 28448 3884 28500 3936
rect 29460 3884 29512 3936
rect 30012 3952 30064 4004
rect 33416 3952 33468 4004
rect 35440 4020 35492 4072
rect 36176 4131 36228 4140
rect 36176 4097 36190 4131
rect 36190 4097 36224 4131
rect 36224 4097 36228 4131
rect 38476 4131 38528 4140
rect 36176 4088 36228 4097
rect 38476 4097 38485 4131
rect 38485 4097 38519 4131
rect 38519 4097 38528 4131
rect 38476 4088 38528 4097
rect 31576 3884 31628 3936
rect 37372 3952 37424 4004
rect 38660 4088 38712 4140
rect 38844 4131 38896 4140
rect 38844 4097 38853 4131
rect 38853 4097 38887 4131
rect 38887 4097 38896 4131
rect 38844 4088 38896 4097
rect 39028 4088 39080 4140
rect 40224 4088 40276 4140
rect 40592 4088 40644 4140
rect 41052 4088 41104 4140
rect 41328 4088 41380 4140
rect 42708 4156 42760 4208
rect 46112 4199 46164 4208
rect 46112 4165 46121 4199
rect 46121 4165 46155 4199
rect 46155 4165 46164 4199
rect 46112 4156 46164 4165
rect 45928 4131 45980 4140
rect 42892 4020 42944 4072
rect 45928 4097 45937 4131
rect 45937 4097 45971 4131
rect 45971 4097 45980 4131
rect 45928 4088 45980 4097
rect 46020 4088 46072 4140
rect 46848 4156 46900 4208
rect 46940 4156 46992 4208
rect 48228 4156 48280 4208
rect 46296 4131 46348 4140
rect 46296 4097 46305 4131
rect 46305 4097 46339 4131
rect 46339 4097 46348 4131
rect 46296 4088 46348 4097
rect 46480 4088 46532 4140
rect 45468 4020 45520 4072
rect 45836 3952 45888 4004
rect 47400 3952 47452 4004
rect 34704 3884 34756 3936
rect 36360 3927 36412 3936
rect 36360 3893 36369 3927
rect 36369 3893 36403 3927
rect 36403 3893 36412 3927
rect 36360 3884 36412 3893
rect 39120 3927 39172 3936
rect 39120 3893 39129 3927
rect 39129 3893 39163 3927
rect 39163 3893 39172 3927
rect 39120 3884 39172 3893
rect 39856 3927 39908 3936
rect 39856 3893 39865 3927
rect 39865 3893 39899 3927
rect 39899 3893 39908 3927
rect 39856 3884 39908 3893
rect 41144 3884 41196 3936
rect 42616 3884 42668 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2136 3680 2188 3732
rect 4804 3680 4856 3732
rect 4988 3680 5040 3732
rect 7564 3680 7616 3732
rect 4896 3612 4948 3664
rect 8208 3680 8260 3732
rect 11152 3680 11204 3732
rect 11796 3680 11848 3732
rect 12072 3680 12124 3732
rect 21916 3680 21968 3732
rect 1860 3519 1912 3528
rect 1860 3485 1869 3519
rect 1869 3485 1903 3519
rect 1903 3485 1912 3519
rect 1860 3476 1912 3485
rect 3516 3476 3568 3528
rect 3884 3476 3936 3528
rect 5080 3544 5132 3596
rect 5264 3587 5316 3596
rect 5264 3553 5273 3587
rect 5273 3553 5307 3587
rect 5307 3553 5316 3587
rect 5264 3544 5316 3553
rect 6736 3544 6788 3596
rect 3700 3408 3752 3460
rect 6920 3476 6972 3528
rect 9864 3544 9916 3596
rect 7472 3519 7524 3528
rect 664 3340 716 3392
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 6368 3408 6420 3460
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 7564 3476 7616 3528
rect 10232 3476 10284 3528
rect 10600 3476 10652 3528
rect 10692 3476 10744 3528
rect 11336 3544 11388 3596
rect 12072 3544 12124 3596
rect 15108 3612 15160 3664
rect 15568 3655 15620 3664
rect 15568 3621 15577 3655
rect 15577 3621 15611 3655
rect 15611 3621 15620 3655
rect 15568 3612 15620 3621
rect 16396 3612 16448 3664
rect 23664 3655 23716 3664
rect 23664 3621 23673 3655
rect 23673 3621 23707 3655
rect 23707 3621 23716 3655
rect 23664 3612 23716 3621
rect 26240 3612 26292 3664
rect 27252 3680 27304 3732
rect 33324 3680 33376 3732
rect 33416 3680 33468 3732
rect 35532 3680 35584 3732
rect 37464 3680 37516 3732
rect 40224 3723 40276 3732
rect 40224 3689 40233 3723
rect 40233 3689 40267 3723
rect 40267 3689 40276 3723
rect 40224 3680 40276 3689
rect 33048 3612 33100 3664
rect 6644 3383 6696 3392
rect 6644 3349 6653 3383
rect 6653 3349 6687 3383
rect 6687 3349 6696 3383
rect 6644 3340 6696 3349
rect 6828 3340 6880 3392
rect 11888 3476 11940 3528
rect 13360 3476 13412 3528
rect 11244 3408 11296 3460
rect 12900 3408 12952 3460
rect 14004 3408 14056 3460
rect 9864 3383 9916 3392
rect 9864 3349 9873 3383
rect 9873 3349 9907 3383
rect 9907 3349 9916 3383
rect 9864 3340 9916 3349
rect 11152 3340 11204 3392
rect 11704 3340 11756 3392
rect 12164 3383 12216 3392
rect 12164 3349 12173 3383
rect 12173 3349 12207 3383
rect 12207 3349 12216 3383
rect 12164 3340 12216 3349
rect 13820 3340 13872 3392
rect 14556 3340 14608 3392
rect 15016 3519 15068 3528
rect 15016 3485 15026 3519
rect 15026 3485 15060 3519
rect 15060 3485 15068 3519
rect 16304 3544 16356 3596
rect 15016 3476 15068 3485
rect 15568 3476 15620 3528
rect 16028 3519 16080 3528
rect 16028 3485 16037 3519
rect 16037 3485 16071 3519
rect 16071 3485 16080 3519
rect 16028 3476 16080 3485
rect 16212 3519 16264 3528
rect 16212 3485 16219 3519
rect 16219 3485 16264 3519
rect 16212 3476 16264 3485
rect 16488 3519 16540 3528
rect 16488 3485 16502 3519
rect 16502 3485 16536 3519
rect 16536 3485 16540 3519
rect 16488 3476 16540 3485
rect 17132 3476 17184 3528
rect 17408 3544 17460 3596
rect 18696 3476 18748 3528
rect 20260 3519 20312 3528
rect 20260 3485 20269 3519
rect 20269 3485 20303 3519
rect 20303 3485 20312 3519
rect 20260 3476 20312 3485
rect 21088 3476 21140 3528
rect 21548 3544 21600 3596
rect 22560 3544 22612 3596
rect 28172 3544 28224 3596
rect 30564 3544 30616 3596
rect 23480 3476 23532 3528
rect 23572 3476 23624 3528
rect 14832 3408 14884 3460
rect 15200 3451 15252 3460
rect 15200 3417 15209 3451
rect 15209 3417 15243 3451
rect 15243 3417 15252 3451
rect 15200 3408 15252 3417
rect 16028 3340 16080 3392
rect 16488 3340 16540 3392
rect 16580 3340 16632 3392
rect 19156 3408 19208 3460
rect 21824 3408 21876 3460
rect 23664 3408 23716 3460
rect 24952 3476 25004 3528
rect 26148 3476 26200 3528
rect 26332 3476 26384 3528
rect 27436 3476 27488 3528
rect 33140 3544 33192 3596
rect 34060 3612 34112 3664
rect 35532 3544 35584 3596
rect 36912 3544 36964 3596
rect 31116 3519 31168 3528
rect 31116 3485 31125 3519
rect 31125 3485 31159 3519
rect 31159 3485 31168 3519
rect 31116 3476 31168 3485
rect 31300 3519 31352 3528
rect 31300 3485 31309 3519
rect 31309 3485 31343 3519
rect 31343 3485 31352 3519
rect 31300 3476 31352 3485
rect 33416 3519 33468 3528
rect 33416 3485 33425 3519
rect 33425 3485 33459 3519
rect 33459 3485 33468 3519
rect 33416 3476 33468 3485
rect 25412 3408 25464 3460
rect 33324 3408 33376 3460
rect 17500 3340 17552 3392
rect 20168 3340 20220 3392
rect 21180 3383 21232 3392
rect 21180 3349 21189 3383
rect 21189 3349 21223 3383
rect 21223 3349 21232 3383
rect 21180 3340 21232 3349
rect 22192 3340 22244 3392
rect 22836 3340 22888 3392
rect 27988 3340 28040 3392
rect 28080 3383 28132 3392
rect 28080 3349 28089 3383
rect 28089 3349 28123 3383
rect 28123 3349 28132 3383
rect 30472 3383 30524 3392
rect 28080 3340 28132 3349
rect 30472 3349 30481 3383
rect 30481 3349 30515 3383
rect 30515 3349 30524 3383
rect 30472 3340 30524 3349
rect 33692 3340 33744 3392
rect 33784 3340 33836 3392
rect 34796 3476 34848 3528
rect 35348 3476 35400 3528
rect 37188 3476 37240 3528
rect 37556 3544 37608 3596
rect 38844 3544 38896 3596
rect 39120 3544 39172 3596
rect 37464 3519 37516 3528
rect 37464 3485 37473 3519
rect 37473 3485 37507 3519
rect 37507 3485 37516 3519
rect 37464 3476 37516 3485
rect 37740 3476 37792 3528
rect 38292 3519 38344 3528
rect 38292 3485 38301 3519
rect 38301 3485 38335 3519
rect 38335 3485 38344 3519
rect 38292 3476 38344 3485
rect 38384 3476 38436 3528
rect 39948 3476 40000 3528
rect 41420 3519 41472 3528
rect 41420 3485 41429 3519
rect 41429 3485 41463 3519
rect 41463 3485 41472 3519
rect 42156 3519 42208 3528
rect 41420 3476 41472 3485
rect 42156 3485 42165 3519
rect 42165 3485 42199 3519
rect 42199 3485 42208 3519
rect 42156 3476 42208 3485
rect 42248 3476 42300 3528
rect 42708 3476 42760 3528
rect 43996 3612 44048 3664
rect 57152 3612 57204 3664
rect 45744 3544 45796 3596
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 46020 3476 46072 3528
rect 34336 3408 34388 3460
rect 46756 3451 46808 3460
rect 46756 3417 46790 3451
rect 46790 3417 46808 3451
rect 46756 3408 46808 3417
rect 58164 3476 58216 3528
rect 34060 3340 34112 3392
rect 35348 3340 35400 3392
rect 37832 3383 37884 3392
rect 37832 3349 37841 3383
rect 37841 3349 37875 3383
rect 37875 3349 37884 3383
rect 37832 3340 37884 3349
rect 38200 3340 38252 3392
rect 39672 3340 39724 3392
rect 45468 3340 45520 3392
rect 46204 3340 46256 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 3332 3136 3384 3188
rect 3884 3179 3936 3188
rect 3884 3145 3893 3179
rect 3893 3145 3927 3179
rect 3927 3145 3936 3179
rect 3884 3136 3936 3145
rect 6368 3179 6420 3188
rect 3608 3068 3660 3120
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 3516 2975 3568 2984
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 3516 2932 3568 2941
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 4988 3000 5040 3052
rect 7104 3000 7156 3052
rect 6644 2932 6696 2984
rect 21640 3136 21692 3188
rect 33508 3179 33560 3188
rect 9864 3111 9916 3120
rect 7472 3000 7524 3052
rect 9864 3077 9898 3111
rect 9898 3077 9916 3111
rect 9864 3068 9916 3077
rect 10876 3068 10928 3120
rect 11244 3068 11296 3120
rect 12164 3068 12216 3120
rect 11704 3043 11756 3052
rect 7932 2932 7984 2984
rect 8944 2932 8996 2984
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 12808 3043 12860 3052
rect 12808 3009 12817 3043
rect 12817 3009 12851 3043
rect 12851 3009 12860 3043
rect 12808 3000 12860 3009
rect 14464 3068 14516 3120
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 14556 3000 14608 3052
rect 14924 3111 14976 3120
rect 14924 3077 14933 3111
rect 14933 3077 14967 3111
rect 14967 3077 14976 3111
rect 14924 3068 14976 3077
rect 16488 3068 16540 3120
rect 15016 3043 15068 3052
rect 15016 3009 15025 3043
rect 15025 3009 15059 3043
rect 15059 3009 15068 3043
rect 15016 3000 15068 3009
rect 15292 3000 15344 3052
rect 16028 3000 16080 3052
rect 16856 3000 16908 3052
rect 18144 3068 18196 3120
rect 18788 3068 18840 3120
rect 19248 3068 19300 3120
rect 15568 2932 15620 2984
rect 17132 3043 17184 3052
rect 17132 3009 17146 3043
rect 17146 3009 17180 3043
rect 17180 3009 17184 3043
rect 17132 3000 17184 3009
rect 22652 3068 22704 3120
rect 24400 3068 24452 3120
rect 27620 3111 27672 3120
rect 27620 3077 27654 3111
rect 27654 3077 27672 3111
rect 27620 3068 27672 3077
rect 28264 3068 28316 3120
rect 30472 3111 30524 3120
rect 30472 3077 30506 3111
rect 30506 3077 30524 3111
rect 30472 3068 30524 3077
rect 23664 3043 23716 3052
rect 17500 2932 17552 2984
rect 18144 2932 18196 2984
rect 20444 2932 20496 2984
rect 23664 3009 23673 3043
rect 23673 3009 23707 3043
rect 23707 3009 23716 3043
rect 23664 3000 23716 3009
rect 21824 2975 21876 2984
rect 21824 2941 21833 2975
rect 21833 2941 21867 2975
rect 21867 2941 21876 2975
rect 21824 2932 21876 2941
rect 22836 2932 22888 2984
rect 4068 2864 4120 2916
rect 6460 2864 6512 2916
rect 7656 2864 7708 2916
rect 2596 2796 2648 2848
rect 7748 2796 7800 2848
rect 9496 2796 9548 2848
rect 10600 2864 10652 2916
rect 12900 2864 12952 2916
rect 14740 2864 14792 2916
rect 14832 2864 14884 2916
rect 17224 2864 17276 2916
rect 10692 2796 10744 2848
rect 12072 2796 12124 2848
rect 15200 2796 15252 2848
rect 16948 2796 17000 2848
rect 17684 2796 17736 2848
rect 18052 2796 18104 2848
rect 20076 2839 20128 2848
rect 20076 2805 20085 2839
rect 20085 2805 20119 2839
rect 20119 2805 20128 2839
rect 20076 2796 20128 2805
rect 20260 2796 20312 2848
rect 23204 2839 23256 2848
rect 23204 2805 23213 2839
rect 23213 2805 23247 2839
rect 23247 2805 23256 2839
rect 25596 2864 25648 2916
rect 23204 2796 23256 2805
rect 24860 2796 24912 2848
rect 25964 3000 26016 3052
rect 26148 2932 26200 2984
rect 31852 3000 31904 3052
rect 32128 3043 32180 3052
rect 32128 3009 32137 3043
rect 32137 3009 32171 3043
rect 32171 3009 32180 3043
rect 32128 3000 32180 3009
rect 33508 3145 33517 3179
rect 33517 3145 33551 3179
rect 33551 3145 33560 3179
rect 33508 3136 33560 3145
rect 33784 3136 33836 3188
rect 34152 3136 34204 3188
rect 34060 3068 34112 3120
rect 34704 3111 34756 3120
rect 34704 3077 34738 3111
rect 34738 3077 34756 3111
rect 34704 3068 34756 3077
rect 35808 3136 35860 3188
rect 37740 3136 37792 3188
rect 38844 3136 38896 3188
rect 44088 3136 44140 3188
rect 54852 3136 54904 3188
rect 34336 3000 34388 3052
rect 35440 3000 35492 3052
rect 35716 3000 35768 3052
rect 37832 3068 37884 3120
rect 39856 3068 39908 3120
rect 41420 3068 41472 3120
rect 43812 3111 43864 3120
rect 40316 3000 40368 3052
rect 42156 3000 42208 3052
rect 42708 3043 42760 3052
rect 42708 3009 42717 3043
rect 42717 3009 42751 3043
rect 42751 3009 42760 3043
rect 42708 3000 42760 3009
rect 43812 3077 43846 3111
rect 43846 3077 43864 3111
rect 43812 3068 43864 3077
rect 45376 3068 45428 3120
rect 45928 3068 45980 3120
rect 46204 3000 46256 3052
rect 48412 3068 48464 3120
rect 35532 2932 35584 2984
rect 37280 2932 37332 2984
rect 49608 3000 49660 3052
rect 50988 3000 51040 3052
rect 52460 3068 52512 3120
rect 57152 3111 57204 3120
rect 57152 3077 57161 3111
rect 57161 3077 57195 3111
rect 57195 3077 57204 3111
rect 57152 3068 57204 3077
rect 26056 2907 26108 2916
rect 26056 2873 26065 2907
rect 26065 2873 26099 2907
rect 26099 2873 26108 2907
rect 26056 2864 26108 2873
rect 29552 2864 29604 2916
rect 31576 2839 31628 2848
rect 31576 2805 31585 2839
rect 31585 2805 31619 2839
rect 31619 2805 31628 2839
rect 31576 2796 31628 2805
rect 34336 2864 34388 2916
rect 33784 2796 33836 2848
rect 35716 2796 35768 2848
rect 36728 2796 36780 2848
rect 38660 2796 38712 2848
rect 42616 2796 42668 2848
rect 44916 2907 44968 2916
rect 44916 2873 44925 2907
rect 44925 2873 44959 2907
rect 44959 2873 44968 2907
rect 44916 2864 44968 2873
rect 45744 2796 45796 2848
rect 45836 2796 45888 2848
rect 51540 2932 51592 2984
rect 59636 2932 59688 2984
rect 47032 2864 47084 2916
rect 49884 2796 49936 2848
rect 51356 2796 51408 2848
rect 52828 2796 52880 2848
rect 54300 2796 54352 2848
rect 55772 2796 55824 2848
rect 58716 2796 58768 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2044 2592 2096 2644
rect 3056 2592 3108 2644
rect 5448 2592 5500 2644
rect 7012 2592 7064 2644
rect 13268 2592 13320 2644
rect 15384 2592 15436 2644
rect 18420 2592 18472 2644
rect 21364 2592 21416 2644
rect 28816 2635 28868 2644
rect 28816 2601 28825 2635
rect 28825 2601 28859 2635
rect 28859 2601 28868 2635
rect 28816 2592 28868 2601
rect 29368 2592 29420 2644
rect 29828 2592 29880 2644
rect 30288 2635 30340 2644
rect 30288 2601 30297 2635
rect 30297 2601 30331 2635
rect 30331 2601 30340 2635
rect 30288 2592 30340 2601
rect 32864 2592 32916 2644
rect 38660 2592 38712 2644
rect 6000 2524 6052 2576
rect 9404 2524 9456 2576
rect 12348 2524 12400 2576
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 4528 2388 4580 2440
rect 13728 2456 13780 2508
rect 1492 2363 1544 2372
rect 1492 2329 1501 2363
rect 1501 2329 1535 2363
rect 1535 2329 1544 2363
rect 1492 2320 1544 2329
rect 6552 2388 6604 2440
rect 8944 2431 8996 2440
rect 8944 2397 8953 2431
rect 8953 2397 8987 2431
rect 8987 2397 8996 2431
rect 8944 2388 8996 2397
rect 9496 2431 9548 2440
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 10508 2388 10560 2440
rect 12072 2431 12124 2440
rect 7012 2320 7064 2372
rect 3056 2252 3108 2304
rect 5540 2252 5592 2304
rect 6644 2252 6696 2304
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 12992 2431 13044 2440
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 16856 2524 16908 2576
rect 18328 2524 18380 2576
rect 14556 2388 14608 2440
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 15568 2388 15620 2440
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 25044 2524 25096 2576
rect 29644 2524 29696 2576
rect 18788 2456 18840 2508
rect 19248 2499 19300 2508
rect 19248 2465 19257 2499
rect 19257 2465 19291 2499
rect 19291 2465 19300 2499
rect 19248 2456 19300 2465
rect 29460 2456 29512 2508
rect 18420 2388 18472 2397
rect 8484 2252 8536 2304
rect 9220 2252 9272 2304
rect 11336 2252 11388 2304
rect 11888 2252 11940 2304
rect 13728 2252 13780 2304
rect 19248 2320 19300 2372
rect 14280 2252 14332 2304
rect 16764 2252 16816 2304
rect 17224 2252 17276 2304
rect 19156 2252 19208 2304
rect 19524 2431 19576 2440
rect 19524 2397 19558 2431
rect 19558 2397 19576 2431
rect 19524 2388 19576 2397
rect 22284 2388 22336 2440
rect 22560 2431 22612 2440
rect 22560 2397 22569 2431
rect 22569 2397 22603 2431
rect 22603 2397 22612 2431
rect 22560 2388 22612 2397
rect 23296 2431 23348 2440
rect 23296 2397 23305 2431
rect 23305 2397 23339 2431
rect 23339 2397 23348 2431
rect 23296 2388 23348 2397
rect 24768 2388 24820 2440
rect 24860 2388 24912 2440
rect 25688 2388 25740 2440
rect 26240 2388 26292 2440
rect 28080 2431 28132 2440
rect 28080 2397 28089 2431
rect 28089 2397 28123 2431
rect 28123 2397 28132 2431
rect 28080 2388 28132 2397
rect 28908 2388 28960 2440
rect 29552 2431 29604 2440
rect 29552 2397 29561 2431
rect 29561 2397 29595 2431
rect 29595 2397 29604 2431
rect 29552 2388 29604 2397
rect 29736 2388 29788 2440
rect 30380 2388 30432 2440
rect 31392 2456 31444 2508
rect 33324 2456 33376 2508
rect 35164 2524 35216 2576
rect 35072 2456 35124 2508
rect 54392 2456 54444 2508
rect 31852 2388 31904 2440
rect 33600 2388 33652 2440
rect 19432 2320 19484 2372
rect 29828 2320 29880 2372
rect 34152 2388 34204 2440
rect 37372 2388 37424 2440
rect 42432 2388 42484 2440
rect 48504 2388 48556 2440
rect 52368 2388 52420 2440
rect 53840 2388 53892 2440
rect 55220 2388 55272 2440
rect 56692 2388 56744 2440
rect 21640 2252 21692 2304
rect 22100 2252 22152 2304
rect 22836 2252 22888 2304
rect 24032 2252 24084 2304
rect 24676 2252 24728 2304
rect 26516 2252 26568 2304
rect 27988 2252 28040 2304
rect 29460 2252 29512 2304
rect 30840 2252 30892 2304
rect 32312 2252 32364 2304
rect 36268 2320 36320 2372
rect 37740 2320 37792 2372
rect 39212 2320 39264 2372
rect 40592 2320 40644 2372
rect 42064 2320 42116 2372
rect 43536 2320 43588 2372
rect 45008 2320 45060 2372
rect 46480 2320 46532 2372
rect 47952 2320 48004 2372
rect 49424 2320 49476 2372
rect 50896 2320 50948 2372
rect 53012 2363 53064 2372
rect 53012 2329 53021 2363
rect 53021 2329 53055 2363
rect 53055 2329 53064 2363
rect 53012 2320 53064 2329
rect 54208 2363 54260 2372
rect 54208 2329 54217 2363
rect 54217 2329 54251 2363
rect 54251 2329 54260 2363
rect 54208 2320 54260 2329
rect 55588 2363 55640 2372
rect 55588 2329 55597 2363
rect 55597 2329 55631 2363
rect 55631 2329 55640 2363
rect 55588 2320 55640 2329
rect 57060 2363 57112 2372
rect 57060 2329 57069 2363
rect 57069 2329 57103 2363
rect 57103 2329 57112 2363
rect 57060 2320 57112 2329
rect 40500 2252 40552 2304
rect 43812 2295 43864 2304
rect 43812 2261 43821 2295
rect 43821 2261 43855 2295
rect 43855 2261 43864 2295
rect 43812 2252 43864 2261
rect 45560 2295 45612 2304
rect 45560 2261 45569 2295
rect 45569 2261 45603 2295
rect 45603 2261 45612 2295
rect 46756 2295 46808 2304
rect 45560 2252 45612 2261
rect 46756 2261 46765 2295
rect 46765 2261 46799 2295
rect 46799 2261 46808 2295
rect 46756 2252 46808 2261
rect 48228 2295 48280 2304
rect 48228 2261 48237 2295
rect 48237 2261 48271 2295
rect 48271 2261 48280 2295
rect 48228 2252 48280 2261
rect 48412 2252 48464 2304
rect 50712 2295 50764 2304
rect 50712 2261 50721 2295
rect 50721 2261 50755 2295
rect 50755 2261 50764 2295
rect 50712 2252 50764 2261
rect 51632 2295 51684 2304
rect 51632 2261 51641 2295
rect 51641 2261 51675 2295
rect 51675 2261 51684 2295
rect 51632 2252 51684 2261
rect 57244 2252 57296 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 10508 2048 10560 2100
rect 34152 2048 34204 2100
rect 34244 2048 34296 2100
rect 12992 1980 13044 2032
rect 35808 1980 35860 2032
rect 35900 1980 35952 2032
rect 40684 1980 40736 2032
rect 46756 1980 46808 2032
rect 8944 1912 8996 1964
rect 16120 1912 16172 1964
rect 16856 1912 16908 1964
rect 22468 1912 22520 1964
rect 33968 1912 34020 1964
rect 48228 1912 48280 1964
rect 9128 1844 9180 1896
rect 55588 1844 55640 1896
rect 12532 1776 12584 1828
rect 51632 1776 51684 1828
rect 12900 1708 12952 1760
rect 50712 1708 50764 1760
rect 10600 1640 10652 1692
rect 53012 1640 53064 1692
rect 8668 1572 8720 1624
rect 54208 1572 54260 1624
rect 9312 1504 9364 1556
rect 57060 1504 57112 1556
rect 15752 1436 15804 1488
rect 23204 1436 23256 1488
rect 23296 1436 23348 1488
rect 33508 1436 33560 1488
rect 33876 1436 33928 1488
rect 5080 1368 5132 1420
rect 6644 1368 6696 1420
rect 19708 1368 19760 1420
rect 20260 1368 20312 1420
rect 33232 1368 33284 1420
rect 40500 1368 40552 1420
rect 40684 1436 40736 1488
rect 43812 1436 43864 1488
rect 45560 1368 45612 1420
<< metal2 >>
rect 2870 41712 2926 41721
rect 2870 41647 2926 41656
rect 2778 40080 2834 40089
rect 2778 40015 2834 40024
rect 2792 39642 2820 40015
rect 2780 39636 2832 39642
rect 2780 39578 2832 39584
rect 1492 39432 1544 39438
rect 1492 39374 1544 39380
rect 1400 32428 1452 32434
rect 1400 32370 1452 32376
rect 1412 32065 1440 32370
rect 1398 32056 1454 32065
rect 1398 31991 1454 32000
rect 1504 30818 1532 39374
rect 1584 39296 1636 39302
rect 1582 39264 1584 39273
rect 1636 39264 1638 39273
rect 1582 39199 1638 39208
rect 1584 38752 1636 38758
rect 1584 38694 1636 38700
rect 1596 38457 1624 38694
rect 2884 38554 2912 41647
rect 3698 41200 3754 42000
rect 11150 41200 11206 42000
rect 18694 41200 18750 42000
rect 26146 41200 26202 42000
rect 33690 41200 33746 42000
rect 41142 41200 41198 42000
rect 48686 41200 48742 42000
rect 56138 41200 56194 42000
rect 3054 40896 3110 40905
rect 3054 40831 3110 40840
rect 3068 39642 3096 40831
rect 3712 39642 3740 41200
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 3056 39636 3108 39642
rect 3056 39578 3108 39584
rect 3700 39636 3752 39642
rect 3700 39578 3752 39584
rect 18708 39506 18736 41200
rect 26160 39658 26188 41200
rect 26160 39642 26280 39658
rect 26160 39636 26292 39642
rect 26160 39630 26240 39636
rect 26240 39578 26292 39584
rect 8852 39500 8904 39506
rect 8852 39442 8904 39448
rect 18696 39500 18748 39506
rect 18696 39442 18748 39448
rect 3240 39432 3292 39438
rect 3240 39374 3292 39380
rect 2872 38548 2924 38554
rect 2872 38490 2924 38496
rect 1582 38448 1638 38457
rect 1582 38383 1638 38392
rect 2412 38344 2464 38350
rect 2412 38286 2464 38292
rect 1768 37868 1820 37874
rect 1768 37810 1820 37816
rect 1584 37664 1636 37670
rect 1582 37632 1584 37641
rect 1636 37632 1638 37641
rect 1582 37567 1638 37576
rect 1676 36780 1728 36786
rect 1676 36722 1728 36728
rect 1582 36680 1638 36689
rect 1582 36615 1584 36624
rect 1636 36615 1638 36624
rect 1584 36586 1636 36592
rect 1584 36032 1636 36038
rect 1584 35974 1636 35980
rect 1596 35873 1624 35974
rect 1582 35864 1638 35873
rect 1582 35799 1638 35808
rect 1582 35048 1638 35057
rect 1582 34983 1638 34992
rect 1596 34746 1624 34983
rect 1584 34740 1636 34746
rect 1584 34682 1636 34688
rect 1584 33856 1636 33862
rect 1582 33824 1584 33833
rect 1636 33824 1638 33833
rect 1582 33759 1638 33768
rect 1584 32768 1636 32774
rect 1584 32710 1636 32716
rect 1596 32473 1624 32710
rect 1582 32464 1638 32473
rect 1582 32399 1638 32408
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1596 31657 1624 31758
rect 1582 31648 1638 31657
rect 1582 31583 1638 31592
rect 1582 31240 1638 31249
rect 1688 31210 1716 36722
rect 1582 31175 1638 31184
rect 1676 31204 1728 31210
rect 1596 30938 1624 31175
rect 1676 31146 1728 31152
rect 1584 30932 1636 30938
rect 1584 30874 1636 30880
rect 1504 30790 1716 30818
rect 1492 30728 1544 30734
rect 1492 30670 1544 30676
rect 1400 30252 1452 30258
rect 1400 30194 1452 30200
rect 1412 29850 1440 30194
rect 1400 29844 1452 29850
rect 1400 29786 1452 29792
rect 1504 27334 1532 30670
rect 1584 30048 1636 30054
rect 1582 30016 1584 30025
rect 1636 30016 1638 30025
rect 1582 29951 1638 29960
rect 1584 27872 1636 27878
rect 1584 27814 1636 27820
rect 1596 27441 1624 27814
rect 1582 27432 1638 27441
rect 1582 27367 1638 27376
rect 1492 27328 1544 27334
rect 1492 27270 1544 27276
rect 1492 27056 1544 27062
rect 1490 27024 1492 27033
rect 1544 27024 1546 27033
rect 1490 26959 1546 26968
rect 1584 26240 1636 26246
rect 1584 26182 1636 26188
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1412 25809 1440 25842
rect 1398 25800 1454 25809
rect 1398 25735 1454 25744
rect 1596 24993 1624 26182
rect 1688 25974 1716 30790
rect 1676 25968 1728 25974
rect 1676 25910 1728 25916
rect 1780 25498 1808 37810
rect 2424 35894 2452 38286
rect 2424 35866 2544 35894
rect 1860 35012 1912 35018
rect 1860 34954 1912 34960
rect 1872 34649 1900 34954
rect 1952 34944 2004 34950
rect 1952 34886 2004 34892
rect 1858 34640 1914 34649
rect 1858 34575 1914 34584
rect 1860 33516 1912 33522
rect 1860 33458 1912 33464
rect 1872 33425 1900 33458
rect 1858 33416 1914 33425
rect 1858 33351 1914 33360
rect 1860 31340 1912 31346
rect 1860 31282 1912 31288
rect 1872 30841 1900 31282
rect 1858 30832 1914 30841
rect 1858 30767 1914 30776
rect 1858 29608 1914 29617
rect 1858 29543 1914 29552
rect 1872 29238 1900 29543
rect 1860 29232 1912 29238
rect 1860 29174 1912 29180
rect 1860 28484 1912 28490
rect 1860 28426 1912 28432
rect 1872 28393 1900 28426
rect 1858 28384 1914 28393
rect 1858 28319 1914 28328
rect 1860 27464 1912 27470
rect 1860 27406 1912 27412
rect 1872 26314 1900 27406
rect 1860 26308 1912 26314
rect 1860 26250 1912 26256
rect 1768 25492 1820 25498
rect 1768 25434 1820 25440
rect 1872 25362 1900 26250
rect 1860 25356 1912 25362
rect 1860 25298 1912 25304
rect 1582 24984 1638 24993
rect 1582 24919 1638 24928
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1412 24585 1440 24754
rect 1398 24576 1454 24585
rect 1398 24511 1454 24520
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 24041 1440 24142
rect 1584 24064 1636 24070
rect 1398 24032 1454 24041
rect 1584 24006 1636 24012
rect 1398 23967 1454 23976
rect 1596 23769 1624 24006
rect 1582 23760 1638 23769
rect 1400 23724 1452 23730
rect 1582 23695 1638 23704
rect 1400 23666 1452 23672
rect 1412 23225 1440 23666
rect 1584 23520 1636 23526
rect 1584 23462 1636 23468
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 21593 1440 23054
rect 1596 22778 1624 23462
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1584 22432 1636 22438
rect 1582 22400 1584 22409
rect 1636 22400 1638 22409
rect 1582 22335 1638 22344
rect 1860 22024 1912 22030
rect 1858 21992 1860 22001
rect 1912 21992 1914 22001
rect 1858 21927 1914 21936
rect 1398 21584 1454 21593
rect 1398 21519 1454 21528
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 21185 1624 21286
rect 1582 21176 1638 21185
rect 1582 21111 1638 21120
rect 1676 20868 1728 20874
rect 1676 20810 1728 20816
rect 1688 20777 1716 20810
rect 1674 20768 1730 20777
rect 1674 20703 1730 20712
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 19961 1624 20198
rect 1582 19952 1638 19961
rect 1582 19887 1638 19896
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1412 19553 1440 19790
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 1398 19544 1454 19553
rect 1398 19479 1454 19488
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 18970 1440 19314
rect 1492 19304 1544 19310
rect 1492 19246 1544 19252
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1504 18834 1532 19246
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1492 18828 1544 18834
rect 1492 18770 1544 18776
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 18193 1440 18226
rect 1398 18184 1454 18193
rect 1398 18119 1454 18128
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1412 16454 1440 17614
rect 1504 16658 1532 18770
rect 1596 18601 1624 19110
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1582 18592 1638 18601
rect 1582 18527 1638 18536
rect 1688 18426 1716 18702
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1400 16448 1452 16454
rect 1400 16390 1452 16396
rect 1596 16153 1624 17478
rect 1582 16144 1638 16153
rect 1492 16108 1544 16114
rect 1582 16079 1638 16088
rect 1492 16050 1544 16056
rect 1504 15745 1532 16050
rect 1490 15736 1546 15745
rect 1490 15671 1546 15680
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1412 14521 1440 14962
rect 1596 14929 1624 15302
rect 1582 14920 1638 14929
rect 1582 14855 1638 14864
rect 1398 14512 1454 14521
rect 1398 14447 1454 14456
rect 1780 14278 1808 19654
rect 1964 18358 1992 34886
rect 2320 34604 2372 34610
rect 2320 34546 2372 34552
rect 2332 34241 2360 34546
rect 2318 34232 2374 34241
rect 2318 34167 2374 34176
rect 2044 33380 2096 33386
rect 2044 33322 2096 33328
rect 2056 19786 2084 33322
rect 2228 32224 2280 32230
rect 2228 32166 2280 32172
rect 2136 28416 2188 28422
rect 2136 28358 2188 28364
rect 2148 28218 2176 28358
rect 2136 28212 2188 28218
rect 2136 28154 2188 28160
rect 2136 27872 2188 27878
rect 2136 27814 2188 27820
rect 2148 27470 2176 27814
rect 2136 27464 2188 27470
rect 2136 27406 2188 27412
rect 2240 26234 2268 32166
rect 2320 31204 2372 31210
rect 2320 31146 2372 31152
rect 2332 27010 2360 31146
rect 2412 28076 2464 28082
rect 2412 28018 2464 28024
rect 2424 27130 2452 28018
rect 2412 27124 2464 27130
rect 2412 27066 2464 27072
rect 2332 26982 2452 27010
rect 2148 26206 2268 26234
rect 2320 26240 2372 26246
rect 2318 26208 2320 26217
rect 2372 26208 2374 26217
rect 2044 19780 2096 19786
rect 2044 19722 2096 19728
rect 1952 18352 2004 18358
rect 1952 18294 2004 18300
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 1872 16969 1900 17138
rect 1858 16960 1914 16969
rect 1858 16895 1914 16904
rect 2148 16574 2176 26206
rect 2318 26143 2374 26152
rect 2320 25900 2372 25906
rect 2320 25842 2372 25848
rect 2332 25401 2360 25842
rect 2318 25392 2374 25401
rect 2318 25327 2374 25336
rect 2320 25220 2372 25226
rect 2320 25162 2372 25168
rect 2332 24954 2360 25162
rect 2320 24948 2372 24954
rect 2320 24890 2372 24896
rect 2228 24812 2280 24818
rect 2228 24754 2280 24760
rect 2240 24410 2268 24754
rect 2424 24682 2452 26982
rect 2412 24676 2464 24682
rect 2412 24618 2464 24624
rect 2228 24404 2280 24410
rect 2228 24346 2280 24352
rect 2516 23254 2544 35866
rect 2872 33516 2924 33522
rect 2872 33458 2924 33464
rect 2884 33017 2912 33458
rect 2870 33008 2926 33017
rect 2870 32943 2926 32952
rect 3252 31754 3280 39374
rect 4436 39296 4488 39302
rect 4436 39238 4488 39244
rect 4448 39098 4476 39238
rect 4436 39092 4488 39098
rect 4436 39034 4488 39040
rect 7196 38956 7248 38962
rect 7196 38898 7248 38904
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 7208 35894 7236 38898
rect 8864 35894 8892 39442
rect 33704 39438 33732 41200
rect 41156 39930 41184 41200
rect 41156 39902 41460 39930
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 41432 39642 41460 39902
rect 48700 39642 48728 41200
rect 56152 39642 56180 41200
rect 41420 39636 41472 39642
rect 41420 39578 41472 39584
rect 48688 39636 48740 39642
rect 48688 39578 48740 39584
rect 56140 39636 56192 39642
rect 56140 39578 56192 39584
rect 26976 39432 27028 39438
rect 26976 39374 27028 39380
rect 33692 39432 33744 39438
rect 33692 39374 33744 39380
rect 55404 39432 55456 39438
rect 55404 39374 55456 39380
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 26988 39098 27016 39374
rect 34244 39296 34296 39302
rect 34244 39238 34296 39244
rect 26976 39092 27028 39098
rect 26976 39034 27028 39040
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 12808 36168 12860 36174
rect 12808 36110 12860 36116
rect 7208 35866 7328 35894
rect 8864 35866 8984 35894
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 5632 34740 5684 34746
rect 5632 34682 5684 34688
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 5540 33312 5592 33318
rect 5540 33254 5592 33260
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4988 31952 5040 31958
rect 4988 31894 5040 31900
rect 3252 31726 3372 31754
rect 2964 30728 3016 30734
rect 2964 30670 3016 30676
rect 2872 30660 2924 30666
rect 2872 30602 2924 30608
rect 2780 30592 2832 30598
rect 2780 30534 2832 30540
rect 2792 30394 2820 30534
rect 2780 30388 2832 30394
rect 2780 30330 2832 30336
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2700 29510 2728 30194
rect 2688 29504 2740 29510
rect 2688 29446 2740 29452
rect 2884 29209 2912 30602
rect 2976 30433 3004 30670
rect 2962 30424 3018 30433
rect 2962 30359 3018 30368
rect 2964 30184 3016 30190
rect 2964 30126 3016 30132
rect 2976 29714 3004 30126
rect 2964 29708 3016 29714
rect 2964 29650 3016 29656
rect 2870 29200 2926 29209
rect 2870 29135 2926 29144
rect 2596 29028 2648 29034
rect 2596 28970 2648 28976
rect 2872 29028 2924 29034
rect 2872 28970 2924 28976
rect 2504 23248 2556 23254
rect 2504 23190 2556 23196
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2240 22817 2268 23054
rect 2226 22808 2282 22817
rect 2226 22743 2282 22752
rect 2504 22024 2556 22030
rect 2504 21966 2556 21972
rect 2516 21146 2544 21966
rect 2504 21140 2556 21146
rect 2504 21082 2556 21088
rect 2608 19990 2636 28970
rect 2884 28801 2912 28970
rect 2870 28792 2926 28801
rect 2870 28727 2926 28736
rect 3056 28076 3108 28082
rect 3056 28018 3108 28024
rect 2872 27872 2924 27878
rect 3068 27849 3096 28018
rect 2872 27814 2924 27820
rect 3054 27840 3110 27849
rect 2884 27130 2912 27814
rect 3054 27775 3110 27784
rect 2964 27396 3016 27402
rect 2964 27338 3016 27344
rect 2872 27124 2924 27130
rect 2872 27066 2924 27072
rect 2976 26926 3004 27338
rect 3148 27328 3200 27334
rect 3148 27270 3200 27276
rect 3160 27130 3188 27270
rect 3148 27124 3200 27130
rect 3148 27066 3200 27072
rect 2964 26920 3016 26926
rect 2964 26862 3016 26868
rect 3056 26920 3108 26926
rect 3056 26862 3108 26868
rect 3344 26874 3372 31726
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4896 30864 4948 30870
rect 4896 30806 4948 30812
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 4712 30592 4764 30598
rect 4712 30534 4764 30540
rect 4724 30258 4752 30534
rect 4712 30252 4764 30258
rect 4712 30194 4764 30200
rect 4068 30184 4120 30190
rect 4068 30126 4120 30132
rect 3608 30048 3660 30054
rect 3608 29990 3660 29996
rect 3424 29572 3476 29578
rect 3424 29514 3476 29520
rect 3436 29306 3464 29514
rect 3424 29300 3476 29306
rect 3424 29242 3476 29248
rect 3620 29170 3648 29990
rect 4080 29730 4108 30126
rect 4620 30048 4672 30054
rect 4620 29990 4672 29996
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4080 29702 4200 29730
rect 4172 29646 4200 29702
rect 4632 29646 4660 29990
rect 4816 29866 4844 30670
rect 4724 29838 4844 29866
rect 4724 29782 4752 29838
rect 4712 29776 4764 29782
rect 4712 29718 4764 29724
rect 4804 29708 4856 29714
rect 4804 29650 4856 29656
rect 4160 29640 4212 29646
rect 4160 29582 4212 29588
rect 4620 29640 4672 29646
rect 4620 29582 4672 29588
rect 4172 29322 4200 29582
rect 3988 29294 4200 29322
rect 3608 29164 3660 29170
rect 3608 29106 3660 29112
rect 3988 29102 4016 29294
rect 4160 29164 4212 29170
rect 4160 29106 4212 29112
rect 3976 29096 4028 29102
rect 3976 29038 4028 29044
rect 3988 28082 4016 29038
rect 4172 29016 4200 29106
rect 4080 28988 4200 29016
rect 4620 29028 4672 29034
rect 4080 28762 4108 28988
rect 4620 28970 4672 28976
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 4632 28150 4660 28970
rect 4816 28626 4844 29650
rect 4804 28620 4856 28626
rect 4804 28562 4856 28568
rect 4620 28144 4672 28150
rect 4620 28086 4672 28092
rect 3976 28076 4028 28082
rect 3976 28018 4028 28024
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4816 27402 4844 28562
rect 4908 28558 4936 30806
rect 5000 29646 5028 31894
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 5448 29096 5500 29102
rect 5448 29038 5500 29044
rect 4896 28552 4948 28558
rect 4896 28494 4948 28500
rect 4804 27396 4856 27402
rect 4804 27338 4856 27344
rect 3792 27328 3844 27334
rect 3792 27270 3844 27276
rect 3804 27062 3832 27270
rect 3792 27056 3844 27062
rect 3792 26998 3844 27004
rect 3700 26988 3752 26994
rect 3700 26930 3752 26936
rect 3068 26382 3096 26862
rect 3344 26846 3648 26874
rect 3516 26784 3568 26790
rect 3516 26726 3568 26732
rect 3424 26580 3476 26586
rect 3424 26522 3476 26528
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3252 26042 3280 26318
rect 3240 26036 3292 26042
rect 3240 25978 3292 25984
rect 3436 25974 3464 26522
rect 3528 26042 3556 26726
rect 3516 26036 3568 26042
rect 3516 25978 3568 25984
rect 3424 25968 3476 25974
rect 3424 25910 3476 25916
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2700 24274 2728 24550
rect 2688 24268 2740 24274
rect 2688 24210 2740 24216
rect 2884 22642 2912 25638
rect 3240 25152 3292 25158
rect 3240 25094 3292 25100
rect 3148 24812 3200 24818
rect 3148 24754 3200 24760
rect 3056 24268 3108 24274
rect 3056 24210 3108 24216
rect 3068 24018 3096 24210
rect 3160 24177 3188 24754
rect 3252 24614 3280 25094
rect 3436 24750 3464 25910
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 3240 24608 3292 24614
rect 3240 24550 3292 24556
rect 3252 24206 3280 24550
rect 3240 24200 3292 24206
rect 3146 24168 3202 24177
rect 3240 24142 3292 24148
rect 3146 24103 3202 24112
rect 3068 23990 3188 24018
rect 3160 23594 3188 23990
rect 3516 23656 3568 23662
rect 3516 23598 3568 23604
rect 3148 23588 3200 23594
rect 3148 23530 3200 23536
rect 2964 22976 3016 22982
rect 2964 22918 3016 22924
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2792 22166 2820 22578
rect 2780 22160 2832 22166
rect 2780 22102 2832 22108
rect 2688 21888 2740 21894
rect 2688 21830 2740 21836
rect 2700 21622 2728 21830
rect 2688 21616 2740 21622
rect 2688 21558 2740 21564
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 2596 19984 2648 19990
rect 2596 19926 2648 19932
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2608 19446 2636 19654
rect 2596 19440 2648 19446
rect 2596 19382 2648 19388
rect 2700 19378 2728 21286
rect 2976 21010 3004 22918
rect 3160 22574 3188 23530
rect 3528 23322 3556 23598
rect 3620 23526 3648 26846
rect 3712 26625 3740 26930
rect 3698 26616 3754 26625
rect 3698 26551 3754 26560
rect 3700 26512 3752 26518
rect 3700 26454 3752 26460
rect 3712 26246 3740 26454
rect 3700 26240 3752 26246
rect 3700 26182 3752 26188
rect 3804 24818 3832 26998
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4816 25974 4844 27338
rect 5460 26926 5488 29038
rect 5552 28626 5580 33254
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 5644 27538 5672 34682
rect 5724 34536 5776 34542
rect 5724 34478 5776 34484
rect 5632 27532 5684 27538
rect 5632 27474 5684 27480
rect 5736 27402 5764 34478
rect 7300 31754 7328 35866
rect 7208 31726 7328 31754
rect 6828 29844 6880 29850
rect 6828 29786 6880 29792
rect 6840 29510 6868 29786
rect 7012 29640 7064 29646
rect 7012 29582 7064 29588
rect 6828 29504 6880 29510
rect 6828 29446 6880 29452
rect 7024 28422 7052 29582
rect 7012 28416 7064 28422
rect 7012 28358 7064 28364
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6644 27872 6696 27878
rect 6644 27814 6696 27820
rect 5724 27396 5776 27402
rect 5724 27338 5776 27344
rect 6656 27062 6684 27814
rect 6840 27674 6868 28018
rect 7024 27946 7052 28358
rect 7012 27940 7064 27946
rect 7012 27882 7064 27888
rect 6828 27668 6880 27674
rect 6828 27610 6880 27616
rect 7012 27328 7064 27334
rect 7012 27270 7064 27276
rect 7024 27130 7052 27270
rect 7012 27124 7064 27130
rect 7012 27066 7064 27072
rect 6644 27056 6696 27062
rect 6644 26998 6696 27004
rect 5448 26920 5500 26926
rect 5448 26862 5500 26868
rect 5908 26920 5960 26926
rect 5908 26862 5960 26868
rect 4804 25968 4856 25974
rect 4804 25910 4856 25916
rect 4816 25838 4844 25910
rect 5920 25906 5948 26862
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 5908 25900 5960 25906
rect 5908 25842 5960 25848
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 3884 25288 3936 25294
rect 3884 25230 3936 25236
rect 3792 24812 3844 24818
rect 3792 24754 3844 24760
rect 3896 24070 3924 25230
rect 5552 25158 5580 25842
rect 5920 25362 5948 25842
rect 5908 25356 5960 25362
rect 5908 25298 5960 25304
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 4080 24410 4108 24754
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 3884 24064 3936 24070
rect 3804 24024 3884 24052
rect 3608 23520 3660 23526
rect 3608 23462 3660 23468
rect 3516 23316 3568 23322
rect 3516 23258 3568 23264
rect 3804 22642 3832 24024
rect 3884 24006 3936 24012
rect 4080 23866 4108 24346
rect 4160 24132 4212 24138
rect 4160 24074 4212 24080
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4172 23798 4200 24074
rect 5448 24064 5500 24070
rect 5446 24032 5448 24041
rect 5500 24032 5502 24041
rect 5446 23967 5502 23976
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 5552 23730 5580 25094
rect 5632 24880 5684 24886
rect 5632 24822 5684 24828
rect 5644 24206 5672 24822
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 5632 24200 5684 24206
rect 5632 24142 5684 24148
rect 5540 23724 5592 23730
rect 5540 23666 5592 23672
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 4896 22772 4948 22778
rect 4896 22714 4948 22720
rect 3792 22636 3844 22642
rect 3792 22578 3844 22584
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 3148 22568 3200 22574
rect 3148 22510 3200 22516
rect 3160 21010 3188 22510
rect 3804 21350 3832 22578
rect 3896 22234 3924 22578
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3884 22228 3936 22234
rect 3884 22170 3936 22176
rect 3988 22030 4016 22374
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 4908 21622 4936 22714
rect 4896 21616 4948 21622
rect 4896 21558 4948 21564
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3160 20398 3188 20946
rect 4080 20942 4108 21286
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 3148 20392 3200 20398
rect 3148 20334 3200 20340
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2792 19854 2820 20198
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 3712 19514 3740 20402
rect 3896 20369 3924 20402
rect 3882 20360 3938 20369
rect 3882 20295 3938 20304
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 4908 19446 4936 19654
rect 4896 19440 4948 19446
rect 4896 19382 4948 19388
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 2332 18426 2360 18634
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 2516 17746 2544 19246
rect 3974 19136 4030 19145
rect 3974 19071 4030 19080
rect 2688 18964 2740 18970
rect 2688 18906 2740 18912
rect 2700 18426 2728 18906
rect 3988 18766 4016 19071
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 5092 18970 5120 19790
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2596 18284 2648 18290
rect 2596 18226 2648 18232
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2332 17377 2360 17478
rect 2318 17368 2374 17377
rect 2318 17303 2374 17312
rect 2148 16546 2268 16574
rect 2240 15706 2268 16546
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2412 16516 2464 16522
rect 2412 16458 2464 16464
rect 2332 16250 2360 16458
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2424 16182 2452 16458
rect 2608 16182 2636 18226
rect 2792 17270 2820 18226
rect 3436 17785 3464 18226
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 3422 17776 3478 17785
rect 3422 17711 3478 17720
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2700 16250 2728 16390
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2412 16176 2464 16182
rect 2412 16118 2464 16124
rect 2596 16176 2648 16182
rect 2596 16118 2648 16124
rect 2792 16114 2820 17206
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2884 16561 2912 17138
rect 2870 16552 2926 16561
rect 2870 16487 2926 16496
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2780 16108 2832 16114
rect 2832 16068 2912 16096
rect 2780 16050 2832 16056
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 1964 14618 1992 15438
rect 2332 15337 2360 15438
rect 2318 15328 2374 15337
rect 2318 15263 2374 15272
rect 2516 15094 2544 16050
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 2332 14074 2360 14282
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13569 1624 13670
rect 1582 13560 1638 13569
rect 1582 13495 1638 13504
rect 2608 13394 2636 14350
rect 2700 14074 2728 14554
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2792 13977 2820 14962
rect 2778 13968 2834 13977
rect 2884 13938 2912 16068
rect 3804 16046 3832 17614
rect 3884 17604 3936 17610
rect 3884 17546 3936 17552
rect 3896 17338 3924 17546
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4172 17338 4200 17478
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3988 16726 4016 17138
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3804 15502 3832 15982
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 2778 13903 2834 13912
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 3804 13394 3832 15438
rect 4632 15162 4660 16050
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4724 15502 4752 15846
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1582 13288 1638 13297
rect 1412 13161 1440 13262
rect 1582 13223 1638 13232
rect 1596 13190 1624 13223
rect 1584 13184 1636 13190
rect 1398 13152 1454 13161
rect 1584 13126 1636 13132
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 1398 13087 1454 13096
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1872 11937 1900 12786
rect 1858 11928 1914 11937
rect 2148 11898 2176 13126
rect 2608 12170 2636 13330
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2792 12753 2820 13262
rect 3988 12866 4016 13874
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 4080 12986 4108 13194
rect 4632 13190 4660 13806
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4632 12986 4660 13126
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 3988 12850 4384 12866
rect 5276 12850 5304 21286
rect 5644 17610 5672 22918
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 18630 6040 19110
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 5632 17604 5684 17610
rect 5632 17546 5684 17552
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5460 15026 5488 15302
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5460 14618 5488 14962
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 3608 12844 3660 12850
rect 3988 12844 4396 12850
rect 3988 12838 4344 12844
rect 3608 12786 3660 12792
rect 4344 12786 4396 12792
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 2778 12744 2834 12753
rect 2778 12679 2834 12688
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 2884 12345 2912 12582
rect 3240 12368 3292 12374
rect 2870 12336 2926 12345
rect 3240 12310 3292 12316
rect 2870 12271 2926 12280
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 1858 11863 1914 11872
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11121 1624 11494
rect 2608 11218 2636 12106
rect 3252 11762 3280 12310
rect 3436 12238 3464 12582
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 1582 11112 1638 11121
rect 1582 11047 1638 11056
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1872 10713 1900 11018
rect 1858 10704 1914 10713
rect 1584 10668 1636 10674
rect 2056 10674 2084 11154
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 1858 10639 1914 10648
rect 2044 10668 2096 10674
rect 1584 10610 1636 10616
rect 2044 10610 2096 10616
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 9722 1440 10406
rect 1596 10305 1624 10610
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 1400 9716 1452 9722
rect 2056 9674 2084 10610
rect 2148 10266 2176 11086
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2516 10742 2544 10950
rect 2608 10742 2636 11018
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2700 10130 2728 11630
rect 3332 11552 3384 11558
rect 3528 11529 3556 11698
rect 3620 11626 3648 12786
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3332 11494 3384 11500
rect 3514 11520 3570 11529
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 1400 9658 1452 9664
rect 1872 9646 2084 9674
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 1636 9344 1638 9353
rect 1582 9279 1638 9288
rect 1872 9042 1900 9646
rect 2700 9518 2728 10066
rect 3344 10062 3372 11494
rect 3514 11455 3570 11464
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 5460 11354 5488 12582
rect 5644 11830 5672 17546
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5828 17202 5856 17478
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5908 15564 5960 15570
rect 5908 15506 5960 15512
rect 5920 14958 5948 15506
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 6012 12306 6040 18566
rect 6196 15094 6224 24550
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6472 18290 6500 23666
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6184 15088 6236 15094
rect 6184 15030 6236 15036
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5632 11824 5684 11830
rect 5632 11766 5684 11772
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4908 10810 4936 11018
rect 5460 10810 5488 11290
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5736 10674 5764 11494
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10266 3464 10406
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 5092 9722 5120 10610
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8537 1624 8910
rect 1582 8528 1638 8537
rect 1872 8498 1900 8978
rect 2424 8974 2452 9318
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 1582 8463 1638 8472
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1398 8120 1454 8129
rect 1398 8055 1454 8064
rect 1412 7954 1440 8055
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 7313 1532 7346
rect 1490 7304 1546 7313
rect 1490 7239 1546 7248
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 7002 1624 7142
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6497 1440 6734
rect 1398 6488 1454 6497
rect 1398 6423 1454 6432
rect 1584 6112 1636 6118
rect 1582 6080 1584 6089
rect 1636 6080 1638 6089
rect 1582 6015 1638 6024
rect 1872 5794 1900 8434
rect 2056 7546 2084 8774
rect 2240 8566 2268 8774
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2700 8022 2728 9454
rect 3056 8968 3108 8974
rect 3054 8936 3056 8945
rect 3108 8936 3110 8945
rect 3054 8871 3110 8880
rect 3344 8362 3372 9590
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2700 7342 2728 7958
rect 4632 7954 4660 8910
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 2872 7744 2924 7750
rect 2870 7712 2872 7721
rect 2924 7712 2926 7721
rect 2870 7647 2926 7656
rect 4908 7478 4936 9454
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5184 8634 5212 8842
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5736 8498 5764 10610
rect 5920 9178 5948 11698
rect 6012 10062 6040 12242
rect 6380 10130 6408 17478
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8634 5856 8774
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5920 8566 5948 9114
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5276 7546 5304 7754
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 1872 5778 2084 5794
rect 1860 5772 2084 5778
rect 1912 5766 2084 5772
rect 1860 5714 1912 5720
rect 1858 5672 1914 5681
rect 2056 5642 2084 5766
rect 2608 5710 2636 6598
rect 2700 6254 2728 7278
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 2884 6798 2912 7142
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 3344 6458 3372 7142
rect 3528 6905 3556 7346
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3514 6896 3570 6905
rect 3514 6831 3570 6840
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3528 6390 3556 6666
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 1858 5607 1914 5616
rect 2044 5636 2096 5642
rect 1872 5302 1900 5607
rect 2044 5578 2096 5584
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 1860 5296 1912 5302
rect 1860 5238 1912 5244
rect 1584 4752 1636 4758
rect 1584 4694 1636 4700
rect 1124 4480 1176 4486
rect 1124 4422 1176 4428
rect 204 3936 256 3942
rect 204 3878 256 3884
rect 216 800 244 3878
rect 664 3392 716 3398
rect 664 3334 716 3340
rect 676 800 704 3334
rect 1136 800 1164 4422
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1412 1873 1440 2994
rect 1492 2372 1544 2378
rect 1492 2314 1544 2320
rect 1398 1864 1454 1873
rect 1398 1799 1454 1808
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1504 649 1532 2314
rect 1596 800 1624 4694
rect 2056 4162 2084 5578
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2148 4282 2176 4966
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2700 4457 2728 4558
rect 2780 4480 2832 4486
rect 2686 4448 2742 4457
rect 2780 4422 2832 4428
rect 2686 4383 2742 4392
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 2056 4146 2176 4162
rect 2056 4140 2188 4146
rect 2056 4134 2136 4140
rect 1858 3904 1914 3913
rect 1858 3839 1914 3848
rect 1872 3534 1900 3839
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 2056 2650 2084 4134
rect 2136 4082 2188 4088
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2148 800 2176 3674
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2608 800 2636 2790
rect 1490 640 1546 649
rect 1490 575 1546 584
rect 1582 0 1638 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 2792 241 2820 4422
rect 2884 4321 2912 4966
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2870 4312 2926 4321
rect 2870 4247 2926 4256
rect 2976 1465 3004 4558
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3054 2680 3110 2689
rect 3054 2615 3056 2624
rect 3108 2615 3110 2624
rect 3056 2586 3108 2592
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 2962 1456 3018 1465
rect 2962 1391 3018 1400
rect 3068 800 3096 2246
rect 3160 1057 3188 4490
rect 3344 3194 3372 5578
rect 3528 5114 3556 6326
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 3620 5234 3648 6054
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4816 5710 4844 6054
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4172 5234 4200 5646
rect 4908 5574 4936 7414
rect 5552 7342 5580 7686
rect 5736 7410 5764 8434
rect 6012 8090 6040 9386
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6012 7478 6040 8026
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5736 6866 5764 7346
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5736 6322 5764 6802
rect 6288 6798 6316 7822
rect 6472 7342 6500 18226
rect 6748 18154 6776 18770
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6932 18358 6960 18566
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6564 17746 6592 18022
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6748 17678 6776 18090
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6748 17202 6776 17614
rect 6840 17542 6868 18022
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6564 15638 6592 16526
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6748 15570 6776 17138
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6840 16114 6868 16390
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6932 15910 6960 18158
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 7024 15162 7052 27066
rect 7208 25430 7236 31726
rect 7472 29844 7524 29850
rect 7472 29786 7524 29792
rect 7288 29572 7340 29578
rect 7288 29514 7340 29520
rect 7300 29306 7328 29514
rect 7380 29504 7432 29510
rect 7380 29446 7432 29452
rect 7288 29300 7340 29306
rect 7288 29242 7340 29248
rect 7300 28558 7328 29242
rect 7392 29170 7420 29446
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 7288 25764 7340 25770
rect 7288 25706 7340 25712
rect 7196 25424 7248 25430
rect 7196 25366 7248 25372
rect 7208 24750 7236 25366
rect 7300 24954 7328 25706
rect 7288 24948 7340 24954
rect 7288 24890 7340 24896
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 7116 23118 7144 23598
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 7116 20874 7144 23054
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7300 20942 7328 21286
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 7116 20398 7144 20810
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7116 19378 7144 20334
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7116 17882 7144 18702
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7024 14414 7052 15098
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 7208 14346 7236 19450
rect 7484 15026 7512 29786
rect 7932 29640 7984 29646
rect 7932 29582 7984 29588
rect 7944 28762 7972 29582
rect 7932 28756 7984 28762
rect 7932 28698 7984 28704
rect 7564 28620 7616 28626
rect 7564 28562 7616 28568
rect 7576 27538 7604 28562
rect 7656 27940 7708 27946
rect 7656 27882 7708 27888
rect 7564 27532 7616 27538
rect 7564 27474 7616 27480
rect 7668 22094 7696 27882
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 7748 25220 7800 25226
rect 7748 25162 7800 25168
rect 7760 24614 7788 25162
rect 8128 25158 8156 27474
rect 8576 25288 8628 25294
rect 8576 25230 8628 25236
rect 8116 25152 8168 25158
rect 8116 25094 8168 25100
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7668 22066 7788 22094
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7668 21146 7696 21626
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7576 18426 7604 18566
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7656 17264 7708 17270
rect 7656 17206 7708 17212
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 16794 7604 16934
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7484 14906 7512 14962
rect 7392 14878 7512 14906
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6656 13870 6684 14214
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 13530 6960 13670
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6656 12850 6684 13398
rect 7116 12986 7144 13466
rect 7208 13394 7236 14282
rect 7300 14074 7328 14758
rect 7392 14414 7420 14878
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6656 12442 6684 12786
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6748 8362 6776 9998
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6390 5948 6598
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5356 6248 5408 6254
rect 5276 6208 5356 6236
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 3792 5160 3844 5166
rect 3528 5086 3648 5114
rect 3792 5102 3844 5108
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3436 4146 3464 4966
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3528 3534 3556 4966
rect 3620 3942 3648 5086
rect 3804 4729 3832 5102
rect 4816 5030 4844 5170
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 3976 4752 4028 4758
rect 3790 4720 3846 4729
rect 3976 4694 4028 4700
rect 3790 4655 3846 4664
rect 3988 4146 4016 4694
rect 4816 4622 4844 4966
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3620 3346 3648 3878
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3528 3318 3648 3346
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3528 2990 3556 3318
rect 3608 3120 3660 3126
rect 3608 3062 3660 3068
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3146 1048 3202 1057
rect 3146 983 3202 992
rect 3620 800 3648 3062
rect 3712 3058 3740 3402
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3804 2446 3832 3334
rect 3896 3194 3924 3470
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 4080 3097 4108 4014
rect 4632 4010 4660 4422
rect 4724 4146 4752 4422
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4816 3738 4844 4082
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4908 3670 4936 5510
rect 5276 5030 5304 6208
rect 5356 6190 5408 6196
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5460 5914 5488 6122
rect 6288 6118 6316 6734
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5552 5370 5580 5714
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4066 3088 4122 3097
rect 5000 3058 5028 3674
rect 5092 3602 5120 4082
rect 5276 3602 5304 4966
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 4066 3023 4122 3032
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 4080 2281 4108 2858
rect 5368 2774 5396 4490
rect 6288 4010 6684 4026
rect 6276 4004 6684 4010
rect 6328 3998 6684 4004
rect 6276 3946 6328 3952
rect 6656 3942 6684 3998
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6380 3194 6408 3402
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 5368 2746 5488 2774
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 5460 2650 5488 2746
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 6000 2576 6052 2582
rect 6000 2518 6052 2524
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4066 2272 4122 2281
rect 4066 2207 4122 2216
rect 4540 800 4568 2382
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5080 1420 5132 1426
rect 5080 1362 5132 1368
rect 5092 800 5120 1362
rect 5552 800 5580 2246
rect 6012 800 6040 2518
rect 6472 800 6500 2858
rect 6564 2446 6592 3878
rect 6748 3602 6776 8298
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6840 3398 6868 10066
rect 6932 3534 6960 11018
rect 7024 11014 7052 12650
rect 7208 12374 7236 13126
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7300 12238 7328 13738
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7392 12850 7420 12922
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7484 12238 7512 14758
rect 7668 14498 7696 17206
rect 7576 14470 7696 14498
rect 7576 13326 7604 14470
rect 7760 14362 7788 22066
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7852 20058 7880 20402
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 8128 19922 8156 25094
rect 8588 24818 8616 25230
rect 8668 25220 8720 25226
rect 8668 25162 8720 25168
rect 8576 24812 8628 24818
rect 8576 24754 8628 24760
rect 8588 23186 8616 24754
rect 8576 23180 8628 23186
rect 8576 23122 8628 23128
rect 8588 22642 8616 23122
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8220 19718 8248 20470
rect 8312 19854 8340 21558
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8220 18290 8248 19314
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8220 17898 8248 18226
rect 8220 17870 8340 17898
rect 8312 17746 8340 17870
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7852 17338 7880 17546
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8128 15366 8156 15846
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7852 14414 7880 14554
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7668 14334 7788 14362
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7668 13530 7696 14334
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 14006 7788 14214
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7760 13462 7788 13738
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7564 13320 7616 13326
rect 7616 13268 7788 13274
rect 7564 13262 7788 13268
rect 7576 13246 7788 13262
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7576 12850 7604 13126
rect 7760 12986 7788 13246
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7760 12782 7788 12922
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7852 12646 7880 14350
rect 7944 14006 7972 14418
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 8036 13802 8064 14894
rect 8128 14618 8156 15302
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8128 14414 8156 14554
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8496 14346 8524 14826
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8036 13326 8064 13466
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 7944 13190 7972 13262
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7484 11830 7512 12038
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7944 11082 7972 12038
rect 8036 11354 8064 13262
rect 8128 12782 8156 13398
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 8036 10674 8064 11290
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7208 10130 7236 10610
rect 7300 10266 7328 10610
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7208 9518 7236 10066
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7300 9450 7328 10202
rect 7484 9994 7512 10474
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7484 9518 7512 9930
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7484 6662 7512 9454
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7300 4826 7328 5170
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6656 2990 6684 3334
rect 7116 3058 7144 4626
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7484 4146 7512 4422
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7484 4010 7512 4082
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7576 3738 7604 3946
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7484 3058 7512 3470
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 7024 2378 7052 2586
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6656 1426 6684 2246
rect 7576 1850 7604 3470
rect 7668 2922 7696 9998
rect 8220 9586 8248 13942
rect 8390 13288 8446 13297
rect 8390 13223 8392 13232
rect 8444 13223 8446 13232
rect 8392 13194 8444 13200
rect 8496 13190 8524 14282
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8496 12850 8524 13126
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8312 11626 8340 12242
rect 8496 11762 8524 12786
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8588 12306 8616 12582
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8220 9178 8248 9522
rect 8312 9450 8340 11562
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8496 9994 8524 10134
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8496 9450 8524 9930
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7760 7410 7788 7890
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7760 4622 7788 7346
rect 8128 6798 8156 7822
rect 8312 7750 8340 9386
rect 8496 7954 8524 9386
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8220 7478 8248 7686
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8128 5642 8156 6734
rect 8680 5914 8708 25162
rect 8852 24812 8904 24818
rect 8772 24772 8852 24800
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8496 4758 8524 5238
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 8588 4690 8616 5510
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 7760 2854 7788 4558
rect 7852 4078 7880 4558
rect 8588 4298 8616 4626
rect 8666 4448 8722 4457
rect 8666 4383 8722 4392
rect 8496 4270 8616 4298
rect 8496 4146 8524 4270
rect 8680 4214 8708 4383
rect 8668 4208 8720 4214
rect 8668 4150 8720 4156
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 8220 3738 8248 4082
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7484 1822 7604 1850
rect 6644 1420 6696 1426
rect 6644 1362 6696 1368
rect 7484 800 7512 1822
rect 7944 800 7972 2926
rect 8772 2774 8800 24772
rect 8852 24754 8904 24760
rect 8956 23866 8984 35866
rect 10876 32904 10928 32910
rect 10876 32846 10928 32852
rect 10888 28558 10916 32846
rect 10876 28552 10928 28558
rect 10876 28494 10928 28500
rect 10968 28552 11020 28558
rect 10968 28494 11020 28500
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 10508 28416 10560 28422
rect 10508 28358 10560 28364
rect 10520 28150 10548 28358
rect 10508 28144 10560 28150
rect 10508 28086 10560 28092
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 9692 27674 9720 28018
rect 10888 27946 10916 28494
rect 10876 27940 10928 27946
rect 10876 27882 10928 27888
rect 9680 27668 9732 27674
rect 9680 27610 9732 27616
rect 9692 27538 9720 27610
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 9312 26036 9364 26042
rect 9312 25978 9364 25984
rect 9324 25294 9352 25978
rect 9692 25974 9720 27474
rect 10980 27402 11008 28494
rect 12544 28082 12572 28494
rect 12532 28076 12584 28082
rect 12532 28018 12584 28024
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12544 27962 12572 28018
rect 12544 27934 12664 27962
rect 12636 27674 12664 27934
rect 12728 27674 12756 28018
rect 12624 27668 12676 27674
rect 12624 27610 12676 27616
rect 12716 27668 12768 27674
rect 12716 27610 12768 27616
rect 10508 27396 10560 27402
rect 10508 27338 10560 27344
rect 10968 27396 11020 27402
rect 10968 27338 11020 27344
rect 10520 27130 10548 27338
rect 10876 27328 10928 27334
rect 10876 27270 10928 27276
rect 10888 27130 10916 27270
rect 10508 27124 10560 27130
rect 10508 27066 10560 27072
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 10980 26994 11008 27338
rect 10692 26988 10744 26994
rect 10692 26930 10744 26936
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10704 26790 10732 26930
rect 10692 26784 10744 26790
rect 10692 26726 10744 26732
rect 9680 25968 9732 25974
rect 9680 25910 9732 25916
rect 12636 25906 12664 27610
rect 12820 26042 12848 36110
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 13820 33992 13872 33998
rect 13820 33934 13872 33940
rect 13452 28484 13504 28490
rect 13452 28426 13504 28432
rect 12900 27396 12952 27402
rect 12900 27338 12952 27344
rect 12808 26036 12860 26042
rect 12808 25978 12860 25984
rect 9496 25900 9548 25906
rect 9496 25842 9548 25848
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 9508 25498 9536 25842
rect 10888 25498 10916 25842
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 10876 25492 10928 25498
rect 10876 25434 10928 25440
rect 10980 25430 11008 25638
rect 10968 25424 11020 25430
rect 10968 25366 11020 25372
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 10416 25288 10468 25294
rect 10416 25230 10468 25236
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 12072 25288 12124 25294
rect 12532 25288 12584 25294
rect 12072 25230 12124 25236
rect 12452 25248 12532 25276
rect 9036 25152 9088 25158
rect 9036 25094 9088 25100
rect 9048 24886 9076 25094
rect 9036 24880 9088 24886
rect 9036 24822 9088 24828
rect 9692 24818 9720 25230
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 8956 23662 8984 23802
rect 9312 23724 9364 23730
rect 9312 23666 9364 23672
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 8944 23656 8996 23662
rect 8944 23598 8996 23604
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 9048 22642 9076 23258
rect 9324 23186 9352 23666
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 9312 23044 9364 23050
rect 9312 22986 9364 22992
rect 9220 22976 9272 22982
rect 9220 22918 9272 22924
rect 9232 22642 9260 22918
rect 9324 22778 9352 22986
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 8864 12434 8892 22578
rect 9416 22094 9444 23666
rect 9600 23050 9628 23666
rect 9588 23044 9640 23050
rect 9588 22986 9640 22992
rect 9600 22574 9628 22986
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9324 22066 9444 22094
rect 10428 22094 10456 25230
rect 10704 24818 10732 25230
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10704 23730 10732 24754
rect 10796 23798 10824 24754
rect 12084 24682 12112 25230
rect 12072 24676 12124 24682
rect 12072 24618 12124 24624
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 10784 23792 10836 23798
rect 10784 23734 10836 23740
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10796 23118 10824 23734
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 10968 23588 11020 23594
rect 10968 23530 11020 23536
rect 10980 23186 11008 23530
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11716 23202 11744 23462
rect 11808 23322 11836 23666
rect 11796 23316 11848 23322
rect 11796 23258 11848 23264
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 11624 23174 11744 23202
rect 11624 23118 11652 23174
rect 11900 23118 11928 24006
rect 10784 23112 10836 23118
rect 11244 23112 11296 23118
rect 10836 23060 11008 23066
rect 10784 23054 11008 23060
rect 11244 23054 11296 23060
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11888 23112 11940 23118
rect 11888 23054 11940 23060
rect 10796 23038 11008 23054
rect 10876 22160 10928 22166
rect 10876 22102 10928 22108
rect 10428 22066 10548 22094
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8956 17882 8984 21422
rect 8944 17876 8996 17882
rect 8944 17818 8996 17824
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8956 16114 8984 17682
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8864 12406 8984 12434
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8864 7886 8892 8910
rect 8956 8294 8984 12406
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8864 6186 8892 7822
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8864 5370 8892 6122
rect 9140 6118 9168 6666
rect 9232 6186 9260 7278
rect 9220 6180 9272 6186
rect 9220 6122 9272 6128
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 8956 5710 8984 6054
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8956 4622 8984 4966
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8956 2990 8984 4558
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8680 2746 8800 2774
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8496 800 8524 2246
rect 8680 1630 8708 2746
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 8956 1970 8984 2382
rect 8944 1964 8996 1970
rect 8944 1906 8996 1912
rect 9140 1902 9168 5850
rect 9232 3942 9260 6122
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9128 1896 9180 1902
rect 9128 1838 9180 1844
rect 8668 1624 8720 1630
rect 8668 1566 8720 1572
rect 8956 870 9076 898
rect 8956 800 8984 870
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9048 762 9076 870
rect 9232 762 9260 2246
rect 9324 1562 9352 22066
rect 10140 21548 10192 21554
rect 10140 21490 10192 21496
rect 9496 21480 9548 21486
rect 9496 21422 9548 21428
rect 9508 19378 9536 21422
rect 10152 21146 10180 21490
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9692 18766 9720 19654
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9496 16108 9548 16114
rect 9784 16096 9812 19654
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9876 18902 9904 19314
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10336 17270 10364 17478
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9496 16050 9548 16056
rect 9692 16068 9812 16096
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9416 11082 9444 11630
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 9178 9444 11018
rect 9508 10470 9536 16050
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9600 12306 9628 12650
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 4146 9444 8230
rect 9692 7818 9720 16068
rect 9968 14278 9996 16662
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9784 14006 9812 14214
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9968 13462 9996 13738
rect 10060 13530 10088 13874
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 10152 13326 10180 13670
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9784 12714 9812 13194
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 10244 12238 10272 13466
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 11150 9996 11494
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7342 9536 7686
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9600 6798 9628 7210
rect 9784 6798 9812 9998
rect 9968 9586 9996 11086
rect 10060 10266 10088 11698
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10152 10742 10180 10950
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10244 10266 10272 11086
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 8974 9904 9318
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9784 5710 9812 6734
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9692 5234 9720 5510
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9876 4078 9904 8910
rect 9968 4214 9996 9522
rect 10336 9178 10364 15302
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10428 12986 10456 13194
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10060 8906 10088 9114
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10060 8090 10088 8842
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10060 7886 10088 8026
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10060 4826 10088 7822
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7410 10272 7686
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10428 7206 10456 7346
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9876 3602 9904 4014
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 10244 3534 10272 6598
rect 10428 6322 10456 7142
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9876 3126 9904 3334
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9416 800 9444 2518
rect 9508 2446 9536 2790
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 10428 800 10456 4082
rect 10520 2774 10548 22066
rect 10888 21690 10916 22102
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 10600 21616 10652 21622
rect 10600 21558 10652 21564
rect 10612 20942 10640 21558
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10888 20874 10916 21626
rect 10876 20868 10928 20874
rect 10876 20810 10928 20816
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10612 15638 10640 16050
rect 10600 15632 10652 15638
rect 10600 15574 10652 15580
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10612 13870 10640 14418
rect 10704 13938 10732 16934
rect 10980 16590 11008 23038
rect 11256 21962 11284 23054
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 15502 10916 16390
rect 10980 16114 11008 16526
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10612 12646 10640 13398
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10612 9654 10640 10474
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10704 4690 10732 13194
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10796 12374 10824 12854
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10888 11762 10916 12718
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10888 11218 10916 11698
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10980 10554 11008 15846
rect 11072 15502 11100 15846
rect 11164 15502 11192 20742
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11256 19718 11284 19790
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12238 11100 12582
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10888 10526 11008 10554
rect 10888 5166 10916 10526
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 7954 11008 10406
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9518 11100 9862
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10980 6322 11008 7890
rect 11164 6662 11192 15438
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11256 12646 11284 12786
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 5710 11008 6258
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11164 5370 11192 5578
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10612 3534 10640 4422
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10612 2922 10640 3470
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 10704 2854 10732 3470
rect 11164 3398 11192 3674
rect 11348 3602 11376 23054
rect 11428 22976 11480 22982
rect 11796 22976 11848 22982
rect 11480 22924 11796 22930
rect 11428 22918 11848 22924
rect 11440 22902 11836 22918
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11532 20942 11560 21966
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11532 19922 11560 20878
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11440 19514 11468 19858
rect 11624 19786 11652 21286
rect 12084 20806 12112 24618
rect 12452 22930 12480 25248
rect 12532 25230 12584 25236
rect 12636 25106 12664 25842
rect 12820 25294 12848 25978
rect 12912 25294 12940 27338
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 13096 25498 13124 25842
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 12900 25152 12952 25158
rect 12636 25078 12848 25106
rect 12900 25094 12952 25100
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12532 24744 12584 24750
rect 12728 24698 12756 24754
rect 12584 24692 12756 24698
rect 12532 24686 12756 24692
rect 12544 24670 12756 24686
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 12544 23050 12572 24142
rect 12532 23044 12584 23050
rect 12532 22986 12584 22992
rect 12452 22902 12572 22930
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12452 22114 12480 22714
rect 12360 22086 12480 22114
rect 12072 20800 12124 20806
rect 12072 20742 12124 20748
rect 12360 20466 12388 22086
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11440 17678 11468 18702
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11440 16658 11468 17614
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11900 15638 11928 16050
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 11612 15428 11664 15434
rect 11612 15370 11664 15376
rect 11624 15094 11652 15370
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 12084 14958 12112 19450
rect 12176 18766 12204 20402
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12544 17678 12572 22902
rect 12636 22094 12664 24670
rect 12820 24562 12848 25078
rect 12912 24818 12940 25094
rect 13188 24886 13216 25230
rect 13176 24880 13228 24886
rect 13176 24822 13228 24828
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12728 24534 12848 24562
rect 12728 23866 12756 24534
rect 12912 24274 12940 24754
rect 12900 24268 12952 24274
rect 12900 24210 12952 24216
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12728 23186 12756 23802
rect 12716 23180 12768 23186
rect 12716 23122 12768 23128
rect 12728 22778 12756 23122
rect 13268 23044 13320 23050
rect 13268 22986 13320 22992
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12636 22066 12756 22094
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12636 18426 12664 18634
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12176 16658 12296 16674
rect 12164 16652 12296 16658
rect 12216 16646 12296 16652
rect 12164 16594 12216 16600
rect 12072 14952 12124 14958
rect 11992 14900 12072 14906
rect 11992 14894 12124 14900
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 11992 14878 12112 14894
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11440 13394 11468 13806
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11532 12850 11560 13126
rect 11808 12850 11836 13262
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11440 11898 11468 12174
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11532 11150 11560 11834
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11808 10674 11836 11018
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11532 10266 11560 10542
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11900 6866 11928 14826
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11992 5914 12020 14878
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 12084 14006 12112 14758
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12176 12434 12204 13806
rect 12268 13326 12296 16646
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12452 16250 12480 16458
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12544 15162 12572 16050
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12176 12406 12296 12434
rect 12268 11762 12296 12406
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12452 11830 12480 12174
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12636 11830 12664 12038
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12268 11150 12296 11698
rect 12452 11354 12480 11766
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12176 9926 12204 10610
rect 12268 10606 12296 11086
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7478 12296 7822
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12360 5914 12388 10474
rect 12452 9586 12480 11290
rect 12544 10713 12572 11494
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12636 11150 12664 11222
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12530 10704 12586 10713
rect 12530 10639 12586 10648
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12452 7750 12480 9522
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12544 7426 12572 9590
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12636 7546 12664 7754
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12452 7398 12572 7426
rect 12452 7342 12480 7398
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11900 4622 11928 5646
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11900 4146 11928 4558
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11808 3738 11836 4014
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11900 3534 11928 4082
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12084 3602 12112 3674
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11256 3126 11284 3402
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10520 2746 10640 2774
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10520 2106 10548 2382
rect 10508 2100 10560 2106
rect 10508 2042 10560 2048
rect 10612 1698 10640 2746
rect 10600 1692 10652 1698
rect 10600 1634 10652 1640
rect 10888 800 10916 3062
rect 11716 3058 11744 3334
rect 12176 3126 12204 3334
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12084 2446 12112 2790
rect 12728 2774 12756 22066
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 13096 20534 13124 20742
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12820 17270 12848 19314
rect 13188 18970 13216 20946
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 13096 18737 13124 18906
rect 13082 18728 13138 18737
rect 13082 18663 13138 18672
rect 13280 18630 13308 22986
rect 13464 21078 13492 28426
rect 13832 28218 13860 33934
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 25320 31136 25372 31142
rect 25320 31078 25372 31084
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 15108 29708 15160 29714
rect 15108 29650 15160 29656
rect 15120 28762 15148 29650
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 17408 29232 17460 29238
rect 17408 29174 17460 29180
rect 15108 28756 15160 28762
rect 15108 28698 15160 28704
rect 14648 28484 14700 28490
rect 14648 28426 14700 28432
rect 14660 28218 14688 28426
rect 15120 28218 15148 28698
rect 17040 28484 17092 28490
rect 17040 28426 17092 28432
rect 17052 28218 17080 28426
rect 17420 28422 17448 29174
rect 17408 28416 17460 28422
rect 17408 28358 17460 28364
rect 17420 28218 17448 28358
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 13820 28212 13872 28218
rect 13820 28154 13872 28160
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 15108 28212 15160 28218
rect 15108 28154 15160 28160
rect 17040 28212 17092 28218
rect 17040 28154 17092 28160
rect 17408 28212 17460 28218
rect 17408 28154 17460 28160
rect 13832 27402 13860 28154
rect 16948 28076 17000 28082
rect 16948 28018 17000 28024
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 16764 28008 16816 28014
rect 16764 27950 16816 27956
rect 13912 27532 13964 27538
rect 13912 27474 13964 27480
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 13636 26240 13688 26246
rect 13636 26182 13688 26188
rect 13648 25974 13676 26182
rect 13636 25968 13688 25974
rect 13636 25910 13688 25916
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 13360 20936 13412 20942
rect 13358 20904 13360 20913
rect 13544 20936 13596 20942
rect 13412 20904 13414 20913
rect 13544 20878 13596 20884
rect 13358 20839 13414 20848
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13464 20602 13492 20742
rect 13452 20596 13504 20602
rect 13452 20538 13504 20544
rect 13556 19922 13584 20878
rect 13648 20874 13676 22578
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13004 18358 13032 18566
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 13556 18290 13584 19858
rect 13740 19378 13768 26726
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13832 24682 13860 25842
rect 13820 24676 13872 24682
rect 13820 24618 13872 24624
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13832 22982 13860 24074
rect 13820 22976 13872 22982
rect 13820 22918 13872 22924
rect 13832 22710 13860 22918
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13832 19310 13860 21490
rect 13924 19514 13952 27474
rect 16580 27056 16632 27062
rect 16580 26998 16632 27004
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 15108 26308 15160 26314
rect 15108 26250 15160 26256
rect 15120 23798 15148 26250
rect 15752 25696 15804 25702
rect 15752 25638 15804 25644
rect 15764 24750 15792 25638
rect 15752 24744 15804 24750
rect 15752 24686 15804 24692
rect 15200 24676 15252 24682
rect 15200 24618 15252 24624
rect 15212 24206 15240 24618
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 15212 23322 15240 24142
rect 15752 24132 15804 24138
rect 15752 24074 15804 24080
rect 15764 23866 15792 24074
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15200 23316 15252 23322
rect 15200 23258 15252 23264
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 14188 23044 14240 23050
rect 14188 22986 14240 22992
rect 14200 22778 14228 22986
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14476 22778 14504 22918
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 15660 22092 15712 22098
rect 15660 22034 15712 22040
rect 14186 21992 14242 22001
rect 14186 21927 14242 21936
rect 14200 21350 14228 21927
rect 15672 21622 15700 22034
rect 15660 21616 15712 21622
rect 15660 21558 15712 21564
rect 15764 21554 15792 23122
rect 15856 22098 15884 26930
rect 16592 26586 16620 26998
rect 16672 26784 16724 26790
rect 16672 26726 16724 26732
rect 16580 26580 16632 26586
rect 16580 26522 16632 26528
rect 16684 26382 16712 26726
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16028 24064 16080 24070
rect 16028 24006 16080 24012
rect 16040 23798 16068 24006
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 16028 23792 16080 23798
rect 16028 23734 16080 23740
rect 15936 22976 15988 22982
rect 15936 22918 15988 22924
rect 15948 22098 15976 22918
rect 16132 22642 16160 23802
rect 16776 23610 16804 27950
rect 16960 26994 16988 28018
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 17132 25288 17184 25294
rect 17132 25230 17184 25236
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16960 24886 16988 25094
rect 16948 24880 17000 24886
rect 16948 24822 17000 24828
rect 16776 23582 16896 23610
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16028 22568 16080 22574
rect 16028 22510 16080 22516
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15936 22092 15988 22098
rect 15936 22034 15988 22040
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 14188 21344 14240 21350
rect 14188 21286 14240 21292
rect 14384 20942 14412 21490
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14554 20904 14610 20913
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 13912 19508 13964 19514
rect 13912 19450 13964 19456
rect 14200 19310 14228 20742
rect 14292 20466 14320 20878
rect 14554 20839 14610 20848
rect 14568 20806 14596 20839
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14660 20602 14688 20946
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15304 20602 15332 20878
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15304 19922 15332 20402
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14476 19514 14504 19790
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14476 19310 14504 19450
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 13832 18290 13860 19246
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12820 12238 12848 12582
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12820 10470 12848 10746
rect 12912 10674 12940 11018
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 3058 12848 4422
rect 12900 3460 12952 3466
rect 12900 3402 12952 3408
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 12912 2922 12940 3402
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 13004 2774 13032 17614
rect 13096 12102 13124 18226
rect 14292 17814 14320 19110
rect 14844 18290 14872 19790
rect 15580 19514 15608 20878
rect 15764 20398 15792 21490
rect 15948 21350 15976 21898
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 15948 20466 15976 20810
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15764 19378 15792 19654
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14280 17808 14332 17814
rect 14280 17750 14332 17756
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13280 14958 13308 15438
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13096 9110 13124 11562
rect 13188 11286 13216 11698
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 13188 9518 13216 11222
rect 13280 10810 13308 14894
rect 13372 11694 13400 17546
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13464 11370 13492 17614
rect 14372 17264 14424 17270
rect 14372 17206 14424 17212
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14292 16794 14320 17070
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14108 14618 14136 14962
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13372 11342 13492 11370
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13266 10704 13322 10713
rect 13266 10639 13322 10648
rect 13280 10606 13308 10639
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13268 10260 13320 10266
rect 13372 10248 13400 11342
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13464 10674 13492 11154
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13320 10220 13400 10248
rect 13268 10202 13320 10208
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 13280 9042 13308 10202
rect 13360 10056 13412 10062
rect 13464 10044 13492 10610
rect 13412 10016 13492 10044
rect 13360 9998 13412 10004
rect 13372 9586 13400 9998
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13464 9110 13492 9862
rect 13556 9178 13584 14350
rect 14292 14006 14320 16730
rect 14384 16454 14412 17206
rect 14844 17134 14872 18226
rect 14936 17490 14964 18770
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 15028 18086 15056 18634
rect 15212 18426 15240 19314
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15304 18834 15332 19246
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15304 18426 15332 18634
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15028 17610 15056 18022
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 15120 17490 15148 18022
rect 15304 17542 15332 18362
rect 14936 17462 15148 17490
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14200 12986 14228 13194
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12434 13860 12786
rect 13832 12406 13952 12434
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13096 8090 13124 8910
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13096 7546 13124 8026
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 12544 2746 12756 2774
rect 12912 2746 13032 2774
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11348 800 11376 2246
rect 11900 800 11928 2246
rect 12360 800 12388 2518
rect 12544 1834 12572 2746
rect 12532 1828 12584 1834
rect 12532 1770 12584 1776
rect 12912 1766 12940 2746
rect 13280 2650 13308 8842
rect 13464 4078 13492 9046
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 8566 13584 8910
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13648 7410 13676 12038
rect 13740 11558 13768 12106
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10470 13768 11086
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10130 13768 10406
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13740 8634 13768 9114
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13924 8022 13952 12406
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14108 10062 14136 11086
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14096 9444 14148 9450
rect 14096 9386 14148 9392
rect 14108 8906 14136 9386
rect 14096 8900 14148 8906
rect 14096 8842 14148 8848
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 14096 7812 14148 7818
rect 14096 7754 14148 7760
rect 14108 7546 14136 7754
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13648 5166 13676 7346
rect 14200 7002 14228 8026
rect 14292 7818 14320 11494
rect 14384 11354 14412 16390
rect 14568 16182 14596 16390
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14476 15638 14504 16118
rect 14464 15632 14516 15638
rect 14464 15574 14516 15580
rect 14556 14544 14608 14550
rect 14554 14512 14556 14521
rect 14608 14512 14610 14521
rect 14554 14447 14610 14456
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14568 14074 14596 14350
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14568 13190 14596 13874
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 12986 14596 13126
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14752 12238 14780 13670
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14752 10742 14780 12174
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14936 9654 14964 17462
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 15028 16522 15056 17070
rect 15396 16522 15424 19246
rect 15948 18970 15976 20402
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15488 18426 15516 18906
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15672 18222 15700 18906
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15856 18698 15884 18838
rect 15844 18692 15896 18698
rect 15844 18634 15896 18640
rect 16040 18630 16068 22510
rect 16304 22160 16356 22166
rect 16304 22102 16356 22108
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16224 21593 16252 21966
rect 16210 21584 16266 21593
rect 16210 21519 16266 21528
rect 16316 20602 16344 22102
rect 16580 22092 16632 22098
rect 16580 22034 16632 22040
rect 16592 21350 16620 22034
rect 16868 21690 16896 23582
rect 17040 22024 17092 22030
rect 17038 21992 17040 22001
rect 17092 21992 17094 22001
rect 17038 21927 17094 21936
rect 16856 21684 16908 21690
rect 16856 21626 16908 21632
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16316 19310 16344 19790
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16132 18766 16160 18906
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16316 18698 16344 19246
rect 16408 19174 16436 21286
rect 16488 21072 16540 21078
rect 16488 21014 16540 21020
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15934 17776 15990 17785
rect 15934 17711 15990 17720
rect 15948 17678 15976 17711
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 15212 15366 15240 16458
rect 15764 15502 15792 16458
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 14936 9450 14964 9590
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14476 7342 14504 7686
rect 14568 7478 14596 7686
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14476 6798 14504 7278
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14108 6390 14136 6598
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13832 4690 13860 6258
rect 14476 6118 14504 6598
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5778 14504 6054
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14844 5370 14872 8774
rect 15028 8430 15056 8774
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 15120 6866 15148 12786
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15212 7426 15240 12310
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15580 11830 15608 12106
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15672 11286 15700 11630
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15764 11132 15792 15438
rect 15856 14498 15884 17478
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15948 16522 15976 17070
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 16040 15910 16068 18158
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 16132 16658 16160 17206
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16040 14618 16068 15846
rect 16132 15162 16160 16594
rect 16316 16454 16344 18634
rect 16408 17746 16436 18634
rect 16500 17746 16528 21014
rect 16592 21010 16620 21286
rect 17144 21078 17172 25230
rect 17236 22778 17264 28018
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 17316 26920 17368 26926
rect 17316 26862 17368 26868
rect 17328 25226 17356 26862
rect 17408 26308 17460 26314
rect 17408 26250 17460 26256
rect 17420 26042 17448 26250
rect 17408 26036 17460 26042
rect 17408 25978 17460 25984
rect 17788 25906 17816 26930
rect 17972 26568 18000 27814
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 24492 26852 24544 26858
rect 24492 26794 24544 26800
rect 18052 26580 18104 26586
rect 17972 26540 18052 26568
rect 17972 26042 18000 26540
rect 18052 26522 18104 26528
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 17960 26036 18012 26042
rect 17960 25978 18012 25984
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17788 25294 17816 25842
rect 19248 25832 19300 25838
rect 19248 25774 19300 25780
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17776 25288 17828 25294
rect 17776 25230 17828 25236
rect 17316 25220 17368 25226
rect 17316 25162 17368 25168
rect 17328 24614 17356 25162
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17420 24206 17448 25230
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17408 23656 17460 23662
rect 17408 23598 17460 23604
rect 17316 23112 17368 23118
rect 17316 23054 17368 23060
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17224 22432 17276 22438
rect 17224 22374 17276 22380
rect 17236 22098 17264 22374
rect 17328 22234 17356 23054
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17236 21554 17264 21830
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17236 21146 17264 21354
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 16592 19922 16620 20946
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16580 18148 16632 18154
rect 16580 18090 16632 18096
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16408 16114 16436 17682
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16500 17338 16528 17478
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16592 16046 16620 18090
rect 16684 18034 16712 19926
rect 16960 19786 16988 20334
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16868 18290 16896 18702
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16684 18006 16804 18034
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16684 17338 16712 17818
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16670 16824 16726 16833
rect 16670 16759 16672 16768
rect 16724 16759 16726 16768
rect 16672 16730 16724 16736
rect 16672 16448 16724 16454
rect 16776 16436 16804 18006
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 16868 17678 16896 17818
rect 16960 17678 16988 19722
rect 17420 19514 17448 23598
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17512 22438 17540 22986
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 17500 22432 17552 22438
rect 17500 22374 17552 22380
rect 17604 21593 17632 22578
rect 17590 21584 17646 21593
rect 17590 21519 17646 21528
rect 17604 21486 17632 21519
rect 17592 21480 17644 21486
rect 17512 21440 17592 21468
rect 17512 20466 17540 21440
rect 17592 21422 17644 21428
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17512 18698 17540 19790
rect 17604 19310 17632 20946
rect 17696 19990 17724 22578
rect 17776 22568 17828 22574
rect 17960 22568 18012 22574
rect 17776 22510 17828 22516
rect 17880 22528 17960 22556
rect 17788 22234 17816 22510
rect 17776 22228 17828 22234
rect 17776 22170 17828 22176
rect 17880 21350 17908 22528
rect 17960 22510 18012 22516
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 18248 22030 18276 22374
rect 18524 22066 18736 22094
rect 18052 22024 18104 22030
rect 18050 21992 18052 22001
rect 18236 22024 18288 22030
rect 18104 21992 18106 22001
rect 18106 21950 18184 21978
rect 18236 21966 18288 21972
rect 18050 21927 18106 21936
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17880 21078 17908 21286
rect 17972 21146 18000 21490
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17972 20602 18000 20878
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17684 19984 17736 19990
rect 17684 19926 17736 19932
rect 18064 19922 18092 21558
rect 18156 21554 18184 21950
rect 18524 21554 18552 22066
rect 18708 22030 18736 22066
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18616 21486 18644 21966
rect 18880 21616 18932 21622
rect 18880 21558 18932 21564
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18248 20466 18276 20878
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18340 20058 18368 21422
rect 18616 20330 18644 21422
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 18708 20602 18736 21082
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18892 20466 18920 21558
rect 19260 21146 19288 25774
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 21640 24948 21692 24954
rect 21640 24890 21692 24896
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19996 22166 20024 23054
rect 20812 23044 20864 23050
rect 20812 22986 20864 22992
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 20364 22710 20392 22918
rect 20824 22778 20852 22986
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19352 20942 19380 21082
rect 19444 21010 19472 21286
rect 19800 21072 19852 21078
rect 19536 21032 19800 21060
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 19536 20942 19564 21032
rect 19800 21014 19852 21020
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19996 20466 20024 22102
rect 20364 22098 20392 22646
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 21180 21480 21232 21486
rect 21284 21468 21312 22578
rect 21232 21440 21312 21468
rect 21180 21422 21232 21428
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 19984 20460 20036 20466
rect 20720 20460 20772 20466
rect 20036 20420 20208 20448
rect 19984 20402 20036 20408
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18604 20324 18656 20330
rect 18604 20266 18656 20272
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 18616 19854 18644 20266
rect 18708 20058 18736 20334
rect 18984 20262 19012 20334
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 17592 19304 17644 19310
rect 18512 19304 18564 19310
rect 17592 19246 17644 19252
rect 18432 19264 18512 19292
rect 17604 19009 17632 19246
rect 17590 19000 17646 19009
rect 17590 18935 17646 18944
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16868 16658 16896 16934
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16724 16408 16804 16436
rect 16672 16390 16724 16396
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 15856 14470 16160 14498
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 15844 12436 15896 12442
rect 16040 12434 16068 12650
rect 15844 12378 15896 12384
rect 15948 12406 16068 12434
rect 15672 11104 15792 11132
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10810 15608 10950
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15580 8566 15608 9318
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15304 7886 15332 8366
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15488 7546 15516 7822
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15212 7398 15332 7426
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15212 6934 15240 7278
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15120 5846 15148 6802
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15212 5710 15240 6870
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14844 5234 14872 5306
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 14660 4622 14688 4966
rect 15028 4826 15056 5170
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 13910 4176 13966 4185
rect 13910 4111 13966 4120
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13004 2038 13032 2382
rect 12992 2032 13044 2038
rect 12992 1974 13044 1980
rect 12900 1760 12952 1766
rect 12900 1702 12952 1708
rect 13372 800 13400 3470
rect 13464 3233 13492 3878
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13450 3224 13506 3233
rect 13450 3159 13506 3168
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13740 2310 13768 2450
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13832 800 13860 3334
rect 13924 3058 13952 4111
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 14016 3466 14044 3878
rect 15028 3534 15056 4762
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 14004 3460 14056 3466
rect 14004 3402 14056 3408
rect 14832 3460 14884 3466
rect 14884 3420 14964 3448
rect 14832 3402 14884 3408
rect 14556 3392 14608 3398
rect 14462 3360 14518 3369
rect 14556 3334 14608 3340
rect 14462 3295 14518 3304
rect 14476 3126 14504 3295
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14568 3058 14596 3334
rect 14936 3126 14964 3420
rect 15014 3224 15070 3233
rect 15014 3159 15070 3168
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14568 2446 14596 2994
rect 14738 2952 14794 2961
rect 14738 2887 14740 2896
rect 14792 2887 14794 2896
rect 14832 2916 14884 2922
rect 14740 2858 14792 2864
rect 14832 2858 14884 2864
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14292 800 14320 2246
rect 14844 800 14872 2858
rect 14936 2446 14964 3062
rect 15028 3058 15056 3159
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15016 2440 15068 2446
rect 15120 2428 15148 3606
rect 15212 3466 15240 4014
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 15304 3058 15332 7398
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15396 6322 15424 6598
rect 15580 6338 15608 7822
rect 15672 6866 15700 11104
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15764 10266 15792 10542
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15856 10062 15884 12378
rect 15948 12238 15976 12406
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 16040 11830 16068 12242
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15948 11286 15976 11698
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15948 9908 15976 10542
rect 15856 9880 15976 9908
rect 15856 9518 15884 9880
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15764 8430 15792 8910
rect 15856 8906 15884 9454
rect 15948 8974 15976 9454
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15844 8900 15896 8906
rect 15844 8842 15896 8848
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15764 7886 15792 8366
rect 15856 7936 15884 8842
rect 15936 7948 15988 7954
rect 15856 7908 15936 7936
rect 15936 7890 15988 7896
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15672 6458 15700 6802
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15488 6310 15608 6338
rect 15764 6322 15792 7822
rect 15948 6798 15976 7890
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15948 6322 15976 6734
rect 15752 6316 15804 6322
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15200 2848 15252 2854
rect 15252 2808 15332 2836
rect 15200 2790 15252 2796
rect 15068 2400 15148 2428
rect 15016 2382 15068 2388
rect 15304 800 15332 2808
rect 15488 2774 15516 6310
rect 15752 6258 15804 6264
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15580 3670 15608 6190
rect 16132 4690 16160 14470
rect 16408 12442 16436 15030
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16500 14074 16528 14350
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16316 10010 16344 12174
rect 16408 11218 16436 12242
rect 16592 12102 16620 15982
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16684 13870 16712 14758
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 14006 16804 14214
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 16776 12434 16804 13738
rect 16684 12406 16804 12434
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16500 10606 16528 11018
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16500 10062 16528 10542
rect 16224 9982 16344 10010
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16224 7750 16252 9982
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 8974 16344 9862
rect 16592 9466 16620 12038
rect 16684 11694 16712 12406
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16776 10674 16804 11698
rect 16868 11354 16896 13806
rect 16960 13802 16988 17614
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17144 16658 17172 17138
rect 17512 16658 17540 18634
rect 17604 18222 17632 18935
rect 18142 18864 18198 18873
rect 18142 18799 18198 18808
rect 18156 18766 18184 18799
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18156 18290 18184 18702
rect 18234 18456 18290 18465
rect 18234 18391 18236 18400
rect 18288 18391 18290 18400
rect 18236 18362 18288 18368
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 17592 18216 17644 18222
rect 17592 18158 17644 18164
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 18142 18184 18198 18193
rect 17604 17134 17632 18158
rect 17696 17746 17724 18158
rect 18142 18119 18198 18128
rect 18156 18086 18184 18119
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 17774 17776 17830 17785
rect 17684 17740 17736 17746
rect 17774 17711 17776 17720
rect 17684 17682 17736 17688
rect 17828 17711 17830 17720
rect 17776 17682 17828 17688
rect 17696 17202 17724 17682
rect 18340 17338 18368 18702
rect 18432 18426 18460 19264
rect 18512 19246 18564 19252
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18510 19000 18566 19009
rect 18708 18986 18736 19246
rect 18566 18958 18736 18986
rect 18510 18935 18566 18944
rect 18524 18834 18552 18935
rect 18892 18873 18920 19994
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18878 18864 18934 18873
rect 18512 18828 18564 18834
rect 18984 18834 19012 19246
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19076 18834 19104 19110
rect 18878 18799 18934 18808
rect 18972 18828 19024 18834
rect 18512 18770 18564 18776
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18524 18306 18552 18634
rect 18432 18278 18552 18306
rect 18432 18154 18460 18278
rect 18892 18222 18920 18799
rect 18972 18770 19024 18776
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19984 18760 20036 18766
rect 18970 18728 19026 18737
rect 19984 18702 20036 18708
rect 18970 18663 18972 18672
rect 19024 18663 19026 18672
rect 18972 18634 19024 18640
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19338 18456 19394 18465
rect 19574 18448 19882 18468
rect 19338 18391 19340 18400
rect 19392 18391 19394 18400
rect 19340 18362 19392 18368
rect 19996 18358 20024 18702
rect 19984 18352 20036 18358
rect 19338 18320 19394 18329
rect 19984 18294 20036 18300
rect 19338 18255 19340 18264
rect 19392 18255 19394 18264
rect 19340 18226 19392 18232
rect 18512 18216 18564 18222
rect 18880 18216 18932 18222
rect 18512 18158 18564 18164
rect 18708 18176 18880 18204
rect 18420 18148 18472 18154
rect 18420 18090 18472 18096
rect 18524 18057 18552 18158
rect 18604 18080 18656 18086
rect 18510 18048 18566 18057
rect 18604 18022 18656 18028
rect 18510 17983 18566 17992
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 17868 17264 17920 17270
rect 17920 17212 18000 17218
rect 17868 17206 18000 17212
rect 17684 17196 17736 17202
rect 17880 17190 18000 17206
rect 17684 17138 17736 17144
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17132 16652 17184 16658
rect 17500 16652 17552 16658
rect 17132 16594 17184 16600
rect 17420 16612 17500 16640
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 17052 15570 17080 16526
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 17144 15094 17172 15370
rect 17132 15088 17184 15094
rect 17132 15030 17184 15036
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 17052 14618 17080 14894
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17144 14414 17172 15030
rect 17236 14958 17264 15506
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17144 13870 17172 14350
rect 17236 14346 17264 14894
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17236 13938 17264 14282
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 16948 13796 17000 13802
rect 16948 13738 17000 13744
rect 17144 11762 17172 13806
rect 17420 12306 17448 16612
rect 17500 16594 17552 16600
rect 17880 16114 17908 17070
rect 17972 16250 18000 17190
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18156 16658 18184 17070
rect 18144 16652 18196 16658
rect 18144 16594 18196 16600
rect 18248 16454 18276 17138
rect 18616 17134 18644 18022
rect 18708 17134 18736 18176
rect 18880 18158 18932 18164
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 19076 18057 19104 18090
rect 19720 18086 19748 18158
rect 19156 18080 19208 18086
rect 19062 18048 19118 18057
rect 19156 18022 19208 18028
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19062 17983 19118 17992
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 18892 17610 18920 17818
rect 18984 17678 19012 17818
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18788 17604 18840 17610
rect 18788 17546 18840 17552
rect 18880 17604 18932 17610
rect 18880 17546 18932 17552
rect 18800 17338 18828 17546
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18972 17196 19024 17202
rect 19076 17184 19104 17983
rect 19024 17156 19104 17184
rect 18972 17138 19024 17144
rect 19168 17134 19196 18022
rect 19984 17808 20036 17814
rect 19984 17750 20036 17756
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19996 17066 20024 17750
rect 20180 17678 20208 20420
rect 20720 20402 20772 20408
rect 20732 20058 20760 20402
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20640 19242 20668 19382
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20732 18086 20760 19858
rect 21100 19854 21128 20198
rect 21192 19854 21220 21422
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21468 19786 21496 19994
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20824 18358 20852 19382
rect 21652 19174 21680 24890
rect 22468 23180 22520 23186
rect 22468 23122 22520 23128
rect 22480 22030 22508 23122
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 21732 21956 21784 21962
rect 21732 21898 21784 21904
rect 21744 21690 21772 21898
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22204 21690 22232 21830
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22100 21616 22152 21622
rect 22100 21558 22152 21564
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 21730 19816 21786 19825
rect 21730 19751 21786 19760
rect 21824 19780 21876 19786
rect 21744 19718 21772 19751
rect 21824 19722 21876 19728
rect 21732 19712 21784 19718
rect 21732 19654 21784 19660
rect 21836 19446 21864 19722
rect 21824 19440 21876 19446
rect 21824 19382 21876 19388
rect 21928 19378 21956 20198
rect 22112 20058 22140 21558
rect 23124 20466 23152 21966
rect 23940 21412 23992 21418
rect 23940 21354 23992 21360
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23112 20460 23164 20466
rect 23296 20460 23348 20466
rect 23164 20420 23244 20448
rect 23112 20402 23164 20408
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 21008 18426 21036 18906
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20824 18193 20852 18294
rect 20810 18184 20866 18193
rect 20810 18119 20866 18128
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 20180 16658 20208 17614
rect 20548 17202 20576 17682
rect 20810 17640 20866 17649
rect 20810 17575 20866 17584
rect 20904 17604 20956 17610
rect 20824 17542 20852 17575
rect 20904 17546 20956 17552
rect 20812 17536 20864 17542
rect 20916 17513 20944 17546
rect 20812 17478 20864 17484
rect 20902 17504 20958 17513
rect 20902 17439 20958 17448
rect 20628 17264 20680 17270
rect 20628 17206 20680 17212
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 18248 16114 18276 16390
rect 18432 16114 18460 16594
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 17776 15632 17828 15638
rect 17776 15574 17828 15580
rect 17788 15502 17816 15574
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17604 15162 17632 15438
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17880 15026 17908 16050
rect 20180 15502 20208 16594
rect 20640 16454 20668 17206
rect 20810 16824 20866 16833
rect 20810 16759 20866 16768
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17512 14414 17540 14962
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17604 14482 17632 14554
rect 17788 14482 17816 14894
rect 17972 14618 18000 15030
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17866 14512 17922 14521
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17776 14476 17828 14482
rect 17866 14447 17868 14456
rect 17776 14418 17828 14424
rect 17920 14447 17922 14456
rect 17868 14418 17920 14424
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17512 13938 17540 14350
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17788 13802 17816 14418
rect 17972 13870 18000 14554
rect 19444 13938 19472 15438
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 18064 12306 18092 13738
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18156 13326 18184 13670
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18156 12918 18184 13262
rect 18524 12918 18552 13874
rect 19444 13734 19472 13874
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19996 13530 20024 13874
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16868 10674 16896 11086
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 9722 16712 10406
rect 16868 10130 16896 10610
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16592 9438 16712 9466
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16316 7274 16344 8910
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 16040 3534 16068 4014
rect 16408 3670 16436 4082
rect 16396 3664 16448 3670
rect 16396 3606 16448 3612
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 15568 3528 15620 3534
rect 15566 3496 15568 3505
rect 16028 3528 16080 3534
rect 15620 3496 15622 3505
rect 16212 3528 16264 3534
rect 16028 3470 16080 3476
rect 16132 3488 16212 3516
rect 15566 3431 15622 3440
rect 15580 2990 15608 3431
rect 16040 3398 16068 3470
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16040 3058 16068 3334
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15396 2746 15516 2774
rect 15396 2650 15424 2746
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15580 2446 15608 2926
rect 16132 2825 16160 3488
rect 16212 3470 16264 3476
rect 16118 2816 16174 2825
rect 16118 2751 16174 2760
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15764 1494 15792 2382
rect 16132 1970 16160 2751
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 16316 1816 16344 3538
rect 16500 3534 16528 4558
rect 16488 3528 16540 3534
rect 16486 3496 16488 3505
rect 16540 3496 16542 3505
rect 16486 3431 16542 3440
rect 16592 3398 16620 8774
rect 16684 8430 16712 9438
rect 16868 8906 16896 10066
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16868 8498 16896 8842
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16684 7342 16712 8366
rect 16868 7410 16896 8434
rect 16960 8362 16988 11630
rect 17052 11558 17080 11630
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 18064 11218 18092 12242
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 17144 10606 17172 11154
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 17052 8634 17080 8842
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 17040 7268 17092 7274
rect 17040 7210 17092 7216
rect 17052 6984 17080 7210
rect 17132 6996 17184 7002
rect 17052 6956 17132 6984
rect 17132 6938 17184 6944
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16868 5914 16896 6190
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16500 3126 16528 3334
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16868 2582 16896 2994
rect 16960 2854 16988 6190
rect 17144 5710 17172 6938
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17144 3058 17172 3470
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17236 2922 17264 9590
rect 17420 8974 17448 10542
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17420 7342 17448 8910
rect 17880 8634 17908 10678
rect 18064 10130 18092 11154
rect 18156 10606 18184 12854
rect 18524 12714 18552 12854
rect 19444 12850 19472 13194
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 19352 12374 19380 12718
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18984 11762 19012 12242
rect 19444 11762 19472 12786
rect 20088 12434 20116 14214
rect 20640 14074 20668 14282
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20088 12406 20300 12434
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 10742 18828 11494
rect 18788 10736 18840 10742
rect 18788 10678 18840 10684
rect 19168 10674 19196 11698
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18156 9586 18184 10542
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 18156 9382 18184 9522
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 18156 8498 18184 9318
rect 19168 9178 19196 9522
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19352 9042 19380 9522
rect 19444 9450 19472 11086
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19444 8838 19472 9386
rect 19996 8974 20024 11698
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17420 6866 17448 7278
rect 17512 6866 17540 8026
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17328 6458 17356 6734
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17420 5778 17448 6802
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17420 3369 17448 3538
rect 17500 3392 17552 3398
rect 17406 3360 17462 3369
rect 17500 3334 17552 3340
rect 17406 3295 17462 3304
rect 17512 2990 17540 3334
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 17604 2446 17632 7958
rect 18156 6322 18184 8434
rect 19260 8090 19288 8434
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19260 7478 19288 7890
rect 19996 7886 20024 8910
rect 20088 8634 20116 9998
rect 20168 9104 20220 9110
rect 20168 9046 20220 9052
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19168 6730 19196 7346
rect 19352 7206 19380 7686
rect 19444 7342 19472 7822
rect 20088 7818 20116 8570
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 20180 7274 20208 9046
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19708 6996 19760 7002
rect 19708 6938 19760 6944
rect 19432 6928 19484 6934
rect 19432 6870 19484 6876
rect 19444 6798 19472 6870
rect 19720 6798 19748 6938
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18156 3126 18184 6258
rect 19168 6118 19196 6666
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19260 6390 19288 6598
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 19352 5846 19380 6598
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 19338 5672 19394 5681
rect 19338 5607 19394 5616
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18248 4146 18276 4490
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18144 3120 18196 3126
rect 18144 3062 18196 3068
rect 18156 2990 18184 3062
rect 18144 2984 18196 2990
rect 18050 2952 18106 2961
rect 18144 2926 18196 2932
rect 18050 2887 18106 2896
rect 18064 2854 18092 2887
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16224 1788 16344 1816
rect 15752 1488 15804 1494
rect 15752 1430 15804 1436
rect 16224 800 16252 1788
rect 16776 800 16804 2246
rect 16868 1970 16896 2382
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 17236 800 17264 2246
rect 17696 800 17724 2790
rect 18340 2582 18368 5170
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18524 4622 18552 4966
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18524 4146 18552 4558
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 18708 4146 18736 4422
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18788 3936 18840 3942
rect 18786 3904 18788 3913
rect 18840 3904 18842 3913
rect 18786 3839 18842 3848
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18420 2644 18472 2650
rect 18420 2586 18472 2592
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 18432 2446 18460 2586
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18708 800 18736 3470
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 18800 2514 18828 3062
rect 19168 2774 19196 3402
rect 19260 3126 19288 4422
rect 19352 4214 19380 5607
rect 19444 5370 19472 6734
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19444 4690 19472 4966
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19996 4622 20024 7210
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 20088 5030 20116 5170
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 20088 4554 20116 4966
rect 20076 4548 20128 4554
rect 20076 4490 20128 4496
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 19444 4146 19472 4422
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19432 3936 19484 3942
rect 19524 3936 19576 3942
rect 19432 3878 19484 3884
rect 19522 3904 19524 3913
rect 19576 3904 19578 3913
rect 19248 3120 19300 3126
rect 19248 3062 19300 3068
rect 19444 2774 19472 3878
rect 19522 3839 19578 3848
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 20088 2854 20116 4490
rect 20180 4078 20208 7210
rect 20272 7206 20300 12406
rect 20350 9480 20406 9489
rect 20350 9415 20406 9424
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20272 4826 20300 5102
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20272 4622 20300 4762
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20364 4486 20392 9415
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20272 3534 20300 4014
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20076 2848 20128 2854
rect 20074 2816 20076 2825
rect 20128 2816 20130 2825
rect 19168 2746 19288 2774
rect 19444 2746 19564 2774
rect 20074 2751 20130 2760
rect 19260 2514 19288 2746
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19536 2446 19564 2746
rect 19524 2440 19576 2446
rect 19260 2378 19472 2394
rect 19524 2382 19576 2388
rect 19248 2372 19484 2378
rect 19300 2366 19432 2372
rect 19248 2314 19300 2320
rect 19432 2314 19484 2320
rect 19156 2304 19208 2310
rect 19156 2246 19208 2252
rect 19168 800 19196 2246
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19708 1420 19760 1426
rect 19708 1362 19760 1368
rect 19720 800 19748 1362
rect 20180 800 20208 3334
rect 20456 2990 20484 13398
rect 20640 13190 20668 14010
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20824 12442 20852 16759
rect 21008 13870 21036 18362
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21560 15026 21588 15302
rect 21548 15020 21600 15026
rect 21548 14962 21600 14968
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 20812 12436 20864 12442
rect 21192 12434 21220 14418
rect 21456 12708 21508 12714
rect 21456 12650 21508 12656
rect 20812 12378 20864 12384
rect 21100 12406 21220 12434
rect 21364 12436 21416 12442
rect 21100 12170 21128 12406
rect 21364 12378 21416 12384
rect 21088 12164 21140 12170
rect 21088 12106 21140 12112
rect 21100 7954 21128 12106
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 21192 10742 21220 11018
rect 21180 10736 21232 10742
rect 21284 10713 21312 11630
rect 21180 10678 21232 10684
rect 21270 10704 21326 10713
rect 21270 10639 21326 10648
rect 21180 8560 21232 8566
rect 21180 8502 21232 8508
rect 21088 7948 21140 7954
rect 21088 7890 21140 7896
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20548 7342 20576 7686
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20640 6322 20668 6734
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20548 4282 20576 4422
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20272 1426 20300 2790
rect 20260 1420 20312 1426
rect 20260 1362 20312 1368
rect 21100 800 21128 3470
rect 21192 3398 21220 8502
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 21284 7274 21312 8434
rect 21376 8294 21404 12378
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21272 7268 21324 7274
rect 21272 7210 21324 7216
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21284 4826 21312 5850
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 21376 2650 21404 6258
rect 21468 5642 21496 12650
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21560 12209 21588 12242
rect 21546 12200 21602 12209
rect 21546 12135 21602 12144
rect 21548 11688 21600 11694
rect 21548 11630 21600 11636
rect 21560 11354 21588 11630
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21652 7750 21680 19110
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21928 18193 21956 18226
rect 21914 18184 21970 18193
rect 21914 18119 21970 18128
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21836 17678 21864 18022
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 21836 16250 21864 16458
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21836 15162 21864 15370
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21744 12170 21772 13126
rect 21928 12850 21956 13262
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21928 12442 21956 12786
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21732 12164 21784 12170
rect 21732 12106 21784 12112
rect 21836 12073 21864 12174
rect 21822 12064 21878 12073
rect 21822 11999 21878 12008
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21744 10674 21772 10950
rect 21732 10668 21784 10674
rect 21732 10610 21784 10616
rect 21744 10470 21772 10610
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21744 9994 21772 10406
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 21744 9110 21772 9930
rect 21836 9654 21864 11494
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 21824 9648 21876 9654
rect 21824 9590 21876 9596
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21928 8906 21956 9998
rect 22020 9738 22048 19994
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 22112 19378 22140 19722
rect 22204 19514 22232 19858
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22112 13818 22140 19314
rect 22192 18352 22244 18358
rect 22190 18320 22192 18329
rect 22244 18320 22246 18329
rect 22190 18255 22246 18264
rect 22376 18284 22428 18290
rect 22204 17814 22232 18255
rect 22376 18226 22428 18232
rect 22192 17808 22244 17814
rect 22192 17750 22244 17756
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22204 16250 22232 16390
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22388 16114 22416 18226
rect 23216 18222 23244 20420
rect 23296 20402 23348 20408
rect 23308 20058 23336 20402
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23664 19916 23716 19922
rect 23664 19858 23716 19864
rect 23676 18850 23704 19858
rect 23768 19854 23796 20470
rect 23756 19848 23808 19854
rect 23848 19848 23900 19854
rect 23756 19790 23808 19796
rect 23846 19816 23848 19825
rect 23900 19816 23902 19825
rect 23846 19751 23902 19760
rect 23860 19514 23888 19751
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 23676 18822 23796 18850
rect 23664 18692 23716 18698
rect 23664 18634 23716 18640
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 23216 17270 23244 18158
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22204 13938 22232 16050
rect 22468 14000 22520 14006
rect 22468 13942 22520 13948
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22112 13790 22232 13818
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 22112 13258 22140 13466
rect 22100 13252 22152 13258
rect 22100 13194 22152 13200
rect 22204 13190 22232 13790
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22204 11830 22232 12718
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 22296 11762 22324 12378
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22112 10810 22140 11698
rect 22284 11144 22336 11150
rect 22204 11092 22284 11098
rect 22204 11086 22336 11092
rect 22204 11070 22324 11086
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22204 10742 22232 11070
rect 22192 10736 22244 10742
rect 22192 10678 22244 10684
rect 22284 10736 22336 10742
rect 22284 10678 22336 10684
rect 22020 9710 22140 9738
rect 22112 8945 22140 9710
rect 22098 8936 22154 8945
rect 21916 8900 21968 8906
rect 22098 8871 22154 8880
rect 21916 8842 21968 8848
rect 21732 8492 21784 8498
rect 21928 8480 21956 8842
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22112 8498 22140 8774
rect 21784 8452 21956 8480
rect 22100 8492 22152 8498
rect 21732 8434 21784 8440
rect 22100 8434 22152 8440
rect 21824 8356 21876 8362
rect 21824 8298 21876 8304
rect 21730 8256 21786 8265
rect 21730 8191 21786 8200
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21744 6934 21772 8191
rect 21732 6928 21784 6934
rect 21732 6870 21784 6876
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 21836 5166 21864 8298
rect 22100 6384 22152 6390
rect 22100 6326 22152 6332
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 21640 5092 21692 5098
rect 21640 5034 21692 5040
rect 21652 4690 21680 5034
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21836 4622 21864 5102
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 22020 4146 22048 5714
rect 22112 5710 22140 6326
rect 22204 5846 22232 10678
rect 22296 9722 22324 10678
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22296 6322 22324 9658
rect 22388 7410 22416 12174
rect 22480 10198 22508 13942
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22664 12782 22692 13330
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22756 12434 22784 16730
rect 23032 16658 23060 17138
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23020 16108 23072 16114
rect 23020 16050 23072 16056
rect 23032 15570 23060 16050
rect 23020 15564 23072 15570
rect 23020 15506 23072 15512
rect 23032 15094 23060 15506
rect 23020 15088 23072 15094
rect 23020 15030 23072 15036
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22848 14414 22876 14962
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22848 13530 22876 14350
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 22836 13524 22888 13530
rect 22836 13466 22888 13472
rect 23032 13410 23060 13806
rect 23124 13530 23152 16526
rect 23216 16114 23244 17206
rect 23480 16516 23532 16522
rect 23480 16458 23532 16464
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 23400 15026 23428 15370
rect 23492 15162 23520 16458
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23400 14770 23428 14962
rect 23216 14742 23428 14770
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23032 13382 23152 13410
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22848 12782 22876 13262
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22664 12406 22784 12434
rect 22560 11212 22612 11218
rect 22560 11154 22612 11160
rect 22572 10674 22600 11154
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22468 10192 22520 10198
rect 22468 10134 22520 10140
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22480 9382 22508 9998
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22480 8498 22508 9318
rect 22560 9172 22612 9178
rect 22560 9114 22612 9120
rect 22572 8974 22600 9114
rect 22664 8974 22692 12406
rect 22848 12238 22876 12718
rect 23124 12646 23152 13382
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 23112 12640 23164 12646
rect 23112 12582 23164 12588
rect 22836 12232 22888 12238
rect 22742 12200 22798 12209
rect 22940 12209 22968 12582
rect 23124 12442 23152 12582
rect 23112 12436 23164 12442
rect 23112 12378 23164 12384
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 22836 12174 22888 12180
rect 22926 12200 22982 12209
rect 22742 12135 22798 12144
rect 22926 12135 22982 12144
rect 22756 12102 22784 12135
rect 22744 12096 22796 12102
rect 22940 12084 22968 12135
rect 22940 12056 23060 12084
rect 22744 12038 22796 12044
rect 22928 11280 22980 11286
rect 22926 11248 22928 11257
rect 22980 11248 22982 11257
rect 22926 11183 22982 11192
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22468 8356 22520 8362
rect 22468 8298 22520 8304
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22480 7206 22508 8298
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22572 6390 22600 8910
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22572 6236 22600 6326
rect 22480 6208 22600 6236
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 22192 5840 22244 5846
rect 22192 5782 22244 5788
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 22112 5370 22140 5646
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22204 4826 22232 5170
rect 22192 4820 22244 4826
rect 22192 4762 22244 4768
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21560 3602 21588 3878
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21928 3641 21956 3674
rect 21914 3632 21970 3641
rect 21548 3596 21600 3602
rect 21914 3567 21970 3576
rect 21548 3538 21600 3544
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21652 2836 21680 3130
rect 21836 2990 21864 3402
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22204 3074 22232 3334
rect 22020 3046 22232 3074
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 22020 2836 22048 3046
rect 21652 2808 22048 2836
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 22296 2446 22324 6054
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 21652 800 21680 2246
rect 22112 800 22140 2246
rect 22480 1970 22508 6208
rect 22664 5681 22692 8910
rect 22756 8838 22784 9862
rect 23032 9110 23060 12056
rect 23124 11286 23152 12242
rect 23112 11280 23164 11286
rect 23112 11222 23164 11228
rect 23124 10810 23152 11222
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 23112 9716 23164 9722
rect 23112 9658 23164 9664
rect 23020 9104 23072 9110
rect 23020 9046 23072 9052
rect 23124 8888 23152 9658
rect 23216 9654 23244 14742
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23296 13456 23348 13462
rect 23296 13398 23348 13404
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 23204 9376 23256 9382
rect 23204 9318 23256 9324
rect 23216 9178 23244 9318
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 23204 8900 23256 8906
rect 23124 8860 23204 8888
rect 23204 8842 23256 8848
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22756 6798 22784 7142
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22848 6662 22876 7482
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22650 5672 22706 5681
rect 22650 5607 22706 5616
rect 23124 4486 23152 8026
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23216 6934 23244 7346
rect 23204 6928 23256 6934
rect 23204 6870 23256 6876
rect 23308 5710 23336 13398
rect 23400 9926 23428 14554
rect 23492 14006 23520 15098
rect 23676 14074 23704 18634
rect 23768 15706 23796 18822
rect 23756 15700 23808 15706
rect 23756 15642 23808 15648
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23480 14000 23532 14006
rect 23480 13942 23532 13948
rect 23492 13258 23520 13942
rect 23676 13734 23704 14010
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23768 13682 23796 15642
rect 23952 15162 23980 21354
rect 24504 21350 24532 26794
rect 24584 24404 24636 24410
rect 24584 24346 24636 24352
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24492 20324 24544 20330
rect 24492 20266 24544 20272
rect 24504 19922 24532 20266
rect 24492 19916 24544 19922
rect 24492 19858 24544 19864
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24228 19378 24256 19654
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24216 19236 24268 19242
rect 24216 19178 24268 19184
rect 24228 18222 24256 19178
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 24412 17814 24440 18226
rect 24596 18170 24624 24346
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 24688 22778 24716 22986
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 25056 22778 25084 22918
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 25044 22772 25096 22778
rect 25044 22714 25096 22720
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 25056 22030 25084 22578
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 24688 21554 24716 21966
rect 25136 21956 25188 21962
rect 25136 21898 25188 21904
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 24952 21616 25004 21622
rect 24952 21558 25004 21564
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24688 20058 24716 21490
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 24504 18142 24624 18170
rect 24400 17808 24452 17814
rect 24400 17750 24452 17756
rect 24398 16960 24454 16969
rect 24398 16895 24454 16904
rect 24412 16794 24440 16895
rect 24504 16794 24532 18142
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24596 17542 24624 18022
rect 24964 17762 24992 21558
rect 25056 21486 25084 21830
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 25056 20754 25084 21422
rect 25148 21350 25176 21898
rect 25332 21350 25360 31078
rect 25504 28008 25556 28014
rect 25504 27950 25556 27956
rect 25516 22234 25544 27950
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 33508 23112 33560 23118
rect 33508 23054 33560 23060
rect 25688 22704 25740 22710
rect 25688 22646 25740 22652
rect 25700 22234 25728 22646
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25792 22234 25820 22510
rect 27632 22438 27660 23054
rect 27988 23044 28040 23050
rect 27988 22986 28040 22992
rect 28000 22778 28028 22986
rect 29552 22976 29604 22982
rect 29552 22918 29604 22924
rect 27988 22772 28040 22778
rect 27988 22714 28040 22720
rect 28172 22772 28224 22778
rect 28172 22714 28224 22720
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 25504 22228 25556 22234
rect 25504 22170 25556 22176
rect 25688 22228 25740 22234
rect 25688 22170 25740 22176
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 25412 21888 25464 21894
rect 25412 21830 25464 21836
rect 25424 21622 25452 21830
rect 25412 21616 25464 21622
rect 25412 21558 25464 21564
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 25148 20942 25176 21286
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 25056 20726 25176 20754
rect 25148 20534 25176 20726
rect 25136 20528 25188 20534
rect 25136 20470 25188 20476
rect 24964 17734 25084 17762
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24492 16788 24544 16794
rect 24492 16730 24544 16736
rect 24780 16590 24808 17614
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24676 16516 24728 16522
rect 24676 16458 24728 16464
rect 24688 16402 24716 16458
rect 24688 16374 24900 16402
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24412 15706 24440 16050
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24504 15502 24532 15642
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24688 15162 24716 15438
rect 24780 15366 24808 15846
rect 24872 15366 24900 16374
rect 24964 15502 24992 17614
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24860 15360 24912 15366
rect 24860 15302 24912 15308
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 23848 14952 23900 14958
rect 23848 14894 23900 14900
rect 23860 13870 23888 14894
rect 23952 14822 23980 15098
rect 24308 15088 24360 15094
rect 24308 15030 24360 15036
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 23480 13252 23532 13258
rect 23480 13194 23532 13200
rect 23492 12170 23520 13194
rect 23676 12434 23704 13670
rect 23768 13654 23888 13682
rect 23676 12406 23796 12434
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23584 11354 23612 11698
rect 23572 11348 23624 11354
rect 23572 11290 23624 11296
rect 23664 9988 23716 9994
rect 23664 9930 23716 9936
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23400 9382 23428 9590
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23400 7002 23428 7414
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 23400 6458 23428 6938
rect 23388 6452 23440 6458
rect 23388 6394 23440 6400
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23112 4480 23164 4486
rect 23112 4422 23164 4428
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22572 2446 22600 3538
rect 22664 3126 22692 3878
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22652 3120 22704 3126
rect 22652 3062 22704 3068
rect 22848 2990 22876 3334
rect 22836 2984 22888 2990
rect 22836 2926 22888 2932
rect 23216 2854 23244 4558
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23492 3534 23520 3878
rect 23676 3670 23704 9930
rect 23768 7002 23796 12406
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 23860 6186 23888 13654
rect 24044 13190 24072 14962
rect 24320 14482 24348 15030
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24308 14476 24360 14482
rect 24308 14418 24360 14424
rect 24400 14340 24452 14346
rect 24400 14282 24452 14288
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 24044 12442 24072 12922
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 24136 11830 24164 13806
rect 24308 13728 24360 13734
rect 24308 13670 24360 13676
rect 24124 11824 24176 11830
rect 24124 11766 24176 11772
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24228 11558 24256 11630
rect 24216 11552 24268 11558
rect 24216 11494 24268 11500
rect 24320 8022 24348 13670
rect 24412 8566 24440 14282
rect 24504 13546 24532 14758
rect 24584 14544 24636 14550
rect 24584 14486 24636 14492
rect 24596 13734 24624 14486
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24504 13518 24624 13546
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24504 11830 24532 12922
rect 24492 11824 24544 11830
rect 24492 11766 24544 11772
rect 24504 11286 24532 11766
rect 24492 11280 24544 11286
rect 24492 11222 24544 11228
rect 24596 10146 24624 13518
rect 24688 12986 24716 13874
rect 24780 13326 24808 14010
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24780 12986 24808 13262
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24688 12050 24716 12378
rect 24780 12186 24808 12922
rect 24872 12646 24900 15302
rect 24952 14884 25004 14890
rect 24952 14826 25004 14832
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24964 12434 24992 14826
rect 25056 13394 25084 17734
rect 25148 13954 25176 20470
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25332 14074 25360 18226
rect 25412 17604 25464 17610
rect 25412 17546 25464 17552
rect 25424 17270 25452 17546
rect 25412 17264 25464 17270
rect 25412 17206 25464 17212
rect 25424 15570 25452 17206
rect 25412 15564 25464 15570
rect 25412 15506 25464 15512
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25148 13926 25360 13954
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24964 12406 25084 12434
rect 24780 12170 24900 12186
rect 24780 12164 24912 12170
rect 24780 12158 24860 12164
rect 24860 12106 24912 12112
rect 24688 12022 24808 12050
rect 24504 10118 24624 10146
rect 24400 8560 24452 8566
rect 24400 8502 24452 8508
rect 24504 8378 24532 10118
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24596 8974 24624 9998
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24688 9042 24716 9454
rect 24780 9110 24808 12022
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24872 10810 24900 11018
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24964 10674 24992 11494
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 24952 10532 25004 10538
rect 24952 10474 25004 10480
rect 24964 10062 24992 10474
rect 25056 10146 25084 12406
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25240 11082 25268 12038
rect 25228 11076 25280 11082
rect 25228 11018 25280 11024
rect 25056 10118 25176 10146
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24676 9036 24728 9042
rect 24676 8978 24728 8984
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24596 8498 24624 8910
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24504 8350 24624 8378
rect 24308 8016 24360 8022
rect 24308 7958 24360 7964
rect 24398 7984 24454 7993
rect 24398 7919 24454 7928
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24136 7478 24164 7686
rect 24124 7472 24176 7478
rect 24124 7414 24176 7420
rect 24412 7274 24440 7919
rect 24490 7848 24546 7857
rect 24490 7783 24492 7792
rect 24544 7783 24546 7792
rect 24492 7754 24544 7760
rect 24400 7268 24452 7274
rect 24400 7210 24452 7216
rect 24492 7200 24544 7206
rect 24492 7142 24544 7148
rect 23848 6180 23900 6186
rect 23848 6122 23900 6128
rect 24504 4826 24532 7142
rect 24596 6458 24624 8350
rect 24676 8084 24728 8090
rect 24676 8026 24728 8032
rect 24688 7206 24716 8026
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 24492 4820 24544 4826
rect 24492 4762 24544 4768
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 23664 3664 23716 3670
rect 23664 3606 23716 3612
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 22468 1964 22520 1970
rect 22468 1906 22520 1912
rect 22572 870 22692 898
rect 22572 800 22600 870
rect 9048 734 9260 762
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15750 0 15806 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 22664 762 22692 870
rect 22848 762 22876 2246
rect 23216 1494 23244 2790
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23308 1494 23336 2382
rect 23204 1488 23256 1494
rect 23204 1430 23256 1436
rect 23296 1488 23348 1494
rect 23296 1430 23348 1436
rect 23584 800 23612 3470
rect 23664 3460 23716 3466
rect 23664 3402 23716 3408
rect 23676 3058 23704 3402
rect 24412 3126 24440 4422
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 24780 2446 24808 8434
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 24872 7546 24900 7686
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 24964 6118 24992 9998
rect 25056 8974 25084 9998
rect 25148 9178 25176 10118
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 25240 9518 25268 9998
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 25240 8974 25268 9454
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 25056 8634 25084 8910
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 25240 8498 25268 8910
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25332 8378 25360 13926
rect 25412 13388 25464 13394
rect 25412 13330 25464 13336
rect 25424 12782 25452 13330
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25056 8350 25360 8378
rect 25056 7857 25084 8350
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 25042 7848 25098 7857
rect 25042 7783 25098 7792
rect 25148 7546 25176 7890
rect 25228 7880 25280 7886
rect 25424 7834 25452 12718
rect 25280 7828 25452 7834
rect 25228 7822 25452 7828
rect 25240 7806 25452 7822
rect 25412 7744 25464 7750
rect 25412 7686 25464 7692
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 25240 7410 25268 7482
rect 25424 7478 25452 7686
rect 25516 7478 25544 22170
rect 26160 21690 26188 22170
rect 26148 21684 26200 21690
rect 26148 21626 26200 21632
rect 26056 21616 26108 21622
rect 26056 21558 26108 21564
rect 25596 21412 25648 21418
rect 25596 21354 25648 21360
rect 25608 16674 25636 21354
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25700 20466 25728 20742
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25780 16992 25832 16998
rect 25780 16934 25832 16940
rect 25686 16824 25742 16833
rect 25792 16794 25820 16934
rect 25884 16810 25912 21286
rect 26068 20534 26096 21558
rect 27632 21486 27660 22374
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 26056 20528 26108 20534
rect 26056 20470 26108 20476
rect 25964 17604 26016 17610
rect 25964 17546 26016 17552
rect 25976 16998 26004 17546
rect 26068 17082 26096 20470
rect 27632 19854 27660 21422
rect 27908 21146 27936 21490
rect 27896 21140 27948 21146
rect 27896 21082 27948 21088
rect 28184 20942 28212 22714
rect 28264 22500 28316 22506
rect 28264 22442 28316 22448
rect 28172 20936 28224 20942
rect 28172 20878 28224 20884
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 26976 19780 27028 19786
rect 26976 19722 27028 19728
rect 26988 19514 27016 19722
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 27080 19514 27108 19654
rect 26976 19508 27028 19514
rect 26976 19450 27028 19456
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 27988 19372 28040 19378
rect 27988 19314 28040 19320
rect 27160 19304 27212 19310
rect 27160 19246 27212 19252
rect 26884 19168 26936 19174
rect 26884 19110 26936 19116
rect 26896 18834 26924 19110
rect 27172 18970 27200 19246
rect 27160 18964 27212 18970
rect 27160 18906 27212 18912
rect 27712 18896 27764 18902
rect 27712 18838 27764 18844
rect 27804 18896 27856 18902
rect 27804 18838 27856 18844
rect 26884 18828 26936 18834
rect 26884 18770 26936 18776
rect 27252 18760 27304 18766
rect 27252 18702 27304 18708
rect 27160 18692 27212 18698
rect 27160 18634 27212 18640
rect 27172 18290 27200 18634
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 26422 18184 26478 18193
rect 26422 18119 26478 18128
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26160 17202 26188 17478
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26068 17054 26188 17082
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25686 16759 25688 16768
rect 25740 16759 25742 16768
rect 25780 16788 25832 16794
rect 25688 16730 25740 16736
rect 25884 16782 26004 16810
rect 25780 16730 25832 16736
rect 25608 16646 25912 16674
rect 25688 16516 25740 16522
rect 25688 16458 25740 16464
rect 25700 16182 25728 16458
rect 25780 16448 25832 16454
rect 25778 16416 25780 16425
rect 25832 16416 25834 16425
rect 25778 16351 25834 16360
rect 25688 16176 25740 16182
rect 25688 16118 25740 16124
rect 25780 15904 25832 15910
rect 25780 15846 25832 15852
rect 25688 14408 25740 14414
rect 25688 14350 25740 14356
rect 25700 13938 25728 14350
rect 25688 13932 25740 13938
rect 25688 13874 25740 13880
rect 25688 13796 25740 13802
rect 25688 13738 25740 13744
rect 25596 13728 25648 13734
rect 25596 13670 25648 13676
rect 25608 12442 25636 13670
rect 25700 13326 25728 13738
rect 25688 13320 25740 13326
rect 25688 13262 25740 13268
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25596 12164 25648 12170
rect 25596 12106 25648 12112
rect 25608 10538 25636 12106
rect 25596 10532 25648 10538
rect 25596 10474 25648 10480
rect 25700 9518 25728 12582
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 25594 7984 25650 7993
rect 25594 7919 25596 7928
rect 25648 7919 25650 7928
rect 25596 7890 25648 7896
rect 25700 7834 25728 9454
rect 25608 7806 25728 7834
rect 25412 7472 25464 7478
rect 25412 7414 25464 7420
rect 25504 7472 25556 7478
rect 25504 7414 25556 7420
rect 25608 7410 25636 7806
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25412 7200 25464 7206
rect 25332 7160 25412 7188
rect 25228 6860 25280 6866
rect 25228 6802 25280 6808
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 25056 4826 25084 5510
rect 25240 5234 25268 6802
rect 25332 5642 25360 7160
rect 25412 7142 25464 7148
rect 25608 6730 25636 7346
rect 25596 6724 25648 6730
rect 25596 6666 25648 6672
rect 25700 6322 25728 7686
rect 25688 6316 25740 6322
rect 25688 6258 25740 6264
rect 25792 6118 25820 15846
rect 25780 6112 25832 6118
rect 25780 6054 25832 6060
rect 25884 5778 25912 16646
rect 25976 15910 26004 16782
rect 25964 15904 26016 15910
rect 25964 15846 26016 15852
rect 25964 15428 26016 15434
rect 25964 15370 26016 15376
rect 25976 8634 26004 15370
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 26068 14618 26096 14894
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 26054 11248 26110 11257
rect 26054 11183 26056 11192
rect 26108 11183 26110 11192
rect 26056 11154 26108 11160
rect 26160 9382 26188 17054
rect 26330 16416 26386 16425
rect 26330 16351 26386 16360
rect 26240 15428 26292 15434
rect 26240 15370 26292 15376
rect 26252 15162 26280 15370
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26252 13258 26280 13670
rect 26240 13252 26292 13258
rect 26240 13194 26292 13200
rect 26344 10130 26372 16351
rect 26436 15094 26464 18119
rect 27160 17808 27212 17814
rect 27160 17750 27212 17756
rect 27172 17649 27200 17750
rect 27158 17640 27214 17649
rect 26516 17604 26568 17610
rect 27158 17575 27214 17584
rect 26516 17546 26568 17552
rect 26528 17513 26556 17546
rect 26514 17504 26570 17513
rect 26514 17439 26570 17448
rect 27264 16998 27292 18702
rect 27724 18086 27752 18838
rect 27816 18358 27844 18838
rect 28000 18698 28028 19314
rect 27988 18692 28040 18698
rect 27988 18634 28040 18640
rect 27804 18352 27856 18358
rect 27804 18294 27856 18300
rect 28172 18148 28224 18154
rect 28172 18090 28224 18096
rect 27528 18080 27580 18086
rect 27528 18022 27580 18028
rect 27712 18080 27764 18086
rect 27712 18022 27764 18028
rect 27540 17678 27568 18022
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 27252 16992 27304 16998
rect 27252 16934 27304 16940
rect 27528 16720 27580 16726
rect 27528 16662 27580 16668
rect 27540 15910 27568 16662
rect 28080 16584 28132 16590
rect 28080 16526 28132 16532
rect 28092 16130 28120 16526
rect 28184 16250 28212 18090
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 28092 16102 28212 16130
rect 28184 16046 28212 16102
rect 28172 16040 28224 16046
rect 28172 15982 28224 15988
rect 27528 15904 27580 15910
rect 27528 15846 27580 15852
rect 27160 15360 27212 15366
rect 27160 15302 27212 15308
rect 26424 15088 26476 15094
rect 26424 15030 26476 15036
rect 27172 15026 27200 15302
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26884 14952 26936 14958
rect 26884 14894 26936 14900
rect 26436 14074 26464 14894
rect 26896 14414 26924 14894
rect 26884 14408 26936 14414
rect 26884 14350 26936 14356
rect 27172 14346 27200 14962
rect 28184 14414 28212 15982
rect 28172 14408 28224 14414
rect 28172 14350 28224 14356
rect 27160 14340 27212 14346
rect 27160 14282 27212 14288
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26436 11762 26464 14010
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 26608 13184 26660 13190
rect 26608 13126 26660 13132
rect 26620 12170 26648 13126
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 26608 12164 26660 12170
rect 26608 12106 26660 12112
rect 26974 12064 27030 12073
rect 26974 11999 27030 12008
rect 26988 11898 27016 11999
rect 26884 11892 26936 11898
rect 26884 11834 26936 11840
rect 26976 11892 27028 11898
rect 26976 11834 27028 11840
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26516 11756 26568 11762
rect 26516 11698 26568 11704
rect 26332 10124 26384 10130
rect 26332 10066 26384 10072
rect 26148 9376 26200 9382
rect 26148 9318 26200 9324
rect 26056 8900 26108 8906
rect 26056 8842 26108 8848
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 25872 5772 25924 5778
rect 25872 5714 25924 5720
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25320 5636 25372 5642
rect 25320 5578 25372 5584
rect 25700 5370 25728 5646
rect 25688 5364 25740 5370
rect 25688 5306 25740 5312
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 25504 5228 25556 5234
rect 25504 5170 25556 5176
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25516 4622 25544 5170
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 25504 4616 25556 4622
rect 25504 4558 25556 4564
rect 24872 4282 24900 4558
rect 24952 4480 25004 4486
rect 24952 4422 25004 4428
rect 24860 4276 24912 4282
rect 24860 4218 24912 4224
rect 24964 3534 24992 4422
rect 25410 3632 25466 3641
rect 25410 3567 25466 3576
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 25424 3466 25452 3567
rect 25412 3460 25464 3466
rect 25412 3402 25464 3408
rect 25596 2916 25648 2922
rect 25700 2904 25728 5306
rect 25964 3052 26016 3058
rect 25964 2994 26016 3000
rect 25648 2876 25728 2904
rect 25596 2858 25648 2864
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24872 2446 24900 2790
rect 25044 2576 25096 2582
rect 25044 2518 25096 2524
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24032 2304 24084 2310
rect 24676 2304 24728 2310
rect 24032 2246 24084 2252
rect 24596 2264 24676 2292
rect 24044 800 24072 2246
rect 24596 800 24624 2264
rect 24676 2246 24728 2252
rect 25056 800 25084 2518
rect 25700 2446 25728 2876
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 25976 800 26004 2994
rect 26068 2922 26096 8842
rect 26160 8362 26188 9318
rect 26528 8786 26556 11698
rect 26896 11286 26924 11834
rect 26884 11280 26936 11286
rect 26884 11222 26936 11228
rect 27448 11150 27476 12378
rect 27436 11144 27488 11150
rect 27436 11086 27488 11092
rect 27448 10130 27476 11086
rect 27908 10713 27936 13262
rect 28184 13240 28212 14350
rect 28276 13308 28304 22442
rect 29564 21554 29592 22918
rect 29644 22636 29696 22642
rect 29644 22578 29696 22584
rect 29656 22098 29684 22578
rect 29748 22234 29776 23054
rect 33048 22976 33100 22982
rect 33048 22918 33100 22924
rect 33416 22976 33468 22982
rect 33416 22918 33468 22924
rect 33060 22710 33088 22918
rect 33428 22778 33456 22918
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33048 22704 33100 22710
rect 33048 22646 33100 22652
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 30852 22234 30880 22578
rect 32036 22432 32088 22438
rect 32036 22374 32088 22380
rect 29736 22228 29788 22234
rect 29736 22170 29788 22176
rect 30840 22228 30892 22234
rect 30840 22170 30892 22176
rect 29644 22092 29696 22098
rect 32048 22094 32076 22374
rect 29644 22034 29696 22040
rect 31956 22066 32076 22094
rect 32496 22092 32548 22098
rect 29736 22024 29788 22030
rect 29736 21966 29788 21972
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31300 22024 31352 22030
rect 31300 21966 31352 21972
rect 29748 21690 29776 21966
rect 30104 21956 30156 21962
rect 30104 21898 30156 21904
rect 29736 21684 29788 21690
rect 29736 21626 29788 21632
rect 29460 21548 29512 21554
rect 29460 21490 29512 21496
rect 29552 21548 29604 21554
rect 29552 21490 29604 21496
rect 29184 21344 29236 21350
rect 29184 21286 29236 21292
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 29092 20936 29144 20942
rect 29092 20878 29144 20884
rect 28448 20528 28500 20534
rect 28448 20470 28500 20476
rect 28460 19922 28488 20470
rect 28552 20058 28580 20878
rect 28908 20528 28960 20534
rect 28736 20476 28908 20482
rect 28736 20470 28960 20476
rect 28736 20454 28948 20470
rect 28632 20256 28684 20262
rect 28632 20198 28684 20204
rect 28540 20052 28592 20058
rect 28540 19994 28592 20000
rect 28448 19916 28500 19922
rect 28448 19858 28500 19864
rect 28540 19712 28592 19718
rect 28540 19654 28592 19660
rect 28552 19378 28580 19654
rect 28540 19372 28592 19378
rect 28540 19314 28592 19320
rect 28448 17536 28500 17542
rect 28448 17478 28500 17484
rect 28460 17134 28488 17478
rect 28448 17128 28500 17134
rect 28448 17070 28500 17076
rect 28460 16726 28488 17070
rect 28448 16720 28500 16726
rect 28448 16662 28500 16668
rect 28460 16182 28488 16662
rect 28540 16516 28592 16522
rect 28540 16458 28592 16464
rect 28448 16176 28500 16182
rect 28448 16118 28500 16124
rect 28552 16114 28580 16458
rect 28540 16108 28592 16114
rect 28540 16050 28592 16056
rect 28540 14816 28592 14822
rect 28540 14758 28592 14764
rect 28448 13320 28500 13326
rect 28276 13280 28448 13308
rect 28448 13262 28500 13268
rect 28184 13212 28396 13240
rect 27894 10704 27950 10713
rect 27894 10639 27896 10648
rect 27948 10639 27950 10648
rect 27896 10610 27948 10616
rect 27620 10600 27672 10606
rect 27620 10542 27672 10548
rect 27436 10124 27488 10130
rect 27436 10066 27488 10072
rect 26882 8936 26938 8945
rect 26882 8871 26938 8880
rect 26436 8758 26556 8786
rect 26148 8356 26200 8362
rect 26148 8298 26200 8304
rect 26436 8242 26464 8758
rect 26160 8214 26464 8242
rect 26160 6866 26188 8214
rect 26330 7848 26386 7857
rect 26240 7812 26292 7818
rect 26330 7783 26386 7792
rect 26240 7754 26292 7760
rect 26252 7546 26280 7754
rect 26344 7750 26372 7783
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26252 7274 26280 7482
rect 26516 7472 26568 7478
rect 26516 7414 26568 7420
rect 26240 7268 26292 7274
rect 26240 7210 26292 7216
rect 26148 6860 26200 6866
rect 26148 6802 26200 6808
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 26344 5846 26372 6802
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 26332 5840 26384 5846
rect 26332 5782 26384 5788
rect 26344 5710 26372 5782
rect 26332 5704 26384 5710
rect 26436 5688 26464 6598
rect 26332 5646 26384 5652
rect 26424 5682 26476 5688
rect 26528 5642 26556 7414
rect 26896 5778 26924 8871
rect 27632 8378 27660 10542
rect 27988 10464 28040 10470
rect 27988 10406 28040 10412
rect 28000 9586 28028 10406
rect 28080 9988 28132 9994
rect 28080 9930 28132 9936
rect 28092 9722 28120 9930
rect 28172 9920 28224 9926
rect 28172 9862 28224 9868
rect 28080 9716 28132 9722
rect 28080 9658 28132 9664
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 27804 8968 27856 8974
rect 27804 8910 27856 8916
rect 27712 8900 27764 8906
rect 27712 8842 27764 8848
rect 27724 8566 27752 8842
rect 27712 8560 27764 8566
rect 27712 8502 27764 8508
rect 27540 8350 27660 8378
rect 27436 7812 27488 7818
rect 27540 7800 27568 8350
rect 27620 8288 27672 8294
rect 27620 8230 27672 8236
rect 27632 8090 27660 8230
rect 27620 8084 27672 8090
rect 27620 8026 27672 8032
rect 27724 7818 27752 8502
rect 27816 7993 27844 8910
rect 27896 8832 27948 8838
rect 27896 8774 27948 8780
rect 27908 8294 27936 8774
rect 27896 8288 27948 8294
rect 27896 8230 27948 8236
rect 27908 8090 27936 8230
rect 27896 8084 27948 8090
rect 27896 8026 27948 8032
rect 27802 7984 27858 7993
rect 27802 7919 27858 7928
rect 27908 7886 27936 8026
rect 28184 7970 28212 9862
rect 28092 7942 28212 7970
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 27488 7772 27568 7800
rect 27712 7812 27764 7818
rect 27436 7754 27488 7760
rect 27712 7754 27764 7760
rect 27712 7336 27764 7342
rect 27710 7304 27712 7313
rect 27804 7336 27856 7342
rect 27764 7304 27766 7313
rect 27804 7278 27856 7284
rect 27710 7239 27766 7248
rect 27816 7206 27844 7278
rect 27908 7206 27936 7822
rect 27988 7744 28040 7750
rect 27988 7686 28040 7692
rect 28000 7478 28028 7686
rect 27988 7472 28040 7478
rect 27988 7414 28040 7420
rect 27804 7200 27856 7206
rect 27804 7142 27856 7148
rect 27896 7200 27948 7206
rect 27896 7142 27948 7148
rect 27802 7032 27858 7041
rect 27908 7002 27936 7142
rect 27802 6967 27804 6976
rect 27856 6967 27858 6976
rect 27896 6996 27948 7002
rect 27804 6938 27856 6944
rect 27896 6938 27948 6944
rect 28000 6662 28028 7414
rect 27528 6656 27580 6662
rect 27528 6598 27580 6604
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 27436 5908 27488 5914
rect 27436 5850 27488 5856
rect 26976 5840 27028 5846
rect 26976 5782 27028 5788
rect 26792 5772 26844 5778
rect 26792 5714 26844 5720
rect 26884 5772 26936 5778
rect 26884 5714 26936 5720
rect 26424 5624 26476 5630
rect 26516 5636 26568 5642
rect 26516 5578 26568 5584
rect 26148 5568 26200 5574
rect 26148 5510 26200 5516
rect 26160 5234 26188 5510
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 26332 5024 26384 5030
rect 26332 4966 26384 4972
rect 26240 4548 26292 4554
rect 26240 4490 26292 4496
rect 26252 3670 26280 4490
rect 26240 3664 26292 3670
rect 26240 3606 26292 3612
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 26160 2990 26188 3470
rect 26148 2984 26200 2990
rect 26148 2926 26200 2932
rect 26056 2916 26108 2922
rect 26056 2858 26108 2864
rect 26252 2446 26280 3606
rect 26344 3534 26372 4966
rect 26804 4622 26832 5714
rect 26988 5642 27016 5782
rect 27448 5710 27476 5850
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 27540 5642 27568 6598
rect 28000 5914 28028 6598
rect 27988 5908 28040 5914
rect 27988 5850 28040 5856
rect 27896 5704 27948 5710
rect 27896 5646 27948 5652
rect 26976 5636 27028 5642
rect 26976 5578 27028 5584
rect 27528 5636 27580 5642
rect 27528 5578 27580 5584
rect 27528 5160 27580 5166
rect 27528 5102 27580 5108
rect 27540 4826 27568 5102
rect 27620 5024 27672 5030
rect 27620 4966 27672 4972
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 27252 4004 27304 4010
rect 27252 3946 27304 3952
rect 27264 3738 27292 3946
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 27436 3528 27488 3534
rect 27436 3470 27488 3476
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 26528 800 26556 2246
rect 27448 800 27476 3470
rect 27632 3126 27660 4966
rect 27908 4570 27936 5646
rect 27988 5568 28040 5574
rect 27988 5510 28040 5516
rect 28000 5234 28028 5510
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 27908 4554 28028 4570
rect 27908 4548 28040 4554
rect 27908 4542 27988 4548
rect 27988 4490 28040 4496
rect 28000 3398 28028 4490
rect 28092 3398 28120 7942
rect 28172 7880 28224 7886
rect 28172 7822 28224 7828
rect 28184 7546 28212 7822
rect 28264 7744 28316 7750
rect 28264 7686 28316 7692
rect 28172 7540 28224 7546
rect 28172 7482 28224 7488
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 28184 6186 28212 7142
rect 28276 7041 28304 7686
rect 28262 7032 28318 7041
rect 28262 6967 28318 6976
rect 28368 6390 28396 13212
rect 28460 7478 28488 13262
rect 28552 12356 28580 14758
rect 28644 12434 28672 20198
rect 28736 19836 28764 20454
rect 29104 20330 29132 20878
rect 28816 20324 28868 20330
rect 28816 20266 28868 20272
rect 29092 20324 29144 20330
rect 29092 20266 29144 20272
rect 28828 20058 28856 20266
rect 28908 20256 28960 20262
rect 28908 20198 28960 20204
rect 29000 20256 29052 20262
rect 29000 20198 29052 20204
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28816 19848 28868 19854
rect 28736 19808 28816 19836
rect 28816 19790 28868 19796
rect 28828 19446 28856 19790
rect 28920 19718 28948 20198
rect 29012 19990 29040 20198
rect 29000 19984 29052 19990
rect 29000 19926 29052 19932
rect 29196 19922 29224 21286
rect 29472 20942 29500 21490
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29184 19916 29236 19922
rect 29184 19858 29236 19864
rect 29564 19786 29592 21490
rect 30116 20058 30144 21898
rect 31036 21690 31064 21966
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 30196 21072 30248 21078
rect 30196 21014 30248 21020
rect 30208 20058 30236 21014
rect 31220 20874 31248 21966
rect 31312 21622 31340 21966
rect 31956 21962 31984 22066
rect 32496 22034 32548 22040
rect 31852 21956 31904 21962
rect 31852 21898 31904 21904
rect 31944 21956 31996 21962
rect 31944 21898 31996 21904
rect 31300 21616 31352 21622
rect 31300 21558 31352 21564
rect 31864 21554 31892 21898
rect 31956 21622 31984 21898
rect 32508 21690 32536 22034
rect 32496 21684 32548 21690
rect 32496 21626 32548 21632
rect 31944 21616 31996 21622
rect 31944 21558 31996 21564
rect 31852 21548 31904 21554
rect 31852 21490 31904 21496
rect 31956 21010 31984 21558
rect 33324 21480 33376 21486
rect 33324 21422 33376 21428
rect 31944 21004 31996 21010
rect 31944 20946 31996 20952
rect 33048 21004 33100 21010
rect 33048 20946 33100 20952
rect 30380 20868 30432 20874
rect 30380 20810 30432 20816
rect 31208 20868 31260 20874
rect 31208 20810 31260 20816
rect 31668 20868 31720 20874
rect 31668 20810 31720 20816
rect 30104 20052 30156 20058
rect 30104 19994 30156 20000
rect 30196 20052 30248 20058
rect 30196 19994 30248 20000
rect 29736 19916 29788 19922
rect 29736 19858 29788 19864
rect 29552 19780 29604 19786
rect 29552 19722 29604 19728
rect 29644 19780 29696 19786
rect 29644 19722 29696 19728
rect 28908 19712 28960 19718
rect 28908 19654 28960 19660
rect 28816 19440 28868 19446
rect 28816 19382 28868 19388
rect 28828 18834 28856 19382
rect 28920 19378 28948 19654
rect 29564 19446 29592 19722
rect 29552 19440 29604 19446
rect 29552 19382 29604 19388
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 28816 18828 28868 18834
rect 28816 18770 28868 18776
rect 28920 18766 28948 19314
rect 29656 18766 29684 19722
rect 29748 19718 29776 19858
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 29644 18760 29696 18766
rect 29644 18702 29696 18708
rect 28920 17746 28948 18702
rect 28908 17740 28960 17746
rect 28908 17682 28960 17688
rect 29012 16794 29040 18702
rect 29748 18578 29776 19654
rect 30392 19242 30420 20810
rect 31680 20466 31708 20810
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 31760 20460 31812 20466
rect 31760 20402 31812 20408
rect 31772 19854 31800 20402
rect 31956 19854 31984 20946
rect 32772 20800 32824 20806
rect 32772 20742 32824 20748
rect 32680 20528 32732 20534
rect 32680 20470 32732 20476
rect 32034 19952 32090 19961
rect 32692 19922 32720 20470
rect 32034 19887 32090 19896
rect 32680 19916 32732 19922
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 31772 19334 31800 19790
rect 31772 19310 31892 19334
rect 31772 19306 31904 19310
rect 31852 19304 31904 19306
rect 31852 19246 31904 19252
rect 30380 19236 30432 19242
rect 30380 19178 30432 19184
rect 29656 18550 29776 18578
rect 30196 18624 30248 18630
rect 30196 18566 30248 18572
rect 29184 18352 29236 18358
rect 29184 18294 29236 18300
rect 29092 17672 29144 17678
rect 29092 17614 29144 17620
rect 29104 17202 29132 17614
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 29000 16788 29052 16794
rect 29000 16730 29052 16736
rect 29000 16584 29052 16590
rect 29000 16526 29052 16532
rect 28722 16416 28778 16425
rect 28722 16351 28778 16360
rect 28736 16046 28764 16351
rect 29012 16250 29040 16526
rect 29000 16244 29052 16250
rect 29000 16186 29052 16192
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 29012 15366 29040 16186
rect 29104 16114 29132 17138
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 29092 15428 29144 15434
rect 29092 15370 29144 15376
rect 29000 15360 29052 15366
rect 29000 15302 29052 15308
rect 29104 15026 29132 15370
rect 29092 15020 29144 15026
rect 29092 14962 29144 14968
rect 29196 12434 29224 18294
rect 29656 18290 29684 18550
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 29644 18284 29696 18290
rect 29644 18226 29696 18232
rect 29736 18284 29788 18290
rect 29736 18226 29788 18232
rect 30012 18284 30064 18290
rect 30012 18226 30064 18232
rect 29472 17678 29500 18226
rect 29748 17898 29776 18226
rect 29748 17870 29868 17898
rect 29736 17740 29788 17746
rect 29736 17682 29788 17688
rect 29460 17672 29512 17678
rect 29460 17614 29512 17620
rect 29460 17196 29512 17202
rect 29460 17138 29512 17144
rect 29552 17196 29604 17202
rect 29552 17138 29604 17144
rect 29274 16824 29330 16833
rect 29274 16759 29330 16768
rect 29288 16726 29316 16759
rect 29276 16720 29328 16726
rect 29276 16662 29328 16668
rect 29472 16454 29500 17138
rect 29460 16448 29512 16454
rect 29460 16390 29512 16396
rect 29276 15496 29328 15502
rect 29276 15438 29328 15444
rect 29288 15162 29316 15438
rect 29276 15156 29328 15162
rect 29276 15098 29328 15104
rect 29276 15020 29328 15026
rect 29276 14962 29328 14968
rect 29288 14929 29316 14962
rect 29274 14920 29330 14929
rect 29274 14855 29330 14864
rect 29288 14618 29316 14855
rect 29276 14612 29328 14618
rect 29276 14554 29328 14560
rect 29460 14408 29512 14414
rect 29460 14350 29512 14356
rect 29472 12442 29500 14350
rect 29460 12436 29512 12442
rect 28644 12406 28764 12434
rect 29196 12406 29408 12434
rect 28552 12328 28672 12356
rect 28540 12232 28592 12238
rect 28540 12174 28592 12180
rect 28552 11082 28580 12174
rect 28644 11830 28672 12328
rect 28632 11824 28684 11830
rect 28632 11766 28684 11772
rect 28632 11552 28684 11558
rect 28632 11494 28684 11500
rect 28644 11150 28672 11494
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 28540 11076 28592 11082
rect 28540 11018 28592 11024
rect 28632 9512 28684 9518
rect 28630 9480 28632 9489
rect 28684 9480 28686 9489
rect 28630 9415 28686 9424
rect 28540 8900 28592 8906
rect 28540 8842 28592 8848
rect 28552 8362 28580 8842
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28540 8356 28592 8362
rect 28540 8298 28592 8304
rect 28448 7472 28500 7478
rect 28448 7414 28500 7420
rect 28356 6384 28408 6390
rect 28356 6326 28408 6332
rect 28172 6180 28224 6186
rect 28172 6122 28224 6128
rect 28540 5908 28592 5914
rect 28540 5850 28592 5856
rect 28552 5710 28580 5850
rect 28540 5704 28592 5710
rect 28540 5646 28592 5652
rect 28644 5522 28672 8570
rect 28736 8566 28764 12406
rect 28908 12232 28960 12238
rect 28906 12200 28908 12209
rect 28960 12200 28962 12209
rect 28906 12135 28962 12144
rect 28816 12096 28868 12102
rect 28816 12038 28868 12044
rect 28828 11694 28856 12038
rect 28816 11688 28868 11694
rect 28816 11630 28868 11636
rect 29276 11688 29328 11694
rect 29276 11630 29328 11636
rect 29288 11121 29316 11630
rect 29274 11112 29330 11121
rect 29274 11047 29330 11056
rect 28816 9920 28868 9926
rect 28816 9862 28868 9868
rect 28828 9692 28856 9862
rect 28816 9686 28868 9692
rect 28816 9628 28868 9634
rect 28908 9686 28960 9692
rect 28908 9628 28960 9634
rect 28920 9518 28948 9628
rect 28908 9512 28960 9518
rect 28908 9454 28960 9460
rect 28908 9104 28960 9110
rect 28908 9046 28960 9052
rect 28920 8974 28948 9046
rect 28816 8968 28868 8974
rect 28816 8910 28868 8916
rect 28908 8968 28960 8974
rect 28908 8910 28960 8916
rect 28828 8566 28856 8910
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 28724 8560 28776 8566
rect 28724 8502 28776 8508
rect 28816 8560 28868 8566
rect 28816 8502 28868 8508
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 28736 7993 28764 8230
rect 28722 7984 28778 7993
rect 28722 7919 28778 7928
rect 28736 7206 28764 7919
rect 28828 7546 28856 8502
rect 28920 7750 28948 8774
rect 29000 8288 29052 8294
rect 28998 8256 29000 8265
rect 29052 8256 29054 8265
rect 28998 8191 29054 8200
rect 28908 7744 28960 7750
rect 28908 7686 28960 7692
rect 28816 7540 28868 7546
rect 28816 7482 28868 7488
rect 28920 7478 28948 7686
rect 28908 7472 28960 7478
rect 28908 7414 28960 7420
rect 29182 7304 29238 7313
rect 29182 7239 29238 7248
rect 29196 7206 29224 7239
rect 28724 7200 28776 7206
rect 28724 7142 28776 7148
rect 29092 7200 29144 7206
rect 29092 7142 29144 7148
rect 29184 7200 29236 7206
rect 29184 7142 29236 7148
rect 28724 6112 28776 6118
rect 28724 6054 28776 6060
rect 28908 6112 28960 6118
rect 28908 6054 28960 6060
rect 28736 5710 28764 6054
rect 28920 5914 28948 6054
rect 28908 5908 28960 5914
rect 28908 5850 28960 5856
rect 28724 5704 28776 5710
rect 28724 5646 28776 5652
rect 28644 5494 28856 5522
rect 28632 5024 28684 5030
rect 28632 4966 28684 4972
rect 28644 4214 28672 4966
rect 28632 4208 28684 4214
rect 28446 4176 28502 4185
rect 28632 4150 28684 4156
rect 28446 4111 28502 4120
rect 28264 4072 28316 4078
rect 28264 4014 28316 4020
rect 28172 3936 28224 3942
rect 28172 3878 28224 3884
rect 28184 3602 28212 3878
rect 28172 3596 28224 3602
rect 28172 3538 28224 3544
rect 27988 3392 28040 3398
rect 27988 3334 28040 3340
rect 28080 3392 28132 3398
rect 28080 3334 28132 3340
rect 27620 3120 27672 3126
rect 27620 3062 27672 3068
rect 28000 2774 28028 3334
rect 28276 3126 28304 4014
rect 28460 3942 28488 4111
rect 28448 3936 28500 3942
rect 28448 3878 28500 3884
rect 28264 3120 28316 3126
rect 28264 3062 28316 3068
rect 28000 2746 28120 2774
rect 28092 2446 28120 2746
rect 28828 2650 28856 5494
rect 28920 4758 28948 5850
rect 29000 5568 29052 5574
rect 29000 5510 29052 5516
rect 29012 5234 29040 5510
rect 29000 5228 29052 5234
rect 29000 5170 29052 5176
rect 28908 4752 28960 4758
rect 28908 4694 28960 4700
rect 29104 4690 29132 7142
rect 29092 4684 29144 4690
rect 29092 4626 29144 4632
rect 29380 2650 29408 12406
rect 29564 12434 29592 17138
rect 29644 16652 29696 16658
rect 29644 16594 29696 16600
rect 29656 16114 29684 16594
rect 29748 16590 29776 17682
rect 29840 17610 29868 17870
rect 30024 17678 30052 18226
rect 30012 17672 30064 17678
rect 30012 17614 30064 17620
rect 29828 17604 29880 17610
rect 29828 17546 29880 17552
rect 29920 17604 29972 17610
rect 29920 17546 29972 17552
rect 29840 17134 29868 17546
rect 29828 17128 29880 17134
rect 29828 17070 29880 17076
rect 29736 16584 29788 16590
rect 29736 16526 29788 16532
rect 29644 16108 29696 16114
rect 29644 16050 29696 16056
rect 29828 16108 29880 16114
rect 29828 16050 29880 16056
rect 29840 15434 29868 16050
rect 29828 15428 29880 15434
rect 29828 15370 29880 15376
rect 29828 15088 29880 15094
rect 29826 15056 29828 15065
rect 29880 15056 29882 15065
rect 29826 14991 29882 15000
rect 29828 14816 29880 14822
rect 29828 14758 29880 14764
rect 29840 14414 29868 14758
rect 29828 14408 29880 14414
rect 29828 14350 29880 14356
rect 29828 12436 29880 12442
rect 29564 12406 29684 12434
rect 29460 12378 29512 12384
rect 29472 12306 29500 12378
rect 29460 12300 29512 12306
rect 29460 12242 29512 12248
rect 29460 11688 29512 11694
rect 29458 11656 29460 11665
rect 29512 11656 29514 11665
rect 29458 11591 29514 11600
rect 29472 11082 29500 11591
rect 29552 11552 29604 11558
rect 29552 11494 29604 11500
rect 29564 11218 29592 11494
rect 29552 11212 29604 11218
rect 29552 11154 29604 11160
rect 29460 11076 29512 11082
rect 29460 11018 29512 11024
rect 29460 6384 29512 6390
rect 29460 6326 29512 6332
rect 29472 5710 29500 6326
rect 29460 5704 29512 5710
rect 29460 5646 29512 5652
rect 29472 3942 29500 5646
rect 29552 5636 29604 5642
rect 29552 5578 29604 5584
rect 29460 3936 29512 3942
rect 29460 3878 29512 3884
rect 28816 2644 28868 2650
rect 28816 2586 28868 2592
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29472 2514 29500 3878
rect 29564 2922 29592 5578
rect 29552 2916 29604 2922
rect 29552 2858 29604 2864
rect 29460 2508 29512 2514
rect 29460 2450 29512 2456
rect 29564 2446 29592 2858
rect 29656 2582 29684 12406
rect 29932 12434 29960 17546
rect 30024 17202 30052 17614
rect 30208 17542 30236 18566
rect 30392 18306 30420 19178
rect 30392 18278 30512 18306
rect 30380 18216 30432 18222
rect 30380 18158 30432 18164
rect 30392 17610 30420 18158
rect 30380 17604 30432 17610
rect 30380 17546 30432 17552
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30012 17196 30064 17202
rect 30064 17156 30144 17184
rect 30012 17138 30064 17144
rect 30116 16114 30144 17156
rect 30392 17134 30420 17546
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30288 16176 30340 16182
rect 30288 16118 30340 16124
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 30196 15428 30248 15434
rect 30196 15370 30248 15376
rect 30012 15360 30064 15366
rect 30012 15302 30064 15308
rect 30024 15162 30052 15302
rect 30012 15156 30064 15162
rect 30012 15098 30064 15104
rect 30208 14618 30236 15370
rect 30196 14612 30248 14618
rect 30196 14554 30248 14560
rect 29932 12406 30052 12434
rect 29828 12378 29880 12384
rect 29840 11694 29868 12378
rect 29920 11756 29972 11762
rect 29920 11698 29972 11704
rect 29828 11688 29880 11694
rect 29828 11630 29880 11636
rect 29840 11150 29868 11630
rect 29932 11218 29960 11698
rect 29920 11212 29972 11218
rect 29920 11154 29972 11160
rect 29828 11144 29880 11150
rect 29748 11092 29828 11098
rect 29748 11086 29880 11092
rect 29918 11112 29974 11121
rect 29748 11070 29868 11086
rect 29644 2576 29696 2582
rect 29644 2518 29696 2524
rect 29748 2446 29776 11070
rect 29918 11047 29920 11056
rect 29972 11047 29974 11056
rect 29920 11018 29972 11024
rect 29932 10674 29960 11018
rect 29920 10668 29972 10674
rect 29920 10610 29972 10616
rect 29920 7404 29972 7410
rect 29920 7346 29972 7352
rect 29932 7274 29960 7346
rect 29920 7268 29972 7274
rect 29920 7210 29972 7216
rect 29828 6112 29880 6118
rect 29828 6054 29880 6060
rect 29840 5234 29868 6054
rect 29920 5568 29972 5574
rect 29920 5510 29972 5516
rect 29932 5302 29960 5510
rect 29920 5296 29972 5302
rect 29920 5238 29972 5244
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 30024 4010 30052 12406
rect 30104 11620 30156 11626
rect 30104 11562 30156 11568
rect 30116 11150 30144 11562
rect 30104 11144 30156 11150
rect 30104 11086 30156 11092
rect 30196 9376 30248 9382
rect 30196 9318 30248 9324
rect 30208 8498 30236 9318
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 30116 5234 30144 7686
rect 30196 7540 30248 7546
rect 30196 7482 30248 7488
rect 30208 6866 30236 7482
rect 30196 6860 30248 6866
rect 30196 6802 30248 6808
rect 30104 5228 30156 5234
rect 30104 5170 30156 5176
rect 30012 4004 30064 4010
rect 30012 3946 30064 3952
rect 30300 2650 30328 16118
rect 30378 15056 30434 15065
rect 30484 15026 30512 18278
rect 31944 17332 31996 17338
rect 31944 17274 31996 17280
rect 31484 17128 31536 17134
rect 31484 17070 31536 17076
rect 31496 16590 31524 17070
rect 31956 16794 31984 17274
rect 31944 16788 31996 16794
rect 31944 16730 31996 16736
rect 31300 16584 31352 16590
rect 31300 16526 31352 16532
rect 31484 16584 31536 16590
rect 31484 16526 31536 16532
rect 31312 16046 31340 16526
rect 31392 16516 31444 16522
rect 31392 16458 31444 16464
rect 31300 16040 31352 16046
rect 31300 15982 31352 15988
rect 30932 15564 30984 15570
rect 30932 15506 30984 15512
rect 30944 15162 30972 15506
rect 30932 15156 30984 15162
rect 30932 15098 30984 15104
rect 30378 14991 30434 15000
rect 30472 15020 30524 15026
rect 30392 14958 30420 14991
rect 30472 14962 30524 14968
rect 30932 15020 30984 15026
rect 30932 14962 30984 14968
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30392 13734 30420 14894
rect 30484 14074 30512 14962
rect 30944 14929 30972 14962
rect 30930 14920 30986 14929
rect 30930 14855 30986 14864
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30380 13728 30432 13734
rect 30380 13670 30432 13676
rect 30484 13530 30512 14010
rect 30380 13524 30432 13530
rect 30380 13466 30432 13472
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30392 13410 30420 13466
rect 30392 13382 30512 13410
rect 30380 13320 30432 13326
rect 30380 13262 30432 13268
rect 30392 12714 30420 13262
rect 30380 12708 30432 12714
rect 30380 12650 30432 12656
rect 30484 8634 30512 13382
rect 30564 12912 30616 12918
rect 30564 12854 30616 12860
rect 30576 12714 30604 12854
rect 30564 12708 30616 12714
rect 30564 12650 30616 12656
rect 30840 12640 30892 12646
rect 30840 12582 30892 12588
rect 30852 11558 30880 12582
rect 31116 11756 31168 11762
rect 31116 11698 31168 11704
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 30748 10668 30800 10674
rect 30748 10610 30800 10616
rect 30760 9926 30788 10610
rect 30748 9920 30800 9926
rect 30748 9862 30800 9868
rect 30472 8628 30524 8634
rect 30472 8570 30524 8576
rect 30380 8356 30432 8362
rect 30380 8298 30432 8304
rect 30392 7274 30420 8298
rect 30472 7404 30524 7410
rect 30472 7346 30524 7352
rect 30380 7268 30432 7274
rect 30380 7210 30432 7216
rect 30484 5302 30512 7346
rect 30656 6928 30708 6934
rect 30654 6896 30656 6905
rect 30708 6896 30710 6905
rect 30654 6831 30710 6840
rect 30760 6610 30788 9862
rect 30852 9382 30880 11494
rect 30932 10056 30984 10062
rect 30932 9998 30984 10004
rect 30944 9722 30972 9998
rect 30932 9716 30984 9722
rect 30932 9658 30984 9664
rect 30840 9376 30892 9382
rect 30840 9318 30892 9324
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 30944 7478 30972 8434
rect 30932 7472 30984 7478
rect 30932 7414 30984 7420
rect 31128 7410 31156 11698
rect 31208 10532 31260 10538
rect 31208 10474 31260 10480
rect 31220 9722 31248 10474
rect 31208 9716 31260 9722
rect 31208 9658 31260 9664
rect 31116 7404 31168 7410
rect 31116 7346 31168 7352
rect 31128 6934 31156 7346
rect 31116 6928 31168 6934
rect 31116 6870 31168 6876
rect 30840 6724 30892 6730
rect 30840 6666 30892 6672
rect 30576 6582 30788 6610
rect 30472 5296 30524 5302
rect 30472 5238 30524 5244
rect 30576 3602 30604 6582
rect 30852 6254 30880 6666
rect 30840 6248 30892 6254
rect 30840 6190 30892 6196
rect 31116 5296 31168 5302
rect 31116 5238 31168 5244
rect 31128 3641 31156 5238
rect 31220 5030 31248 9658
rect 31298 8392 31354 8401
rect 31298 8327 31354 8336
rect 31312 6390 31340 8327
rect 31300 6384 31352 6390
rect 31300 6326 31352 6332
rect 31312 5642 31340 6326
rect 31300 5636 31352 5642
rect 31300 5578 31352 5584
rect 31312 5302 31340 5578
rect 31300 5296 31352 5302
rect 31300 5238 31352 5244
rect 31208 5024 31260 5030
rect 31208 4966 31260 4972
rect 31300 5024 31352 5030
rect 31300 4966 31352 4972
rect 31312 4486 31340 4966
rect 31300 4480 31352 4486
rect 31300 4422 31352 4428
rect 31114 3632 31170 3641
rect 30564 3596 30616 3602
rect 31114 3567 31170 3576
rect 30564 3538 30616 3544
rect 31128 3534 31156 3567
rect 31116 3528 31168 3534
rect 31300 3528 31352 3534
rect 31116 3470 31168 3476
rect 31298 3496 31300 3505
rect 31352 3496 31354 3505
rect 31298 3431 31354 3440
rect 30472 3392 30524 3398
rect 30472 3334 30524 3340
rect 30484 3126 30512 3334
rect 30472 3120 30524 3126
rect 30472 3062 30524 3068
rect 29828 2644 29880 2650
rect 29828 2586 29880 2592
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 27988 2304 28040 2310
rect 27988 2246 28040 2252
rect 28000 800 28028 2246
rect 28920 800 28948 2382
rect 29840 2378 29868 2586
rect 31404 2514 31432 16458
rect 31576 14000 31628 14006
rect 31576 13942 31628 13948
rect 31588 13002 31616 13942
rect 31852 13320 31904 13326
rect 31852 13262 31904 13268
rect 31668 13184 31720 13190
rect 31668 13126 31720 13132
rect 31496 12986 31616 13002
rect 31484 12980 31616 12986
rect 31536 12974 31616 12980
rect 31484 12922 31536 12928
rect 31588 12434 31616 12974
rect 31680 12918 31708 13126
rect 31668 12912 31720 12918
rect 31668 12854 31720 12860
rect 31864 12442 31892 13262
rect 31496 12406 31616 12434
rect 31852 12436 31904 12442
rect 31496 12238 31524 12406
rect 31852 12378 31904 12384
rect 31484 12232 31536 12238
rect 31484 12174 31536 12180
rect 31496 11762 31524 12174
rect 31484 11756 31536 11762
rect 31484 11698 31536 11704
rect 31484 10464 31536 10470
rect 31484 10406 31536 10412
rect 31496 9654 31524 10406
rect 31668 10124 31720 10130
rect 31668 10066 31720 10072
rect 31680 9674 31708 10066
rect 31484 9648 31536 9654
rect 31680 9646 31892 9674
rect 31484 9590 31536 9596
rect 31864 9518 31892 9646
rect 31852 9512 31904 9518
rect 31852 9454 31904 9460
rect 31864 7750 31892 9454
rect 31852 7744 31904 7750
rect 31852 7686 31904 7692
rect 31864 6254 31892 7686
rect 31852 6248 31904 6254
rect 31574 6216 31630 6225
rect 31852 6190 31904 6196
rect 31574 6151 31630 6160
rect 31588 5914 31616 6151
rect 31576 5908 31628 5914
rect 31576 5850 31628 5856
rect 31576 3936 31628 3942
rect 31576 3878 31628 3884
rect 31588 2854 31616 3878
rect 31864 3058 31892 6190
rect 31852 3052 31904 3058
rect 31852 2994 31904 3000
rect 31576 2848 31628 2854
rect 31576 2790 31628 2796
rect 32048 2774 32076 19887
rect 32680 19858 32732 19864
rect 32220 19712 32272 19718
rect 32220 19654 32272 19660
rect 32680 19712 32732 19718
rect 32680 19654 32732 19660
rect 32128 17536 32180 17542
rect 32128 17478 32180 17484
rect 32140 17202 32168 17478
rect 32128 17196 32180 17202
rect 32128 17138 32180 17144
rect 32128 14272 32180 14278
rect 32128 14214 32180 14220
rect 32140 12850 32168 14214
rect 32128 12844 32180 12850
rect 32128 12786 32180 12792
rect 32128 7812 32180 7818
rect 32128 7754 32180 7760
rect 32140 7546 32168 7754
rect 32128 7540 32180 7546
rect 32128 7482 32180 7488
rect 32128 5296 32180 5302
rect 32126 5264 32128 5273
rect 32180 5264 32182 5273
rect 32126 5199 32182 5208
rect 32128 4616 32180 4622
rect 32126 4584 32128 4593
rect 32180 4584 32182 4593
rect 32126 4519 32182 4528
rect 32126 3088 32182 3097
rect 32126 3023 32128 3032
rect 32180 3023 32182 3032
rect 32128 2994 32180 3000
rect 32232 2774 32260 19654
rect 32692 19378 32720 19654
rect 32496 19372 32548 19378
rect 32496 19314 32548 19320
rect 32680 19372 32732 19378
rect 32680 19314 32732 19320
rect 32404 18216 32456 18222
rect 32404 18158 32456 18164
rect 32416 17814 32444 18158
rect 32404 17808 32456 17814
rect 32404 17750 32456 17756
rect 32416 17610 32444 17750
rect 32404 17604 32456 17610
rect 32404 17546 32456 17552
rect 32312 16992 32364 16998
rect 32310 16960 32312 16969
rect 32364 16960 32366 16969
rect 32310 16895 32366 16904
rect 32508 15008 32536 19314
rect 32784 19242 32812 20742
rect 33060 20466 33088 20946
rect 33336 20942 33364 21422
rect 33324 20936 33376 20942
rect 33324 20878 33376 20884
rect 33140 20800 33192 20806
rect 33140 20742 33192 20748
rect 32956 20460 33008 20466
rect 32956 20402 33008 20408
rect 33048 20460 33100 20466
rect 33048 20402 33100 20408
rect 32968 20346 32996 20402
rect 32968 20318 33088 20346
rect 32864 19848 32916 19854
rect 32916 19808 32996 19836
rect 32864 19790 32916 19796
rect 32864 19712 32916 19718
rect 32864 19654 32916 19660
rect 32876 19446 32904 19654
rect 32864 19440 32916 19446
rect 32864 19382 32916 19388
rect 32588 19236 32640 19242
rect 32588 19178 32640 19184
rect 32772 19236 32824 19242
rect 32772 19178 32824 19184
rect 32600 18766 32628 19178
rect 32680 19168 32732 19174
rect 32680 19110 32732 19116
rect 32692 18970 32720 19110
rect 32680 18964 32732 18970
rect 32680 18906 32732 18912
rect 32588 18760 32640 18766
rect 32588 18702 32640 18708
rect 32600 17746 32628 18702
rect 32876 18698 32904 19382
rect 32968 19310 32996 19808
rect 33060 19718 33088 20318
rect 33048 19712 33100 19718
rect 33048 19654 33100 19660
rect 33060 19378 33088 19654
rect 33152 19514 33180 20742
rect 33232 20392 33284 20398
rect 33428 20346 33456 22714
rect 33520 22234 33548 23054
rect 33692 22432 33744 22438
rect 33692 22374 33744 22380
rect 33508 22228 33560 22234
rect 33508 22170 33560 22176
rect 33508 22024 33560 22030
rect 33508 21966 33560 21972
rect 33520 20942 33548 21966
rect 33704 21078 33732 22374
rect 33692 21072 33744 21078
rect 33692 21014 33744 21020
rect 33600 21004 33652 21010
rect 33600 20946 33652 20952
rect 33508 20936 33560 20942
rect 33508 20878 33560 20884
rect 33612 20534 33640 20946
rect 33692 20936 33744 20942
rect 33692 20878 33744 20884
rect 33704 20602 33732 20878
rect 33876 20868 33928 20874
rect 33876 20810 33928 20816
rect 33888 20602 33916 20810
rect 33692 20596 33744 20602
rect 33692 20538 33744 20544
rect 33876 20596 33928 20602
rect 33876 20538 33928 20544
rect 33600 20528 33652 20534
rect 33600 20470 33652 20476
rect 33232 20334 33284 20340
rect 33244 19961 33272 20334
rect 33336 20318 33456 20346
rect 33612 20330 33640 20470
rect 33600 20324 33652 20330
rect 33230 19952 33286 19961
rect 33230 19887 33286 19896
rect 33232 19780 33284 19786
rect 33232 19722 33284 19728
rect 33140 19508 33192 19514
rect 33140 19450 33192 19456
rect 33048 19372 33100 19378
rect 33048 19314 33100 19320
rect 32956 19304 33008 19310
rect 32956 19246 33008 19252
rect 33060 18766 33088 19314
rect 33048 18760 33100 18766
rect 32968 18720 33048 18748
rect 32864 18692 32916 18698
rect 32864 18634 32916 18640
rect 32876 18290 32904 18634
rect 32968 18358 32996 18720
rect 33048 18702 33100 18708
rect 33048 18624 33100 18630
rect 33048 18566 33100 18572
rect 32956 18352 33008 18358
rect 32956 18294 33008 18300
rect 32864 18284 32916 18290
rect 32864 18226 32916 18232
rect 32588 17740 32640 17746
rect 32588 17682 32640 17688
rect 32772 16448 32824 16454
rect 32772 16390 32824 16396
rect 32784 15910 32812 16390
rect 32956 16176 33008 16182
rect 32956 16118 33008 16124
rect 32864 16108 32916 16114
rect 32864 16050 32916 16056
rect 32772 15904 32824 15910
rect 32772 15846 32824 15852
rect 32784 15502 32812 15846
rect 32772 15496 32824 15502
rect 32772 15438 32824 15444
rect 32876 15162 32904 16050
rect 32864 15156 32916 15162
rect 32864 15098 32916 15104
rect 32508 14980 32812 15008
rect 32680 12844 32732 12850
rect 32680 12786 32732 12792
rect 32692 11762 32720 12786
rect 32680 11756 32732 11762
rect 32680 11698 32732 11704
rect 32692 9518 32720 11698
rect 32680 9512 32732 9518
rect 32680 9454 32732 9460
rect 32312 8356 32364 8362
rect 32312 8298 32364 8304
rect 32324 6798 32352 8298
rect 32588 8084 32640 8090
rect 32588 8026 32640 8032
rect 32600 7750 32628 8026
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 32588 7744 32640 7750
rect 32588 7686 32640 7692
rect 32692 7426 32720 7822
rect 32508 7398 32720 7426
rect 32508 6866 32536 7398
rect 32588 7336 32640 7342
rect 32588 7278 32640 7284
rect 32496 6860 32548 6866
rect 32496 6802 32548 6808
rect 32312 6792 32364 6798
rect 32312 6734 32364 6740
rect 32496 6724 32548 6730
rect 32496 6666 32548 6672
rect 32402 6080 32458 6089
rect 32402 6015 32458 6024
rect 32416 5710 32444 6015
rect 32508 5817 32536 6666
rect 32494 5808 32550 5817
rect 32494 5743 32550 5752
rect 32404 5704 32456 5710
rect 32404 5646 32456 5652
rect 32496 5636 32548 5642
rect 32496 5578 32548 5584
rect 32508 5545 32536 5578
rect 32494 5536 32550 5545
rect 32494 5471 32550 5480
rect 32312 5364 32364 5370
rect 32600 5352 32628 7278
rect 32680 6452 32732 6458
rect 32680 6394 32732 6400
rect 32692 5574 32720 6394
rect 32784 6202 32812 14980
rect 32968 14278 32996 16118
rect 32956 14272 33008 14278
rect 32956 14214 33008 14220
rect 32968 13938 32996 14214
rect 32956 13932 33008 13938
rect 32956 13874 33008 13880
rect 32956 8492 33008 8498
rect 32956 8434 33008 8440
rect 32968 7818 32996 8434
rect 32956 7812 33008 7818
rect 32956 7754 33008 7760
rect 32864 6656 32916 6662
rect 32864 6598 32916 6604
rect 32876 6390 32904 6598
rect 32864 6384 32916 6390
rect 32864 6326 32916 6332
rect 32784 6174 32904 6202
rect 32770 5944 32826 5953
rect 32770 5879 32826 5888
rect 32680 5568 32732 5574
rect 32680 5510 32732 5516
rect 32680 5364 32732 5370
rect 32600 5324 32680 5352
rect 32312 5306 32364 5312
rect 32680 5306 32732 5312
rect 32324 4622 32352 5306
rect 32496 5228 32548 5234
rect 32496 5170 32548 5176
rect 32312 4616 32364 4622
rect 32312 4558 32364 4564
rect 32508 4554 32536 5170
rect 32496 4548 32548 4554
rect 32496 4490 32548 4496
rect 32508 4457 32536 4490
rect 32588 4480 32640 4486
rect 32494 4448 32550 4457
rect 32588 4422 32640 4428
rect 32494 4383 32550 4392
rect 32600 4282 32628 4422
rect 32588 4276 32640 4282
rect 32588 4218 32640 4224
rect 31956 2746 32076 2774
rect 32140 2746 32260 2774
rect 31392 2508 31444 2514
rect 31392 2450 31444 2456
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 31852 2440 31904 2446
rect 31956 2417 31984 2746
rect 32140 2553 32168 2746
rect 32126 2544 32182 2553
rect 32126 2479 32182 2488
rect 31852 2382 31904 2388
rect 31942 2408 31998 2417
rect 29828 2372 29880 2378
rect 29828 2314 29880 2320
rect 29460 2304 29512 2310
rect 29460 2246 29512 2252
rect 29472 800 29500 2246
rect 30392 800 30420 2382
rect 30840 2304 30892 2310
rect 30840 2246 30892 2252
rect 30852 800 30880 2246
rect 31864 800 31892 2382
rect 31942 2343 31998 2352
rect 32312 2304 32364 2310
rect 32312 2246 32364 2252
rect 32324 800 32352 2246
rect 32784 2145 32812 5879
rect 32876 2650 32904 6174
rect 32968 5370 32996 7754
rect 33060 5953 33088 18566
rect 33140 18284 33192 18290
rect 33140 18226 33192 18232
rect 33152 17678 33180 18226
rect 33140 17672 33192 17678
rect 33140 17614 33192 17620
rect 33152 17202 33180 17614
rect 33140 17196 33192 17202
rect 33140 17138 33192 17144
rect 33152 16998 33180 17138
rect 33140 16992 33192 16998
rect 33140 16934 33192 16940
rect 33140 15020 33192 15026
rect 33140 14962 33192 14968
rect 33152 13394 33180 14962
rect 33140 13388 33192 13394
rect 33140 13330 33192 13336
rect 33140 9648 33192 9654
rect 33140 9590 33192 9596
rect 33152 9450 33180 9590
rect 33140 9444 33192 9450
rect 33140 9386 33192 9392
rect 33140 8288 33192 8294
rect 33140 8230 33192 8236
rect 33152 7342 33180 8230
rect 33140 7336 33192 7342
rect 33140 7278 33192 7284
rect 33140 6112 33192 6118
rect 33138 6080 33140 6089
rect 33192 6080 33194 6089
rect 33138 6015 33194 6024
rect 33046 5944 33102 5953
rect 33046 5879 33102 5888
rect 33048 5840 33100 5846
rect 33046 5808 33048 5817
rect 33100 5808 33102 5817
rect 33046 5743 33102 5752
rect 32956 5364 33008 5370
rect 32956 5306 33008 5312
rect 33140 5364 33192 5370
rect 33140 5306 33192 5312
rect 32956 5228 33008 5234
rect 32956 5170 33008 5176
rect 32968 4622 32996 5170
rect 32956 4616 33008 4622
rect 32956 4558 33008 4564
rect 33152 4146 33180 5306
rect 33140 4140 33192 4146
rect 33140 4082 33192 4088
rect 33046 3768 33102 3777
rect 33046 3703 33102 3712
rect 33060 3670 33088 3703
rect 33048 3664 33100 3670
rect 33048 3606 33100 3612
rect 33152 3602 33180 4082
rect 33140 3596 33192 3602
rect 33140 3538 33192 3544
rect 32864 2644 32916 2650
rect 32864 2586 32916 2592
rect 32770 2136 32826 2145
rect 32770 2071 32826 2080
rect 33244 1426 33272 19722
rect 33336 15026 33364 20318
rect 33600 20266 33652 20272
rect 33416 20256 33468 20262
rect 33416 20198 33468 20204
rect 33428 20058 33456 20198
rect 33416 20052 33468 20058
rect 33416 19994 33468 20000
rect 33704 19922 33732 20538
rect 34060 20256 34112 20262
rect 34060 20198 34112 20204
rect 33692 19916 33744 19922
rect 33692 19858 33744 19864
rect 34072 19378 34100 20198
rect 34060 19372 34112 19378
rect 34060 19314 34112 19320
rect 33692 19168 33744 19174
rect 33692 19110 33744 19116
rect 33704 18902 33732 19110
rect 33692 18896 33744 18902
rect 33692 18838 33744 18844
rect 33876 18420 33928 18426
rect 33980 18414 34192 18442
rect 33980 18408 34008 18414
rect 33928 18380 34008 18408
rect 33876 18362 33928 18368
rect 33600 18148 33652 18154
rect 33600 18090 33652 18096
rect 33508 17604 33560 17610
rect 33612 17592 33640 18090
rect 33888 17678 33916 18362
rect 34060 18352 34112 18358
rect 33980 18312 34060 18340
rect 33876 17672 33928 17678
rect 33876 17614 33928 17620
rect 33560 17564 33640 17592
rect 33508 17546 33560 17552
rect 33520 17270 33548 17546
rect 33508 17264 33560 17270
rect 33508 17206 33560 17212
rect 33888 17202 33916 17614
rect 33876 17196 33928 17202
rect 33876 17138 33928 17144
rect 33508 15360 33560 15366
rect 33508 15302 33560 15308
rect 33520 15094 33548 15302
rect 33508 15088 33560 15094
rect 33508 15030 33560 15036
rect 33324 15020 33376 15026
rect 33324 14962 33376 14968
rect 33336 14414 33364 14962
rect 33416 14884 33468 14890
rect 33416 14826 33468 14832
rect 33324 14408 33376 14414
rect 33324 14350 33376 14356
rect 33324 13932 33376 13938
rect 33324 13874 33376 13880
rect 33336 13530 33364 13874
rect 33324 13524 33376 13530
rect 33324 13466 33376 13472
rect 33324 13320 33376 13326
rect 33428 13308 33456 14826
rect 33376 13280 33456 13308
rect 33324 13262 33376 13268
rect 33336 13190 33364 13262
rect 33324 13184 33376 13190
rect 33324 13126 33376 13132
rect 33336 9654 33364 13126
rect 33508 12640 33560 12646
rect 33508 12582 33560 12588
rect 33520 11898 33548 12582
rect 33508 11892 33560 11898
rect 33508 11834 33560 11840
rect 33600 11892 33652 11898
rect 33600 11834 33652 11840
rect 33612 11626 33640 11834
rect 33600 11620 33652 11626
rect 33600 11562 33652 11568
rect 33784 11144 33836 11150
rect 33784 11086 33836 11092
rect 33324 9648 33376 9654
rect 33324 9590 33376 9596
rect 33600 9580 33652 9586
rect 33600 9522 33652 9528
rect 33612 9178 33640 9522
rect 33600 9172 33652 9178
rect 33600 9114 33652 9120
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 33508 8968 33560 8974
rect 33612 8945 33640 8978
rect 33508 8910 33560 8916
rect 33598 8936 33654 8945
rect 33520 8634 33548 8910
rect 33598 8871 33654 8880
rect 33692 8900 33744 8906
rect 33692 8842 33744 8848
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33324 8560 33376 8566
rect 33324 8502 33376 8508
rect 33336 8401 33364 8502
rect 33322 8392 33378 8401
rect 33322 8327 33378 8336
rect 33704 8294 33732 8842
rect 33692 8288 33744 8294
rect 33692 8230 33744 8236
rect 33324 8016 33376 8022
rect 33322 7984 33324 7993
rect 33376 7984 33378 7993
rect 33322 7919 33378 7928
rect 33336 6798 33364 7919
rect 33416 6860 33468 6866
rect 33416 6802 33468 6808
rect 33324 6792 33376 6798
rect 33324 6734 33376 6740
rect 33428 5778 33456 6802
rect 33600 6452 33652 6458
rect 33600 6394 33652 6400
rect 33416 5772 33468 5778
rect 33416 5714 33468 5720
rect 33612 5710 33640 6394
rect 33600 5704 33652 5710
rect 33600 5646 33652 5652
rect 33324 5568 33376 5574
rect 33322 5536 33324 5545
rect 33376 5536 33378 5545
rect 33322 5471 33378 5480
rect 33612 5273 33640 5646
rect 33598 5264 33654 5273
rect 33598 5199 33654 5208
rect 33322 4176 33378 4185
rect 33322 4111 33378 4120
rect 33508 4140 33560 4146
rect 33336 3738 33364 4111
rect 33508 4082 33560 4088
rect 33416 4004 33468 4010
rect 33416 3946 33468 3952
rect 33428 3738 33456 3946
rect 33324 3732 33376 3738
rect 33324 3674 33376 3680
rect 33416 3732 33468 3738
rect 33416 3674 33468 3680
rect 33416 3528 33468 3534
rect 33520 3516 33548 4082
rect 33468 3488 33548 3516
rect 33416 3470 33468 3476
rect 33324 3460 33376 3466
rect 33324 3402 33376 3408
rect 33336 3369 33364 3402
rect 33322 3360 33378 3369
rect 33322 3295 33378 3304
rect 33508 3188 33560 3194
rect 33508 3130 33560 3136
rect 33324 2508 33376 2514
rect 33324 2450 33376 2456
rect 33232 1420 33284 1426
rect 33232 1362 33284 1368
rect 33336 800 33364 2450
rect 33520 1494 33548 3130
rect 33612 2446 33640 5199
rect 33692 4072 33744 4078
rect 33692 4014 33744 4020
rect 33704 3398 33732 4014
rect 33796 3398 33824 11086
rect 33876 9172 33928 9178
rect 33876 9114 33928 9120
rect 33888 8974 33916 9114
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 33876 8628 33928 8634
rect 33876 8570 33928 8576
rect 33888 8430 33916 8570
rect 33876 8424 33928 8430
rect 33876 8366 33928 8372
rect 33876 7540 33928 7546
rect 33876 7482 33928 7488
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 33796 3194 33824 3334
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 33784 2848 33836 2854
rect 33784 2790 33836 2796
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 33508 1488 33560 1494
rect 33508 1430 33560 1436
rect 33796 800 33824 2790
rect 33888 1494 33916 7482
rect 33980 1970 34008 18312
rect 34060 18294 34112 18300
rect 34164 18290 34192 18414
rect 34152 18284 34204 18290
rect 34152 18226 34204 18232
rect 34060 14068 34112 14074
rect 34060 14010 34112 14016
rect 34072 13394 34100 14010
rect 34060 13388 34112 13394
rect 34060 13330 34112 13336
rect 34072 9654 34100 13330
rect 34152 11008 34204 11014
rect 34152 10950 34204 10956
rect 34060 9648 34112 9654
rect 34060 9590 34112 9596
rect 34060 8968 34112 8974
rect 34164 8956 34192 10950
rect 34256 8974 34284 39238
rect 50294 39196 50602 39216
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39120 50602 39140
rect 35808 39024 35860 39030
rect 35808 38966 35860 38972
rect 35716 38956 35768 38962
rect 35716 38898 35768 38904
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34428 22432 34480 22438
rect 34428 22374 34480 22380
rect 34440 22030 34468 22374
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35728 22094 35756 38898
rect 35544 22066 35756 22094
rect 34428 22024 34480 22030
rect 34428 21966 34480 21972
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 34808 20602 34836 21490
rect 35440 21344 35492 21350
rect 35440 21286 35492 21292
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35452 20942 35480 21286
rect 35440 20936 35492 20942
rect 35440 20878 35492 20884
rect 34796 20596 34848 20602
rect 34796 20538 34848 20544
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34704 20460 34756 20466
rect 34704 20402 34756 20408
rect 34532 19514 34560 20402
rect 34716 19990 34744 20402
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34704 19984 34756 19990
rect 34704 19926 34756 19932
rect 34520 19508 34572 19514
rect 34520 19450 34572 19456
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34440 18290 34468 19314
rect 35440 19304 35492 19310
rect 35440 19246 35492 19252
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 35452 18834 35480 19246
rect 35440 18828 35492 18834
rect 35440 18770 35492 18776
rect 35452 18426 35480 18770
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 35440 18420 35492 18426
rect 35440 18362 35492 18368
rect 34428 18284 34480 18290
rect 34428 18226 34480 18232
rect 34808 17678 34836 18362
rect 35452 18290 35480 18362
rect 35440 18284 35492 18290
rect 35440 18226 35492 18232
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34796 17672 34848 17678
rect 34796 17614 34848 17620
rect 34336 17604 34388 17610
rect 34336 17546 34388 17552
rect 34112 8928 34192 8956
rect 34244 8968 34296 8974
rect 34060 8910 34112 8916
rect 34244 8910 34296 8916
rect 34072 7993 34100 8910
rect 34058 7984 34114 7993
rect 34058 7919 34114 7928
rect 34348 7546 34376 17546
rect 34428 17264 34480 17270
rect 34428 17206 34480 17212
rect 34336 7540 34388 7546
rect 34336 7482 34388 7488
rect 34152 5296 34204 5302
rect 34152 5238 34204 5244
rect 34058 3768 34114 3777
rect 34058 3703 34114 3712
rect 34072 3670 34100 3703
rect 34060 3664 34112 3670
rect 34060 3606 34112 3612
rect 34060 3392 34112 3398
rect 34060 3334 34112 3340
rect 34072 3126 34100 3334
rect 34164 3194 34192 5238
rect 34336 3460 34388 3466
rect 34336 3402 34388 3408
rect 34348 3369 34376 3402
rect 34334 3360 34390 3369
rect 34334 3295 34390 3304
rect 34152 3188 34204 3194
rect 34152 3130 34204 3136
rect 34060 3120 34112 3126
rect 34060 3062 34112 3068
rect 34334 3088 34390 3097
rect 34334 3023 34336 3032
rect 34388 3023 34390 3032
rect 34336 2994 34388 3000
rect 34334 2952 34390 2961
rect 34334 2887 34336 2896
rect 34388 2887 34390 2896
rect 34336 2858 34388 2864
rect 34440 2774 34468 17206
rect 34612 17128 34664 17134
rect 34612 17070 34664 17076
rect 34624 13802 34652 17070
rect 34808 16590 34836 17614
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 35544 16810 35572 22066
rect 35716 20936 35768 20942
rect 35716 20878 35768 20884
rect 35728 20806 35756 20878
rect 35716 20800 35768 20806
rect 35716 20742 35768 20748
rect 35820 17354 35848 38966
rect 50294 38108 50602 38128
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38032 50602 38052
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 37648 20936 37700 20942
rect 37648 20878 37700 20884
rect 37372 20800 37424 20806
rect 37372 20742 37424 20748
rect 37464 20800 37516 20806
rect 37464 20742 37516 20748
rect 37384 20534 37412 20742
rect 37372 20528 37424 20534
rect 37372 20470 37424 20476
rect 37476 20058 37504 20742
rect 37660 20058 37688 20878
rect 37740 20868 37792 20874
rect 37740 20810 37792 20816
rect 37752 20534 37780 20810
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 37740 20528 37792 20534
rect 37740 20470 37792 20476
rect 37464 20052 37516 20058
rect 37464 19994 37516 20000
rect 37648 20052 37700 20058
rect 37648 19994 37700 20000
rect 37752 19938 37780 20470
rect 38016 20256 38068 20262
rect 38016 20198 38068 20204
rect 37752 19910 37872 19938
rect 36912 19848 36964 19854
rect 36912 19790 36964 19796
rect 37740 19848 37792 19854
rect 37740 19790 37792 19796
rect 36924 18766 36952 19790
rect 37752 19446 37780 19790
rect 37740 19440 37792 19446
rect 37740 19382 37792 19388
rect 37280 18964 37332 18970
rect 37280 18906 37332 18912
rect 36636 18760 36688 18766
rect 36636 18702 36688 18708
rect 36912 18760 36964 18766
rect 36912 18702 36964 18708
rect 37188 18760 37240 18766
rect 37188 18702 37240 18708
rect 36648 18358 36676 18702
rect 36636 18352 36688 18358
rect 36636 18294 36688 18300
rect 35900 18148 35952 18154
rect 35900 18090 35952 18096
rect 35452 16782 35572 16810
rect 35636 17326 35848 17354
rect 35912 17338 35940 18090
rect 36084 18080 36136 18086
rect 36084 18022 36136 18028
rect 36544 18080 36596 18086
rect 36544 18022 36596 18028
rect 36096 17338 36124 18022
rect 36268 17536 36320 17542
rect 36268 17478 36320 17484
rect 35900 17332 35952 17338
rect 34796 16584 34848 16590
rect 34796 16526 34848 16532
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34704 14544 34756 14550
rect 34704 14486 34756 14492
rect 34612 13796 34664 13802
rect 34612 13738 34664 13744
rect 34520 13456 34572 13462
rect 34520 13398 34572 13404
rect 34532 12238 34560 13398
rect 34624 13258 34652 13738
rect 34612 13252 34664 13258
rect 34612 13194 34664 13200
rect 34716 12434 34744 14486
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 35452 12918 35480 16782
rect 35532 16652 35584 16658
rect 35532 16594 35584 16600
rect 35544 14550 35572 16594
rect 35532 14544 35584 14550
rect 35532 14486 35584 14492
rect 35440 12912 35492 12918
rect 35440 12854 35492 12860
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34624 12406 34744 12434
rect 34520 12232 34572 12238
rect 34520 12174 34572 12180
rect 34624 7154 34652 12406
rect 35636 12102 35664 17326
rect 35900 17274 35952 17280
rect 36084 17332 36136 17338
rect 36084 17274 36136 17280
rect 36096 16572 36124 17274
rect 36280 16590 36308 17478
rect 36452 17264 36504 17270
rect 36452 17206 36504 17212
rect 36464 16726 36492 17206
rect 36556 16998 36584 18022
rect 36924 17746 36952 18702
rect 37200 18290 37228 18702
rect 37188 18284 37240 18290
rect 37188 18226 37240 18232
rect 37004 18216 37056 18222
rect 37004 18158 37056 18164
rect 36912 17740 36964 17746
rect 36912 17682 36964 17688
rect 37016 17678 37044 18158
rect 36728 17672 36780 17678
rect 36728 17614 36780 17620
rect 37004 17672 37056 17678
rect 37004 17614 37056 17620
rect 36636 17196 36688 17202
rect 36636 17138 36688 17144
rect 36544 16992 36596 16998
rect 36544 16934 36596 16940
rect 36452 16720 36504 16726
rect 36452 16662 36504 16668
rect 36173 16584 36225 16590
rect 36096 16544 36173 16572
rect 36173 16526 36225 16532
rect 36268 16584 36320 16590
rect 36268 16526 36320 16532
rect 35808 16448 35860 16454
rect 35808 16390 35860 16396
rect 35820 16182 35848 16390
rect 35808 16176 35860 16182
rect 35808 16118 35860 16124
rect 36452 14884 36504 14890
rect 36452 14826 36504 14832
rect 36360 14340 36412 14346
rect 36360 14282 36412 14288
rect 36372 14006 36400 14282
rect 36464 14074 36492 14826
rect 36648 14618 36676 17138
rect 36740 16250 36768 17614
rect 37016 16454 37044 17614
rect 37200 17542 37228 18226
rect 37292 18222 37320 18906
rect 37280 18216 37332 18222
rect 37280 18158 37332 18164
rect 37292 17814 37320 18158
rect 37280 17808 37332 17814
rect 37280 17750 37332 17756
rect 37188 17536 37240 17542
rect 37188 17478 37240 17484
rect 37556 17536 37608 17542
rect 37556 17478 37608 17484
rect 37096 16992 37148 16998
rect 37096 16934 37148 16940
rect 37108 16590 37136 16934
rect 37372 16788 37424 16794
rect 37372 16730 37424 16736
rect 37096 16584 37148 16590
rect 37096 16526 37148 16532
rect 37004 16448 37056 16454
rect 37004 16390 37056 16396
rect 36728 16244 36780 16250
rect 36728 16186 36780 16192
rect 36636 14612 36688 14618
rect 36636 14554 36688 14560
rect 36544 14340 36596 14346
rect 36544 14282 36596 14288
rect 36452 14068 36504 14074
rect 36452 14010 36504 14016
rect 36360 14000 36412 14006
rect 36360 13942 36412 13948
rect 36176 13864 36228 13870
rect 36176 13806 36228 13812
rect 35992 12844 36044 12850
rect 35992 12786 36044 12792
rect 35900 12776 35952 12782
rect 35900 12718 35952 12724
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 35624 12096 35676 12102
rect 35624 12038 35676 12044
rect 34808 11354 34836 12038
rect 35912 11626 35940 12718
rect 36004 12238 36032 12786
rect 36188 12434 36216 13806
rect 36556 13326 36584 14282
rect 36648 13802 36676 14554
rect 36728 14340 36780 14346
rect 36728 14282 36780 14288
rect 36740 13870 36768 14282
rect 36728 13864 36780 13870
rect 36728 13806 36780 13812
rect 36912 13864 36964 13870
rect 36912 13806 36964 13812
rect 36636 13796 36688 13802
rect 36636 13738 36688 13744
rect 36648 13530 36676 13738
rect 36636 13524 36688 13530
rect 36636 13466 36688 13472
rect 36544 13320 36596 13326
rect 36544 13262 36596 13268
rect 36188 12406 36400 12434
rect 35992 12232 36044 12238
rect 35992 12174 36044 12180
rect 36372 11762 36400 12406
rect 36636 12300 36688 12306
rect 36636 12242 36688 12248
rect 36452 12164 36504 12170
rect 36452 12106 36504 12112
rect 36176 11756 36228 11762
rect 36176 11698 36228 11704
rect 36360 11756 36412 11762
rect 36360 11698 36412 11704
rect 35990 11656 36046 11665
rect 35900 11620 35952 11626
rect 35990 11591 35992 11600
rect 35900 11562 35952 11568
rect 36044 11591 36046 11600
rect 35992 11562 36044 11568
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 36188 11354 36216 11698
rect 34796 11348 34848 11354
rect 34796 11290 34848 11296
rect 35440 11348 35492 11354
rect 35440 11290 35492 11296
rect 36176 11348 36228 11354
rect 36176 11290 36228 11296
rect 35072 11280 35124 11286
rect 35070 11248 35072 11257
rect 35124 11248 35126 11257
rect 35070 11183 35126 11192
rect 35452 11014 35480 11290
rect 36174 11248 36230 11257
rect 36174 11183 36230 11192
rect 36188 11150 36216 11183
rect 36176 11144 36228 11150
rect 35728 11082 36124 11098
rect 36176 11086 36228 11092
rect 36372 11082 36400 11698
rect 35728 11076 36136 11082
rect 35728 11070 36084 11076
rect 35728 11014 35756 11070
rect 36084 11018 36136 11024
rect 36360 11076 36412 11082
rect 36360 11018 36412 11024
rect 35440 11008 35492 11014
rect 35440 10950 35492 10956
rect 35716 11008 35768 11014
rect 35716 10950 35768 10956
rect 36176 11008 36228 11014
rect 36176 10950 36228 10956
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 36188 9382 36216 10950
rect 36464 10062 36492 12106
rect 36544 12096 36596 12102
rect 36544 12038 36596 12044
rect 36556 11762 36584 12038
rect 36544 11756 36596 11762
rect 36544 11698 36596 11704
rect 36544 11552 36596 11558
rect 36544 11494 36596 11500
rect 36556 11218 36584 11494
rect 36544 11212 36596 11218
rect 36544 11154 36596 11160
rect 36544 11008 36596 11014
rect 36544 10950 36596 10956
rect 36452 10056 36504 10062
rect 36452 9998 36504 10004
rect 36556 9994 36584 10950
rect 36544 9988 36596 9994
rect 36544 9930 36596 9936
rect 36452 9920 36504 9926
rect 36452 9862 36504 9868
rect 35348 9376 35400 9382
rect 35348 9318 35400 9324
rect 35808 9376 35860 9382
rect 35808 9318 35860 9324
rect 36176 9376 36228 9382
rect 36176 9318 36228 9324
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34796 8832 34848 8838
rect 34796 8774 34848 8780
rect 34808 8022 34836 8774
rect 35360 8430 35388 9318
rect 35532 8900 35584 8906
rect 35532 8842 35584 8848
rect 35348 8424 35400 8430
rect 35348 8366 35400 8372
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34796 8016 34848 8022
rect 34796 7958 34848 7964
rect 35072 7880 35124 7886
rect 35072 7822 35124 7828
rect 34796 7812 34848 7818
rect 34796 7754 34848 7760
rect 34532 7126 34652 7154
rect 34532 7002 34560 7126
rect 34808 7002 34836 7754
rect 34886 7440 34942 7449
rect 35084 7410 35112 7822
rect 35256 7744 35308 7750
rect 35256 7686 35308 7692
rect 35268 7410 35296 7686
rect 34886 7375 34888 7384
rect 34940 7375 34942 7384
rect 35072 7404 35124 7410
rect 34888 7346 34940 7352
rect 35072 7346 35124 7352
rect 35256 7404 35308 7410
rect 35256 7346 35308 7352
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34520 6996 34572 7002
rect 34520 6938 34572 6944
rect 34796 6996 34848 7002
rect 34796 6938 34848 6944
rect 34704 6792 34756 6798
rect 34704 6734 34756 6740
rect 34716 5166 34744 6734
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34704 5160 34756 5166
rect 34624 5120 34704 5148
rect 34520 5024 34572 5030
rect 34520 4966 34572 4972
rect 34532 4690 34560 4966
rect 34520 4684 34572 4690
rect 34520 4626 34572 4632
rect 34520 4140 34572 4146
rect 34520 4082 34572 4088
rect 34532 4049 34560 4082
rect 34518 4040 34574 4049
rect 34518 3975 34574 3984
rect 34624 3097 34652 5120
rect 34704 5102 34756 5108
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34702 4312 34758 4321
rect 34702 4247 34758 4256
rect 34716 4146 34744 4247
rect 34704 4140 34756 4146
rect 34704 4082 34756 4088
rect 34704 3936 34756 3942
rect 34704 3878 34756 3884
rect 34716 3126 34744 3878
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35360 3534 35388 8366
rect 35440 8288 35492 8294
rect 35440 8230 35492 8236
rect 35452 7886 35480 8230
rect 35544 8022 35572 8842
rect 35820 8294 35848 9318
rect 36266 9072 36322 9081
rect 36266 9007 36322 9016
rect 36280 8974 36308 9007
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 36360 8832 36412 8838
rect 36360 8774 36412 8780
rect 36372 8362 36400 8774
rect 36360 8356 36412 8362
rect 36360 8298 36412 8304
rect 35808 8288 35860 8294
rect 35808 8230 35860 8236
rect 35532 8016 35584 8022
rect 35532 7958 35584 7964
rect 35440 7880 35492 7886
rect 35440 7822 35492 7828
rect 35532 7744 35584 7750
rect 35532 7686 35584 7692
rect 35440 4548 35492 4554
rect 35440 4490 35492 4496
rect 35452 4078 35480 4490
rect 35544 4214 35572 7686
rect 36176 7404 36228 7410
rect 36176 7346 36228 7352
rect 35624 7200 35676 7206
rect 35624 7142 35676 7148
rect 35636 6798 35664 7142
rect 35808 6996 35860 7002
rect 35808 6938 35860 6944
rect 35624 6792 35676 6798
rect 35624 6734 35676 6740
rect 35820 5778 35848 6938
rect 36188 6662 36216 7346
rect 36176 6656 36228 6662
rect 36176 6598 36228 6604
rect 36188 6304 36216 6598
rect 36268 6316 36320 6322
rect 36096 6276 36268 6304
rect 35808 5772 35860 5778
rect 35808 5714 35860 5720
rect 35716 5568 35768 5574
rect 35820 5556 35848 5714
rect 35768 5528 35848 5556
rect 35900 5568 35952 5574
rect 35716 5510 35768 5516
rect 35900 5510 35952 5516
rect 35912 5234 35940 5510
rect 35992 5364 36044 5370
rect 35992 5306 36044 5312
rect 35900 5228 35952 5234
rect 35900 5170 35952 5176
rect 35622 4720 35678 4729
rect 35622 4655 35678 4664
rect 35636 4622 35664 4655
rect 36004 4622 36032 5306
rect 35624 4616 35676 4622
rect 35624 4558 35676 4564
rect 35992 4616 36044 4622
rect 35992 4558 36044 4564
rect 35532 4208 35584 4214
rect 35532 4150 35584 4156
rect 35440 4072 35492 4078
rect 35440 4014 35492 4020
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35348 3528 35400 3534
rect 35348 3470 35400 3476
rect 34704 3120 34756 3126
rect 34610 3088 34666 3097
rect 34704 3062 34756 3068
rect 34610 3023 34666 3032
rect 34256 2746 34468 2774
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 34164 2106 34192 2382
rect 34256 2106 34284 2746
rect 34152 2100 34204 2106
rect 34152 2042 34204 2048
rect 34244 2100 34296 2106
rect 34244 2042 34296 2048
rect 33968 1964 34020 1970
rect 33968 1906 34020 1912
rect 33876 1488 33928 1494
rect 33876 1430 33928 1436
rect 34808 800 34836 3470
rect 35348 3392 35400 3398
rect 35348 3334 35400 3340
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35164 2576 35216 2582
rect 35070 2544 35126 2553
rect 35164 2518 35216 2524
rect 35070 2479 35072 2488
rect 35124 2479 35126 2488
rect 35072 2450 35124 2456
rect 35176 2417 35204 2518
rect 35162 2408 35218 2417
rect 35162 2343 35218 2352
rect 35360 898 35388 3334
rect 35452 3058 35480 4014
rect 35544 3738 35572 4150
rect 35636 4146 35664 4558
rect 35808 4276 35860 4282
rect 35808 4218 35860 4224
rect 35624 4140 35676 4146
rect 35624 4082 35676 4088
rect 35532 3732 35584 3738
rect 35532 3674 35584 3680
rect 35544 3602 35572 3674
rect 35532 3596 35584 3602
rect 35532 3538 35584 3544
rect 35820 3194 35848 4218
rect 36096 4185 36124 6276
rect 36268 6258 36320 6264
rect 36372 6254 36400 8298
rect 36360 6248 36412 6254
rect 36358 6216 36360 6225
rect 36412 6216 36414 6225
rect 36358 6151 36414 6160
rect 36464 5710 36492 9862
rect 36556 9586 36584 9930
rect 36544 9580 36596 9586
rect 36544 9522 36596 9528
rect 36556 8498 36584 9522
rect 36648 8974 36676 12242
rect 36728 12232 36780 12238
rect 36780 12192 36860 12220
rect 36728 12174 36780 12180
rect 36832 11354 36860 12192
rect 36924 12170 36952 13806
rect 37280 12368 37332 12374
rect 37280 12310 37332 12316
rect 36912 12164 36964 12170
rect 36912 12106 36964 12112
rect 37096 11892 37148 11898
rect 37096 11834 37148 11840
rect 36820 11348 36872 11354
rect 36820 11290 36872 11296
rect 36832 11150 36860 11290
rect 36820 11144 36872 11150
rect 36820 11086 36872 11092
rect 37108 11082 37136 11834
rect 37096 11076 37148 11082
rect 37096 11018 37148 11024
rect 36820 9648 36872 9654
rect 36820 9590 36872 9596
rect 36832 9382 36860 9590
rect 36728 9376 36780 9382
rect 36728 9318 36780 9324
rect 36820 9376 36872 9382
rect 36820 9318 36872 9324
rect 36636 8968 36688 8974
rect 36636 8910 36688 8916
rect 36634 8528 36690 8537
rect 36544 8492 36596 8498
rect 36634 8463 36690 8472
rect 36544 8434 36596 8440
rect 36648 7449 36676 8463
rect 36634 7440 36690 7449
rect 36634 7375 36690 7384
rect 36648 7018 36676 7375
rect 36556 6990 36676 7018
rect 36556 6798 36584 6990
rect 36634 6896 36690 6905
rect 36634 6831 36690 6840
rect 36544 6792 36596 6798
rect 36544 6734 36596 6740
rect 36648 6254 36676 6831
rect 36636 6248 36688 6254
rect 36636 6190 36688 6196
rect 36268 5704 36320 5710
rect 36268 5646 36320 5652
rect 36452 5704 36504 5710
rect 36452 5646 36504 5652
rect 36176 5160 36228 5166
rect 36176 5102 36228 5108
rect 36188 5030 36216 5102
rect 36176 5024 36228 5030
rect 36176 4966 36228 4972
rect 36176 4616 36228 4622
rect 36176 4558 36228 4564
rect 36082 4176 36138 4185
rect 36188 4146 36216 4558
rect 36280 4486 36308 5646
rect 36464 5166 36492 5646
rect 36452 5160 36504 5166
rect 36452 5102 36504 5108
rect 36464 4554 36492 5102
rect 36740 4622 36768 9318
rect 36832 8430 36860 9318
rect 37002 8936 37058 8945
rect 37002 8871 37004 8880
rect 37056 8871 37058 8880
rect 37004 8842 37056 8848
rect 36912 8832 36964 8838
rect 36912 8774 36964 8780
rect 36820 8424 36872 8430
rect 36820 8366 36872 8372
rect 36924 7478 36952 8774
rect 37108 8537 37136 11018
rect 37292 9994 37320 12310
rect 37188 9988 37240 9994
rect 37188 9930 37240 9936
rect 37280 9988 37332 9994
rect 37280 9930 37332 9936
rect 37200 8974 37228 9930
rect 37292 9586 37320 9930
rect 37280 9580 37332 9586
rect 37280 9522 37332 9528
rect 37384 9178 37412 16730
rect 37568 16658 37596 17478
rect 37556 16652 37608 16658
rect 37556 16594 37608 16600
rect 37568 16114 37596 16594
rect 37556 16108 37608 16114
rect 37556 16050 37608 16056
rect 37568 14482 37596 16050
rect 37752 14550 37780 19382
rect 37844 18902 37872 19910
rect 38028 19310 38056 20198
rect 38292 19848 38344 19854
rect 38292 19790 38344 19796
rect 38304 19310 38332 19790
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 44088 19372 44140 19378
rect 44088 19314 44140 19320
rect 38016 19304 38068 19310
rect 38016 19246 38068 19252
rect 38292 19304 38344 19310
rect 38292 19246 38344 19252
rect 37832 18896 37884 18902
rect 37832 18838 37884 18844
rect 38304 18630 38332 19246
rect 43904 19168 43956 19174
rect 43904 19110 43956 19116
rect 38568 18896 38620 18902
rect 38568 18838 38620 18844
rect 37832 18624 37884 18630
rect 37832 18566 37884 18572
rect 38292 18624 38344 18630
rect 38292 18566 38344 18572
rect 37844 17746 37872 18566
rect 37832 17740 37884 17746
rect 37832 17682 37884 17688
rect 38016 17672 38068 17678
rect 38016 17614 38068 17620
rect 38200 17672 38252 17678
rect 38200 17614 38252 17620
rect 37832 15088 37884 15094
rect 37832 15030 37884 15036
rect 37740 14544 37792 14550
rect 37740 14486 37792 14492
rect 37556 14476 37608 14482
rect 37556 14418 37608 14424
rect 37568 12850 37596 14418
rect 37752 14278 37780 14486
rect 37844 14414 37872 15030
rect 37832 14408 37884 14414
rect 37832 14350 37884 14356
rect 37740 14272 37792 14278
rect 37740 14214 37792 14220
rect 37844 14074 37872 14350
rect 37832 14068 37884 14074
rect 37832 14010 37884 14016
rect 37924 13728 37976 13734
rect 37924 13670 37976 13676
rect 37556 12844 37608 12850
rect 37556 12786 37608 12792
rect 37648 10056 37700 10062
rect 37648 9998 37700 10004
rect 37464 9920 37516 9926
rect 37464 9862 37516 9868
rect 37372 9172 37424 9178
rect 37372 9114 37424 9120
rect 37476 9042 37504 9862
rect 37660 9654 37688 9998
rect 37936 9994 37964 13670
rect 38028 13530 38056 17614
rect 38212 16794 38240 17614
rect 38304 17610 38332 18566
rect 38580 17678 38608 18838
rect 43916 18766 43944 19110
rect 43076 18760 43128 18766
rect 43076 18702 43128 18708
rect 43904 18760 43956 18766
rect 43904 18702 43956 18708
rect 39212 18692 39264 18698
rect 39212 18634 39264 18640
rect 38936 18624 38988 18630
rect 38936 18566 38988 18572
rect 38948 17746 38976 18566
rect 39224 17882 39252 18634
rect 42616 18352 42668 18358
rect 42616 18294 42668 18300
rect 39212 17876 39264 17882
rect 39212 17818 39264 17824
rect 38936 17740 38988 17746
rect 38936 17682 38988 17688
rect 42628 17678 42656 18294
rect 43088 18290 43116 18702
rect 44100 18426 44128 19314
rect 47492 18760 47544 18766
rect 47492 18702 47544 18708
rect 44364 18624 44416 18630
rect 44364 18566 44416 18572
rect 47308 18624 47360 18630
rect 47308 18566 47360 18572
rect 43168 18420 43220 18426
rect 43168 18362 43220 18368
rect 44088 18420 44140 18426
rect 44088 18362 44140 18368
rect 43076 18284 43128 18290
rect 43076 18226 43128 18232
rect 43088 17882 43116 18226
rect 43076 17876 43128 17882
rect 43076 17818 43128 17824
rect 42800 17808 42852 17814
rect 42800 17750 42852 17756
rect 38568 17672 38620 17678
rect 38568 17614 38620 17620
rect 42616 17672 42668 17678
rect 42616 17614 42668 17620
rect 38292 17604 38344 17610
rect 38292 17546 38344 17552
rect 42156 17536 42208 17542
rect 42156 17478 42208 17484
rect 42524 17536 42576 17542
rect 42524 17478 42576 17484
rect 42168 17202 42196 17478
rect 42536 17338 42564 17478
rect 42524 17332 42576 17338
rect 42524 17274 42576 17280
rect 41696 17196 41748 17202
rect 41696 17138 41748 17144
rect 42156 17196 42208 17202
rect 42156 17138 42208 17144
rect 38200 16788 38252 16794
rect 38200 16730 38252 16736
rect 41708 16590 41736 17138
rect 42536 16658 42564 17274
rect 42524 16652 42576 16658
rect 42524 16594 42576 16600
rect 38752 16584 38804 16590
rect 38752 16526 38804 16532
rect 41696 16584 41748 16590
rect 41696 16526 41748 16532
rect 42248 16584 42300 16590
rect 42248 16526 42300 16532
rect 38476 14816 38528 14822
rect 38476 14758 38528 14764
rect 38660 14816 38712 14822
rect 38660 14758 38712 14764
rect 38488 14414 38516 14758
rect 38672 14618 38700 14758
rect 38660 14612 38712 14618
rect 38660 14554 38712 14560
rect 38476 14408 38528 14414
rect 38476 14350 38528 14356
rect 38568 14068 38620 14074
rect 38568 14010 38620 14016
rect 38384 14000 38436 14006
rect 38476 14000 38528 14006
rect 38436 13960 38476 13988
rect 38384 13942 38436 13948
rect 38476 13942 38528 13948
rect 38580 13938 38608 14010
rect 38764 13938 38792 16526
rect 40316 16108 40368 16114
rect 40316 16050 40368 16056
rect 40408 16108 40460 16114
rect 40408 16050 40460 16056
rect 38936 15156 38988 15162
rect 38936 15098 38988 15104
rect 38844 15020 38896 15026
rect 38844 14962 38896 14968
rect 38856 14074 38884 14962
rect 38948 14958 38976 15098
rect 40328 15026 40356 16050
rect 40420 15434 40448 16050
rect 41512 15632 41564 15638
rect 41512 15574 41564 15580
rect 40408 15428 40460 15434
rect 40408 15370 40460 15376
rect 41524 15162 41552 15574
rect 42260 15434 42288 16526
rect 42524 16448 42576 16454
rect 42524 16390 42576 16396
rect 42536 15570 42564 16390
rect 42628 16250 42656 17614
rect 42616 16244 42668 16250
rect 42616 16186 42668 16192
rect 42524 15564 42576 15570
rect 42352 15524 42524 15552
rect 42248 15428 42300 15434
rect 42248 15370 42300 15376
rect 41512 15156 41564 15162
rect 41512 15098 41564 15104
rect 41052 15088 41104 15094
rect 41052 15030 41104 15036
rect 40316 15020 40368 15026
rect 40316 14962 40368 14968
rect 38936 14952 38988 14958
rect 38936 14894 38988 14900
rect 38844 14068 38896 14074
rect 38844 14010 38896 14016
rect 38568 13932 38620 13938
rect 38568 13874 38620 13880
rect 38752 13932 38804 13938
rect 38752 13874 38804 13880
rect 38016 13524 38068 13530
rect 38016 13466 38068 13472
rect 38476 13524 38528 13530
rect 38476 13466 38528 13472
rect 38014 12336 38070 12345
rect 38014 12271 38016 12280
rect 38068 12271 38070 12280
rect 38016 12242 38068 12248
rect 38488 12102 38516 13466
rect 38660 13320 38712 13326
rect 38660 13262 38712 13268
rect 38568 13184 38620 13190
rect 38568 13126 38620 13132
rect 38580 12918 38608 13126
rect 38568 12912 38620 12918
rect 38568 12854 38620 12860
rect 38568 12232 38620 12238
rect 38568 12174 38620 12180
rect 38384 12096 38436 12102
rect 38384 12038 38436 12044
rect 38476 12096 38528 12102
rect 38476 12038 38528 12044
rect 38396 11218 38424 12038
rect 38384 11212 38436 11218
rect 38384 11154 38436 11160
rect 38476 10668 38528 10674
rect 38476 10610 38528 10616
rect 38488 10266 38516 10610
rect 38580 10470 38608 12174
rect 38672 10742 38700 13262
rect 38764 12442 38792 13874
rect 38844 12640 38896 12646
rect 38844 12582 38896 12588
rect 38752 12436 38804 12442
rect 38752 12378 38804 12384
rect 38750 12336 38806 12345
rect 38750 12271 38806 12280
rect 38764 12238 38792 12271
rect 38856 12238 38884 12582
rect 38752 12232 38804 12238
rect 38752 12174 38804 12180
rect 38844 12232 38896 12238
rect 38844 12174 38896 12180
rect 38948 11150 38976 14894
rect 39028 14612 39080 14618
rect 39028 14554 39080 14560
rect 39040 14278 39068 14554
rect 39028 14272 39080 14278
rect 39028 14214 39080 14220
rect 40328 13870 40356 14962
rect 41064 14958 41092 15030
rect 41052 14952 41104 14958
rect 41052 14894 41104 14900
rect 40408 14272 40460 14278
rect 40408 14214 40460 14220
rect 40420 13938 40448 14214
rect 40408 13932 40460 13938
rect 40408 13874 40460 13880
rect 40316 13864 40368 13870
rect 40316 13806 40368 13812
rect 40420 13326 40448 13874
rect 40776 13864 40828 13870
rect 40776 13806 40828 13812
rect 39028 13320 39080 13326
rect 39028 13262 39080 13268
rect 40408 13320 40460 13326
rect 40408 13262 40460 13268
rect 39040 12918 39068 13262
rect 39120 13184 39172 13190
rect 39120 13126 39172 13132
rect 39028 12912 39080 12918
rect 39028 12854 39080 12860
rect 39132 12646 39160 13126
rect 40788 12850 40816 13806
rect 41064 13258 41092 14894
rect 41524 14414 41552 15098
rect 41604 15020 41656 15026
rect 41604 14962 41656 14968
rect 41616 14482 41644 14962
rect 41696 14544 41748 14550
rect 41696 14486 41748 14492
rect 41604 14476 41656 14482
rect 41604 14418 41656 14424
rect 41512 14408 41564 14414
rect 41512 14350 41564 14356
rect 41420 14068 41472 14074
rect 41420 14010 41472 14016
rect 41432 13530 41460 14010
rect 41708 13938 41736 14486
rect 42260 14414 42288 15370
rect 42248 14408 42300 14414
rect 42248 14350 42300 14356
rect 41880 14272 41932 14278
rect 41880 14214 41932 14220
rect 41892 14074 41920 14214
rect 41880 14068 41932 14074
rect 41880 14010 41932 14016
rect 41696 13932 41748 13938
rect 41696 13874 41748 13880
rect 41420 13524 41472 13530
rect 41420 13466 41472 13472
rect 41052 13252 41104 13258
rect 41052 13194 41104 13200
rect 41064 12918 41092 13194
rect 42260 13190 42288 14350
rect 42248 13184 42300 13190
rect 42248 13126 42300 13132
rect 41052 12912 41104 12918
rect 41052 12854 41104 12860
rect 40776 12844 40828 12850
rect 40776 12786 40828 12792
rect 39120 12640 39172 12646
rect 39120 12582 39172 12588
rect 39132 12238 39160 12582
rect 39948 12436 40000 12442
rect 40788 12434 40816 12786
rect 41052 12776 41104 12782
rect 41052 12718 41104 12724
rect 40788 12406 40908 12434
rect 39948 12378 40000 12384
rect 39120 12232 39172 12238
rect 39120 12174 39172 12180
rect 38936 11144 38988 11150
rect 38936 11086 38988 11092
rect 38660 10736 38712 10742
rect 38660 10678 38712 10684
rect 39132 10674 39160 12174
rect 39960 11286 39988 12378
rect 40776 12232 40828 12238
rect 40776 12174 40828 12180
rect 40316 11552 40368 11558
rect 40316 11494 40368 11500
rect 39948 11280 40000 11286
rect 39948 11222 40000 11228
rect 40328 10810 40356 11494
rect 40592 11280 40644 11286
rect 40592 11222 40644 11228
rect 40316 10804 40368 10810
rect 40316 10746 40368 10752
rect 39120 10668 39172 10674
rect 39120 10610 39172 10616
rect 39580 10668 39632 10674
rect 39580 10610 39632 10616
rect 38568 10464 38620 10470
rect 38568 10406 38620 10412
rect 38844 10464 38896 10470
rect 38844 10406 38896 10412
rect 38016 10260 38068 10266
rect 38016 10202 38068 10208
rect 38476 10260 38528 10266
rect 38476 10202 38528 10208
rect 37924 9988 37976 9994
rect 37924 9930 37976 9936
rect 37648 9648 37700 9654
rect 37648 9590 37700 9596
rect 37556 9172 37608 9178
rect 37556 9114 37608 9120
rect 37568 9081 37596 9114
rect 37554 9072 37610 9081
rect 37464 9036 37516 9042
rect 37554 9007 37610 9016
rect 37464 8978 37516 8984
rect 37660 8974 37688 9590
rect 37188 8968 37240 8974
rect 37188 8910 37240 8916
rect 37648 8968 37700 8974
rect 37648 8910 37700 8916
rect 37740 8968 37792 8974
rect 37740 8910 37792 8916
rect 37094 8528 37150 8537
rect 37094 8463 37150 8472
rect 37004 8424 37056 8430
rect 37200 8378 37228 8910
rect 37004 8366 37056 8372
rect 37016 8294 37044 8366
rect 37108 8350 37228 8378
rect 37004 8288 37056 8294
rect 37004 8230 37056 8236
rect 37108 7698 37136 8350
rect 37188 8288 37240 8294
rect 37188 8230 37240 8236
rect 37200 7750 37228 8230
rect 37752 7954 37780 8910
rect 37922 8392 37978 8401
rect 37922 8327 37924 8336
rect 37976 8327 37978 8336
rect 37924 8298 37976 8304
rect 37740 7948 37792 7954
rect 37740 7890 37792 7896
rect 38028 7886 38056 10202
rect 38856 10062 38884 10406
rect 39132 10266 39160 10610
rect 39592 10470 39620 10610
rect 40604 10470 40632 11222
rect 40788 11082 40816 12174
rect 40880 11150 40908 12406
rect 41064 11558 41092 12718
rect 42352 12374 42380 15524
rect 42524 15506 42576 15512
rect 42812 15094 42840 17750
rect 42984 17264 43036 17270
rect 42984 17206 43036 17212
rect 42892 16720 42944 16726
rect 42892 16662 42944 16668
rect 42904 16522 42932 16662
rect 42892 16516 42944 16522
rect 42892 16458 42944 16464
rect 42892 15360 42944 15366
rect 42892 15302 42944 15308
rect 42904 15162 42932 15302
rect 42892 15156 42944 15162
rect 42892 15098 42944 15104
rect 42800 15088 42852 15094
rect 42800 15030 42852 15036
rect 42524 14952 42576 14958
rect 42524 14894 42576 14900
rect 42536 13870 42564 14894
rect 42800 14340 42852 14346
rect 42800 14282 42852 14288
rect 42524 13864 42576 13870
rect 42524 13806 42576 13812
rect 42432 13320 42484 13326
rect 42432 13262 42484 13268
rect 42444 12918 42472 13262
rect 42432 12912 42484 12918
rect 42432 12854 42484 12860
rect 42536 12442 42564 13806
rect 42812 13734 42840 14282
rect 42800 13728 42852 13734
rect 42800 13670 42852 13676
rect 42812 13530 42840 13670
rect 42800 13524 42852 13530
rect 42800 13466 42852 13472
rect 42892 13320 42944 13326
rect 42892 13262 42944 13268
rect 42616 12844 42668 12850
rect 42616 12786 42668 12792
rect 42524 12436 42576 12442
rect 42524 12378 42576 12384
rect 42340 12368 42392 12374
rect 42340 12310 42392 12316
rect 42524 12232 42576 12238
rect 42524 12174 42576 12180
rect 41696 12164 41748 12170
rect 41696 12106 41748 12112
rect 41880 12164 41932 12170
rect 41880 12106 41932 12112
rect 41708 11898 41736 12106
rect 41696 11892 41748 11898
rect 41696 11834 41748 11840
rect 41892 11830 41920 12106
rect 42536 11937 42564 12174
rect 42522 11928 42578 11937
rect 42522 11863 42578 11872
rect 41880 11824 41932 11830
rect 41880 11766 41932 11772
rect 42536 11626 42564 11863
rect 42628 11762 42656 12786
rect 42904 12782 42932 13262
rect 42892 12776 42944 12782
rect 42892 12718 42944 12724
rect 42708 12096 42760 12102
rect 42708 12038 42760 12044
rect 42616 11756 42668 11762
rect 42616 11698 42668 11704
rect 42524 11620 42576 11626
rect 42524 11562 42576 11568
rect 41052 11552 41104 11558
rect 41052 11494 41104 11500
rect 41064 11150 41092 11494
rect 42720 11150 42748 12038
rect 42904 11830 42932 12718
rect 42892 11824 42944 11830
rect 42892 11766 42944 11772
rect 40868 11144 40920 11150
rect 40868 11086 40920 11092
rect 41052 11144 41104 11150
rect 41052 11086 41104 11092
rect 42708 11144 42760 11150
rect 42708 11086 42760 11092
rect 40776 11076 40828 11082
rect 40776 11018 40828 11024
rect 40788 10538 40816 11018
rect 40880 10810 40908 11086
rect 40868 10804 40920 10810
rect 40868 10746 40920 10752
rect 40776 10532 40828 10538
rect 40776 10474 40828 10480
rect 39580 10464 39632 10470
rect 39580 10406 39632 10412
rect 40592 10464 40644 10470
rect 40592 10406 40644 10412
rect 39120 10260 39172 10266
rect 39120 10202 39172 10208
rect 38844 10056 38896 10062
rect 38844 9998 38896 10004
rect 38936 9920 38988 9926
rect 38936 9862 38988 9868
rect 38948 9586 38976 9862
rect 39592 9586 39620 10406
rect 40788 10266 40816 10474
rect 41328 10464 41380 10470
rect 41328 10406 41380 10412
rect 40776 10260 40828 10266
rect 40776 10202 40828 10208
rect 41340 10062 41368 10406
rect 42248 10192 42300 10198
rect 42248 10134 42300 10140
rect 41236 10056 41288 10062
rect 41236 9998 41288 10004
rect 41328 10056 41380 10062
rect 41328 9998 41380 10004
rect 38936 9580 38988 9586
rect 38936 9522 38988 9528
rect 39580 9580 39632 9586
rect 39580 9522 39632 9528
rect 39764 9580 39816 9586
rect 39764 9522 39816 9528
rect 39776 9450 39804 9522
rect 39764 9444 39816 9450
rect 39764 9386 39816 9392
rect 39856 9444 39908 9450
rect 39856 9386 39908 9392
rect 38476 9376 38528 9382
rect 38476 9318 38528 9324
rect 38384 8016 38436 8022
rect 38106 7984 38162 7993
rect 38384 7958 38436 7964
rect 38106 7919 38162 7928
rect 38016 7880 38068 7886
rect 38016 7822 38068 7828
rect 38120 7818 38148 7919
rect 38108 7812 38160 7818
rect 38108 7754 38160 7760
rect 37016 7670 37136 7698
rect 37188 7744 37240 7750
rect 37188 7686 37240 7692
rect 37280 7744 37332 7750
rect 37280 7686 37332 7692
rect 36912 7472 36964 7478
rect 36912 7414 36964 7420
rect 36924 6798 36952 7414
rect 36912 6792 36964 6798
rect 36912 6734 36964 6740
rect 36820 6724 36872 6730
rect 36820 6666 36872 6672
rect 36832 6458 36860 6666
rect 36820 6452 36872 6458
rect 36820 6394 36872 6400
rect 37016 6202 37044 7670
rect 37096 7540 37148 7546
rect 37096 7482 37148 7488
rect 37108 7274 37136 7482
rect 37096 7268 37148 7274
rect 37096 7210 37148 7216
rect 37200 6866 37228 7686
rect 37188 6860 37240 6866
rect 37188 6802 37240 6808
rect 36924 6174 37044 6202
rect 36728 4616 36780 4622
rect 36542 4584 36598 4593
rect 36452 4548 36504 4554
rect 36728 4558 36780 4564
rect 36542 4519 36598 4528
rect 36452 4490 36504 4496
rect 36268 4480 36320 4486
rect 36268 4422 36320 4428
rect 36556 4214 36584 4519
rect 36924 4321 36952 6174
rect 37004 6112 37056 6118
rect 37004 6054 37056 6060
rect 37016 4622 37044 6054
rect 37004 4616 37056 4622
rect 37004 4558 37056 4564
rect 36910 4312 36966 4321
rect 36910 4247 36966 4256
rect 36544 4208 36596 4214
rect 36544 4150 36596 4156
rect 36082 4111 36138 4120
rect 36176 4140 36228 4146
rect 36176 4082 36228 4088
rect 36360 3936 36412 3942
rect 36360 3878 36412 3884
rect 36372 3505 36400 3878
rect 36924 3602 36952 4247
rect 37292 4049 37320 7686
rect 38396 7410 38424 7958
rect 37464 7404 37516 7410
rect 37464 7346 37516 7352
rect 38384 7404 38436 7410
rect 38384 7346 38436 7352
rect 37476 7002 37504 7346
rect 37740 7336 37792 7342
rect 37740 7278 37792 7284
rect 37752 7002 37780 7278
rect 37464 6996 37516 7002
rect 37464 6938 37516 6944
rect 37740 6996 37792 7002
rect 37740 6938 37792 6944
rect 37372 6860 37424 6866
rect 37372 6802 37424 6808
rect 37464 6860 37516 6866
rect 37464 6802 37516 6808
rect 37384 6662 37412 6802
rect 37372 6656 37424 6662
rect 37372 6598 37424 6604
rect 37278 4040 37334 4049
rect 37384 4010 37412 6598
rect 37476 5778 37504 6802
rect 38292 6452 38344 6458
rect 38292 6394 38344 6400
rect 38304 5846 38332 6394
rect 38292 5840 38344 5846
rect 38292 5782 38344 5788
rect 37464 5772 37516 5778
rect 37464 5714 37516 5720
rect 38292 5296 38344 5302
rect 38292 5238 38344 5244
rect 37556 5160 37608 5166
rect 37556 5102 37608 5108
rect 37568 4622 37596 5102
rect 37556 4616 37608 4622
rect 37556 4558 37608 4564
rect 37568 4282 37596 4558
rect 38304 4486 38332 5238
rect 38488 4729 38516 9318
rect 39578 9208 39634 9217
rect 39578 9143 39634 9152
rect 39120 8968 39172 8974
rect 39120 8910 39172 8916
rect 38752 8832 38804 8838
rect 38752 8774 38804 8780
rect 38764 8498 38792 8774
rect 38752 8492 38804 8498
rect 38752 8434 38804 8440
rect 38568 8356 38620 8362
rect 38568 8298 38620 8304
rect 38580 7886 38608 8298
rect 38764 8022 38792 8434
rect 39132 8430 39160 8910
rect 39592 8634 39620 9143
rect 39580 8628 39632 8634
rect 39580 8570 39632 8576
rect 39776 8498 39804 9386
rect 39868 9178 39896 9386
rect 39856 9172 39908 9178
rect 39856 9114 39908 9120
rect 39764 8492 39816 8498
rect 39764 8434 39816 8440
rect 39120 8424 39172 8430
rect 39120 8366 39172 8372
rect 38752 8016 38804 8022
rect 38752 7958 38804 7964
rect 39132 7954 39160 8366
rect 41248 7954 41276 9998
rect 42260 9722 42288 10134
rect 42432 10124 42484 10130
rect 42432 10066 42484 10072
rect 42444 9722 42472 10066
rect 42248 9716 42300 9722
rect 42248 9658 42300 9664
rect 42432 9716 42484 9722
rect 42432 9658 42484 9664
rect 42800 9648 42852 9654
rect 42800 9590 42852 9596
rect 42616 9580 42668 9586
rect 42616 9522 42668 9528
rect 42708 9580 42760 9586
rect 42708 9522 42760 9528
rect 41696 9376 41748 9382
rect 41696 9318 41748 9324
rect 41512 9036 41564 9042
rect 41512 8978 41564 8984
rect 41524 8498 41552 8978
rect 41604 8628 41656 8634
rect 41604 8570 41656 8576
rect 41512 8492 41564 8498
rect 41512 8434 41564 8440
rect 41524 8378 41552 8434
rect 41432 8350 41552 8378
rect 39120 7948 39172 7954
rect 39120 7890 39172 7896
rect 40040 7948 40092 7954
rect 40040 7890 40092 7896
rect 41236 7948 41288 7954
rect 41236 7890 41288 7896
rect 38568 7880 38620 7886
rect 38568 7822 38620 7828
rect 39120 7200 39172 7206
rect 39120 7142 39172 7148
rect 39132 6662 39160 7142
rect 40052 7002 40080 7890
rect 40040 6996 40092 7002
rect 40040 6938 40092 6944
rect 39120 6656 39172 6662
rect 39120 6598 39172 6604
rect 40052 6474 40080 6938
rect 40684 6724 40736 6730
rect 40684 6666 40736 6672
rect 39868 6446 40080 6474
rect 39672 6180 39724 6186
rect 39672 6122 39724 6128
rect 39684 6089 39712 6122
rect 39670 6080 39726 6089
rect 39670 6015 39726 6024
rect 38752 5908 38804 5914
rect 38752 5850 38804 5856
rect 38568 5704 38620 5710
rect 38568 5646 38620 5652
rect 38580 5234 38608 5646
rect 38764 5370 38792 5850
rect 39868 5778 39896 6446
rect 40040 6316 40092 6322
rect 40040 6258 40092 6264
rect 39948 6112 40000 6118
rect 39948 6054 40000 6060
rect 39856 5772 39908 5778
rect 39856 5714 39908 5720
rect 39868 5574 39896 5714
rect 39960 5710 39988 6054
rect 39948 5704 40000 5710
rect 39948 5646 40000 5652
rect 39856 5568 39908 5574
rect 39856 5510 39908 5516
rect 38752 5364 38804 5370
rect 38752 5306 38804 5312
rect 38568 5228 38620 5234
rect 38568 5170 38620 5176
rect 38474 4720 38530 4729
rect 38474 4655 38530 4664
rect 38292 4480 38344 4486
rect 38290 4448 38292 4457
rect 38344 4448 38346 4457
rect 38290 4383 38346 4392
rect 38290 4312 38346 4321
rect 37556 4276 37608 4282
rect 38290 4247 38346 4256
rect 37556 4218 37608 4224
rect 37278 3975 37334 3984
rect 37372 4004 37424 4010
rect 36912 3596 36964 3602
rect 36912 3538 36964 3544
rect 37188 3528 37240 3534
rect 36358 3496 36414 3505
rect 37292 3516 37320 3975
rect 37372 3946 37424 3952
rect 37240 3488 37320 3516
rect 37188 3470 37240 3476
rect 36358 3431 36414 3440
rect 37384 3346 37412 3946
rect 37464 3732 37516 3738
rect 37464 3674 37516 3680
rect 37476 3534 37504 3674
rect 37556 3596 37608 3602
rect 37556 3538 37608 3544
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 37292 3318 37412 3346
rect 35808 3188 35860 3194
rect 35808 3130 35860 3136
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 35716 3052 35768 3058
rect 35716 2994 35768 3000
rect 35532 2984 35584 2990
rect 35530 2952 35532 2961
rect 35584 2952 35586 2961
rect 35530 2887 35586 2896
rect 35728 2854 35756 2994
rect 35716 2848 35768 2854
rect 35716 2790 35768 2796
rect 35820 2038 35848 3130
rect 37292 2990 37320 3318
rect 37280 2984 37332 2990
rect 37280 2926 37332 2932
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 36268 2372 36320 2378
rect 36268 2314 36320 2320
rect 35898 2136 35954 2145
rect 35898 2071 35954 2080
rect 35912 2038 35940 2071
rect 35808 2032 35860 2038
rect 35808 1974 35860 1980
rect 35900 2032 35952 2038
rect 35900 1974 35952 1980
rect 35268 870 35388 898
rect 35268 800 35296 870
rect 36280 800 36308 2314
rect 36740 800 36768 2790
rect 37568 2774 37596 3538
rect 38304 3534 38332 4247
rect 38488 4146 38516 4655
rect 38580 4622 38608 5170
rect 40052 4622 40080 6258
rect 40592 6248 40644 6254
rect 40592 6190 40644 6196
rect 40316 5568 40368 5574
rect 40316 5510 40368 5516
rect 40408 5568 40460 5574
rect 40408 5510 40460 5516
rect 40224 5296 40276 5302
rect 40224 5238 40276 5244
rect 40132 5228 40184 5234
rect 40132 5170 40184 5176
rect 40144 5030 40172 5170
rect 40132 5024 40184 5030
rect 40132 4966 40184 4972
rect 38568 4616 38620 4622
rect 38568 4558 38620 4564
rect 40040 4616 40092 4622
rect 40040 4558 40092 4564
rect 38476 4140 38528 4146
rect 38580 4128 38608 4558
rect 39028 4548 39080 4554
rect 39028 4490 39080 4496
rect 40132 4548 40184 4554
rect 40132 4490 40184 4496
rect 39040 4282 39068 4490
rect 39028 4276 39080 4282
rect 39028 4218 39080 4224
rect 39040 4146 39068 4218
rect 38660 4140 38712 4146
rect 38580 4100 38660 4128
rect 38476 4082 38528 4088
rect 38660 4082 38712 4088
rect 38844 4140 38896 4146
rect 38844 4082 38896 4088
rect 39028 4140 39080 4146
rect 39028 4082 39080 4088
rect 38382 3632 38438 3641
rect 38856 3602 38884 4082
rect 39120 3936 39172 3942
rect 39120 3878 39172 3884
rect 39856 3936 39908 3942
rect 39856 3878 39908 3884
rect 39132 3602 39160 3878
rect 38382 3567 38438 3576
rect 38844 3596 38896 3602
rect 38396 3534 38424 3567
rect 38844 3538 38896 3544
rect 39120 3596 39172 3602
rect 39120 3538 39172 3544
rect 37740 3528 37792 3534
rect 37740 3470 37792 3476
rect 38292 3528 38344 3534
rect 38292 3470 38344 3476
rect 38384 3528 38436 3534
rect 38384 3470 38436 3476
rect 37752 3194 37780 3470
rect 37832 3392 37884 3398
rect 37832 3334 37884 3340
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 37844 3126 37872 3334
rect 37832 3120 37884 3126
rect 37832 3062 37884 3068
rect 37384 2746 37596 2774
rect 37384 2446 37412 2746
rect 37372 2440 37424 2446
rect 37372 2382 37424 2388
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 37752 800 37780 2314
rect 38212 800 38240 3334
rect 38856 3194 38884 3538
rect 39672 3392 39724 3398
rect 39672 3334 39724 3340
rect 38844 3188 38896 3194
rect 38844 3130 38896 3136
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38672 2650 38700 2790
rect 38660 2644 38712 2650
rect 38660 2586 38712 2592
rect 39212 2372 39264 2378
rect 39212 2314 39264 2320
rect 39224 800 39252 2314
rect 39684 800 39712 3334
rect 39868 3126 39896 3878
rect 39948 3528 40000 3534
rect 40144 3516 40172 4490
rect 40236 4486 40264 5238
rect 40224 4480 40276 4486
rect 40224 4422 40276 4428
rect 40224 4140 40276 4146
rect 40224 4082 40276 4088
rect 40236 3738 40264 4082
rect 40224 3732 40276 3738
rect 40224 3674 40276 3680
rect 40000 3488 40172 3516
rect 39948 3470 40000 3476
rect 39856 3120 39908 3126
rect 39856 3062 39908 3068
rect 40328 3058 40356 5510
rect 40420 5234 40448 5510
rect 40604 5370 40632 6190
rect 40592 5364 40644 5370
rect 40592 5306 40644 5312
rect 40408 5228 40460 5234
rect 40408 5170 40460 5176
rect 40500 5228 40552 5234
rect 40500 5170 40552 5176
rect 40512 5098 40540 5170
rect 40500 5092 40552 5098
rect 40500 5034 40552 5040
rect 40592 4684 40644 4690
rect 40592 4626 40644 4632
rect 40604 4146 40632 4626
rect 40696 4554 40724 6666
rect 41432 6662 41460 8350
rect 41512 8288 41564 8294
rect 41512 8230 41564 8236
rect 41524 7886 41552 8230
rect 41512 7880 41564 7886
rect 41512 7822 41564 7828
rect 41420 6656 41472 6662
rect 41420 6598 41472 6604
rect 41432 6322 41460 6598
rect 41420 6316 41472 6322
rect 41420 6258 41472 6264
rect 41328 5772 41380 5778
rect 41328 5714 41380 5720
rect 41340 5574 41368 5714
rect 41328 5568 41380 5574
rect 41328 5510 41380 5516
rect 40960 5364 41012 5370
rect 40960 5306 41012 5312
rect 40684 4548 40736 4554
rect 40684 4490 40736 4496
rect 40972 4282 41000 5306
rect 40960 4276 41012 4282
rect 40960 4218 41012 4224
rect 41052 4276 41104 4282
rect 41052 4218 41104 4224
rect 41064 4146 41092 4218
rect 41340 4146 41368 5510
rect 41616 5030 41644 8570
rect 41708 8362 41736 9318
rect 41788 9172 41840 9178
rect 41788 9114 41840 9120
rect 42248 9172 42300 9178
rect 42248 9114 42300 9120
rect 41800 8634 41828 9114
rect 42260 8906 42288 9114
rect 42432 8968 42484 8974
rect 42432 8910 42484 8916
rect 41880 8900 41932 8906
rect 41880 8842 41932 8848
rect 42248 8900 42300 8906
rect 42248 8842 42300 8848
rect 41892 8634 41920 8842
rect 42340 8832 42392 8838
rect 42340 8774 42392 8780
rect 41788 8628 41840 8634
rect 41788 8570 41840 8576
rect 41880 8628 41932 8634
rect 41880 8570 41932 8576
rect 42352 8498 42380 8774
rect 42340 8492 42392 8498
rect 42340 8434 42392 8440
rect 41696 8356 41748 8362
rect 41696 8298 41748 8304
rect 42444 8022 42472 8910
rect 42628 8498 42656 9522
rect 42720 9217 42748 9522
rect 42812 9518 42840 9590
rect 42892 9580 42944 9586
rect 42892 9522 42944 9528
rect 42800 9512 42852 9518
rect 42800 9454 42852 9460
rect 42706 9208 42762 9217
rect 42706 9143 42762 9152
rect 42904 8566 42932 9522
rect 42892 8560 42944 8566
rect 42892 8502 42944 8508
rect 42616 8492 42668 8498
rect 42616 8434 42668 8440
rect 42708 8492 42760 8498
rect 42708 8434 42760 8440
rect 42432 8016 42484 8022
rect 42432 7958 42484 7964
rect 42340 7880 42392 7886
rect 42340 7822 42392 7828
rect 42352 7546 42380 7822
rect 42340 7540 42392 7546
rect 42340 7482 42392 7488
rect 41972 7472 42024 7478
rect 41972 7414 42024 7420
rect 41880 6180 41932 6186
rect 41880 6122 41932 6128
rect 41892 5710 41920 6122
rect 41984 5710 42012 7414
rect 42444 7342 42472 7958
rect 42524 7744 42576 7750
rect 42524 7686 42576 7692
rect 42536 7478 42564 7686
rect 42524 7472 42576 7478
rect 42524 7414 42576 7420
rect 42720 7410 42748 8434
rect 42904 7954 42932 8502
rect 42892 7948 42944 7954
rect 42892 7890 42944 7896
rect 42904 7410 42932 7890
rect 42616 7404 42668 7410
rect 42616 7346 42668 7352
rect 42708 7404 42760 7410
rect 42708 7346 42760 7352
rect 42892 7404 42944 7410
rect 42892 7346 42944 7352
rect 42432 7336 42484 7342
rect 42432 7278 42484 7284
rect 41880 5704 41932 5710
rect 41880 5646 41932 5652
rect 41972 5704 42024 5710
rect 41972 5646 42024 5652
rect 41984 5574 42012 5646
rect 41696 5568 41748 5574
rect 41696 5510 41748 5516
rect 41972 5568 42024 5574
rect 41972 5510 42024 5516
rect 41420 5024 41472 5030
rect 41420 4966 41472 4972
rect 41604 5024 41656 5030
rect 41604 4966 41656 4972
rect 40592 4140 40644 4146
rect 40592 4082 40644 4088
rect 41052 4140 41104 4146
rect 41052 4082 41104 4088
rect 41328 4140 41380 4146
rect 41328 4082 41380 4088
rect 41144 3936 41196 3942
rect 41144 3878 41196 3884
rect 40316 3052 40368 3058
rect 40316 2994 40368 3000
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40500 2304 40552 2310
rect 40500 2246 40552 2252
rect 40512 1426 40540 2246
rect 40500 1420 40552 1426
rect 40500 1362 40552 1368
rect 40604 800 40632 2314
rect 40684 2032 40736 2038
rect 40684 1974 40736 1980
rect 40696 1494 40724 1974
rect 40684 1488 40736 1494
rect 40684 1430 40736 1436
rect 41156 800 41184 3878
rect 41432 3534 41460 4966
rect 41616 4826 41644 4966
rect 41708 4826 41736 5510
rect 41604 4820 41656 4826
rect 41604 4762 41656 4768
rect 41696 4820 41748 4826
rect 41696 4762 41748 4768
rect 42248 4480 42300 4486
rect 42248 4422 42300 4428
rect 42260 3534 42288 4422
rect 41420 3528 41472 3534
rect 41420 3470 41472 3476
rect 42156 3528 42208 3534
rect 42156 3470 42208 3476
rect 42248 3528 42300 3534
rect 42248 3470 42300 3476
rect 41432 3126 41460 3470
rect 41420 3120 41472 3126
rect 41420 3062 41472 3068
rect 42168 3058 42196 3470
rect 42156 3052 42208 3058
rect 42156 2994 42208 3000
rect 42444 2446 42472 7278
rect 42628 6186 42656 7346
rect 42616 6180 42668 6186
rect 42616 6122 42668 6128
rect 42522 6080 42578 6089
rect 42522 6015 42578 6024
rect 42536 5846 42564 6015
rect 42524 5840 42576 5846
rect 42524 5782 42576 5788
rect 42720 5642 42748 7346
rect 42892 6180 42944 6186
rect 42892 6122 42944 6128
rect 42904 5710 42932 6122
rect 42892 5704 42944 5710
rect 42892 5646 42944 5652
rect 42708 5636 42760 5642
rect 42708 5578 42760 5584
rect 42996 5574 43024 17206
rect 43088 14958 43116 17818
rect 43180 17678 43208 18362
rect 43904 18080 43956 18086
rect 43904 18022 43956 18028
rect 43916 17882 43944 18022
rect 43904 17876 43956 17882
rect 43904 17818 43956 17824
rect 44376 17678 44404 18566
rect 47320 18358 47348 18566
rect 47308 18352 47360 18358
rect 47308 18294 47360 18300
rect 46664 18284 46716 18290
rect 46664 18226 46716 18232
rect 44456 17740 44508 17746
rect 44456 17682 44508 17688
rect 43168 17672 43220 17678
rect 43168 17614 43220 17620
rect 44088 17672 44140 17678
rect 44088 17614 44140 17620
rect 44364 17672 44416 17678
rect 44364 17614 44416 17620
rect 43180 17338 43208 17614
rect 43168 17332 43220 17338
rect 43168 17274 43220 17280
rect 44100 17270 44128 17614
rect 44088 17264 44140 17270
rect 44088 17206 44140 17212
rect 44100 16794 44128 17206
rect 44376 17202 44404 17614
rect 44468 17270 44496 17682
rect 46676 17678 46704 18226
rect 47032 18080 47084 18086
rect 47032 18022 47084 18028
rect 47044 17882 47072 18022
rect 47504 17882 47532 18702
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 55416 18426 55444 39374
rect 55404 18420 55456 18426
rect 55404 18362 55456 18368
rect 47584 18284 47636 18290
rect 47584 18226 47636 18232
rect 53564 18284 53616 18290
rect 53564 18226 53616 18232
rect 47032 17876 47084 17882
rect 47032 17818 47084 17824
rect 47492 17876 47544 17882
rect 47492 17818 47544 17824
rect 46664 17672 46716 17678
rect 46664 17614 46716 17620
rect 44456 17264 44508 17270
rect 44456 17206 44508 17212
rect 45284 17264 45336 17270
rect 45284 17206 45336 17212
rect 44364 17196 44416 17202
rect 44364 17138 44416 17144
rect 44088 16788 44140 16794
rect 44088 16730 44140 16736
rect 44376 16590 44404 17138
rect 45296 16590 45324 17206
rect 46676 16794 46704 17614
rect 46940 17604 46992 17610
rect 46940 17546 46992 17552
rect 46952 16794 46980 17546
rect 46664 16788 46716 16794
rect 46664 16730 46716 16736
rect 46940 16788 46992 16794
rect 46940 16730 46992 16736
rect 47596 16658 47624 18226
rect 53380 18216 53432 18222
rect 53380 18158 53432 18164
rect 47860 18080 47912 18086
rect 47860 18022 47912 18028
rect 47872 17678 47900 18022
rect 47860 17672 47912 17678
rect 47860 17614 47912 17620
rect 47872 17270 47900 17614
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 47860 17264 47912 17270
rect 47860 17206 47912 17212
rect 51448 17196 51500 17202
rect 51448 17138 51500 17144
rect 51080 16992 51132 16998
rect 51080 16934 51132 16940
rect 47584 16652 47636 16658
rect 47584 16594 47636 16600
rect 50804 16652 50856 16658
rect 50804 16594 50856 16600
rect 44364 16584 44416 16590
rect 44364 16526 44416 16532
rect 45284 16584 45336 16590
rect 45284 16526 45336 16532
rect 45836 16584 45888 16590
rect 45836 16526 45888 16532
rect 45928 16584 45980 16590
rect 45928 16526 45980 16532
rect 45008 16516 45060 16522
rect 45008 16458 45060 16464
rect 45020 16114 45048 16458
rect 45848 16182 45876 16526
rect 45836 16176 45888 16182
rect 45836 16118 45888 16124
rect 45940 16114 45968 16526
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 46756 16448 46808 16454
rect 46756 16390 46808 16396
rect 46768 16250 46796 16390
rect 47688 16250 47716 16458
rect 47860 16448 47912 16454
rect 47860 16390 47912 16396
rect 49240 16448 49292 16454
rect 49240 16390 49292 16396
rect 46756 16244 46808 16250
rect 46756 16186 46808 16192
rect 47676 16244 47728 16250
rect 47676 16186 47728 16192
rect 47872 16114 47900 16390
rect 49252 16182 49280 16390
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 49240 16176 49292 16182
rect 49240 16118 49292 16124
rect 43628 16108 43680 16114
rect 43628 16050 43680 16056
rect 45008 16108 45060 16114
rect 45008 16050 45060 16056
rect 45928 16108 45980 16114
rect 45928 16050 45980 16056
rect 47860 16108 47912 16114
rect 47860 16050 47912 16056
rect 43640 15570 43668 16050
rect 43720 15904 43772 15910
rect 43720 15846 43772 15852
rect 43628 15564 43680 15570
rect 43628 15506 43680 15512
rect 43732 15502 43760 15846
rect 43536 15496 43588 15502
rect 43536 15438 43588 15444
rect 43720 15496 43772 15502
rect 43720 15438 43772 15444
rect 43168 15088 43220 15094
rect 43168 15030 43220 15036
rect 43076 14952 43128 14958
rect 43076 14894 43128 14900
rect 43076 12436 43128 12442
rect 43180 12434 43208 15030
rect 43548 12782 43576 15438
rect 44088 15428 44140 15434
rect 44088 15370 44140 15376
rect 44100 15094 44128 15370
rect 45020 15162 45048 16050
rect 45940 15706 45968 16050
rect 45928 15700 45980 15706
rect 45928 15642 45980 15648
rect 48044 15496 48096 15502
rect 48044 15438 48096 15444
rect 47860 15360 47912 15366
rect 47860 15302 47912 15308
rect 45008 15156 45060 15162
rect 45008 15098 45060 15104
rect 47872 15094 47900 15302
rect 44088 15088 44140 15094
rect 44088 15030 44140 15036
rect 47860 15088 47912 15094
rect 47860 15030 47912 15036
rect 46020 14952 46072 14958
rect 46020 14894 46072 14900
rect 46032 13394 46060 14894
rect 48056 14618 48084 15438
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 49056 14884 49108 14890
rect 49056 14826 49108 14832
rect 48964 14816 49016 14822
rect 48964 14758 49016 14764
rect 48044 14612 48096 14618
rect 48044 14554 48096 14560
rect 48976 14346 49004 14758
rect 49068 14414 49096 14826
rect 50620 14816 50672 14822
rect 50620 14758 50672 14764
rect 49056 14408 49108 14414
rect 49056 14350 49108 14356
rect 48504 14340 48556 14346
rect 48504 14282 48556 14288
rect 48964 14340 49016 14346
rect 48964 14282 49016 14288
rect 47860 14272 47912 14278
rect 47860 14214 47912 14220
rect 47400 13932 47452 13938
rect 47400 13874 47452 13880
rect 46204 13728 46256 13734
rect 46204 13670 46256 13676
rect 46020 13388 46072 13394
rect 46020 13330 46072 13336
rect 44456 12844 44508 12850
rect 44456 12786 44508 12792
rect 43536 12776 43588 12782
rect 43536 12718 43588 12724
rect 43720 12776 43772 12782
rect 43720 12718 43772 12724
rect 43548 12646 43576 12718
rect 43536 12640 43588 12646
rect 43536 12582 43588 12588
rect 43628 12640 43680 12646
rect 43628 12582 43680 12588
rect 43180 12406 43300 12434
rect 43076 12378 43128 12384
rect 43088 11830 43116 12378
rect 43272 12374 43300 12406
rect 43260 12368 43312 12374
rect 43260 12310 43312 12316
rect 43260 12232 43312 12238
rect 43180 12192 43260 12220
rect 43076 11824 43128 11830
rect 43076 11766 43128 11772
rect 43076 11348 43128 11354
rect 43076 11290 43128 11296
rect 43088 11150 43116 11290
rect 43076 11144 43128 11150
rect 43076 11086 43128 11092
rect 43180 11082 43208 12192
rect 43260 12174 43312 12180
rect 43260 11756 43312 11762
rect 43260 11698 43312 11704
rect 43272 11354 43300 11698
rect 43260 11348 43312 11354
rect 43260 11290 43312 11296
rect 43640 11218 43668 12582
rect 43732 12442 43760 12718
rect 43996 12708 44048 12714
rect 43996 12650 44048 12656
rect 43720 12436 43772 12442
rect 43720 12378 43772 12384
rect 43628 11212 43680 11218
rect 43628 11154 43680 11160
rect 43732 11150 43760 12378
rect 44008 12238 44036 12650
rect 43996 12232 44048 12238
rect 43996 12174 44048 12180
rect 43996 12096 44048 12102
rect 43996 12038 44048 12044
rect 44008 11830 44036 12038
rect 43996 11824 44048 11830
rect 43996 11766 44048 11772
rect 44468 11354 44496 12786
rect 46032 11762 46060 13330
rect 46112 13252 46164 13258
rect 46112 13194 46164 13200
rect 46124 12986 46152 13194
rect 46112 12980 46164 12986
rect 46112 12922 46164 12928
rect 46216 12850 46244 13670
rect 47412 13190 47440 13874
rect 47872 13870 47900 14214
rect 47860 13864 47912 13870
rect 47860 13806 47912 13812
rect 48516 13326 48544 14282
rect 48504 13320 48556 13326
rect 48504 13262 48556 13268
rect 48688 13252 48740 13258
rect 48688 13194 48740 13200
rect 47400 13184 47452 13190
rect 47400 13126 47452 13132
rect 48596 13184 48648 13190
rect 48596 13126 48648 13132
rect 46204 12844 46256 12850
rect 46204 12786 46256 12792
rect 47412 12306 47440 13126
rect 48044 12912 48096 12918
rect 48044 12854 48096 12860
rect 47400 12300 47452 12306
rect 47400 12242 47452 12248
rect 47676 12232 47728 12238
rect 47676 12174 47728 12180
rect 46570 11928 46626 11937
rect 46570 11863 46572 11872
rect 46624 11863 46626 11872
rect 46572 11834 46624 11840
rect 46584 11762 46612 11834
rect 46020 11756 46072 11762
rect 46020 11698 46072 11704
rect 46572 11756 46624 11762
rect 46572 11698 46624 11704
rect 44456 11348 44508 11354
rect 44456 11290 44508 11296
rect 47688 11150 47716 12174
rect 47860 12096 47912 12102
rect 47860 12038 47912 12044
rect 43720 11144 43772 11150
rect 43720 11086 43772 11092
rect 47676 11144 47728 11150
rect 47676 11086 47728 11092
rect 43168 11076 43220 11082
rect 43168 11018 43220 11024
rect 47584 10668 47636 10674
rect 47584 10610 47636 10616
rect 47124 10600 47176 10606
rect 47124 10542 47176 10548
rect 46572 10056 46624 10062
rect 46572 9998 46624 10004
rect 44640 9988 44692 9994
rect 44640 9930 44692 9936
rect 46480 9988 46532 9994
rect 46480 9930 46532 9936
rect 43168 9444 43220 9450
rect 43168 9386 43220 9392
rect 43180 8974 43208 9386
rect 44548 9104 44600 9110
rect 44548 9046 44600 9052
rect 43168 8968 43220 8974
rect 43168 8910 43220 8916
rect 44180 8900 44232 8906
rect 44180 8842 44232 8848
rect 44192 7886 44220 8842
rect 44560 8430 44588 9046
rect 44548 8424 44600 8430
rect 44548 8366 44600 8372
rect 44180 7880 44232 7886
rect 44180 7822 44232 7828
rect 44272 7880 44324 7886
rect 44272 7822 44324 7828
rect 44284 7698 44312 7822
rect 44192 7670 44312 7698
rect 43076 7200 43128 7206
rect 43076 7142 43128 7148
rect 43088 6322 43116 7142
rect 44192 6866 44220 7670
rect 44652 7410 44680 9930
rect 45928 9920 45980 9926
rect 45928 9862 45980 9868
rect 45940 9654 45968 9862
rect 45928 9648 45980 9654
rect 45928 9590 45980 9596
rect 45376 9444 45428 9450
rect 45376 9386 45428 9392
rect 45006 9208 45062 9217
rect 45006 9143 45062 9152
rect 44732 9104 44784 9110
rect 44732 9046 44784 9052
rect 44744 8566 44772 9046
rect 45020 9042 45048 9143
rect 45388 9042 45416 9386
rect 46296 9376 46348 9382
rect 46296 9318 46348 9324
rect 46308 9178 46336 9318
rect 46204 9172 46256 9178
rect 46204 9114 46256 9120
rect 46296 9172 46348 9178
rect 46296 9114 46348 9120
rect 46216 9058 46244 9114
rect 45008 9036 45060 9042
rect 45008 8978 45060 8984
rect 45376 9036 45428 9042
rect 46216 9030 46336 9058
rect 45376 8978 45428 8984
rect 44916 8968 44968 8974
rect 44916 8910 44968 8916
rect 44732 8560 44784 8566
rect 44732 8502 44784 8508
rect 44928 8498 44956 8910
rect 45020 8566 45048 8978
rect 46308 8906 46336 9030
rect 45468 8900 45520 8906
rect 45468 8842 45520 8848
rect 46296 8900 46348 8906
rect 46296 8842 46348 8848
rect 45480 8634 45508 8842
rect 46204 8832 46256 8838
rect 46204 8774 46256 8780
rect 45468 8628 45520 8634
rect 45468 8570 45520 8576
rect 45008 8560 45060 8566
rect 45008 8502 45060 8508
rect 44916 8492 44968 8498
rect 44916 8434 44968 8440
rect 45480 7954 45508 8570
rect 46216 8566 46244 8774
rect 46204 8560 46256 8566
rect 46204 8502 46256 8508
rect 46492 8090 46520 9930
rect 46584 8838 46612 9998
rect 47136 9586 47164 10542
rect 47596 10266 47624 10610
rect 47872 10266 47900 12038
rect 47584 10260 47636 10266
rect 47584 10202 47636 10208
rect 47860 10260 47912 10266
rect 47860 10202 47912 10208
rect 48056 10130 48084 12854
rect 48608 12442 48636 13126
rect 48700 12850 48728 13194
rect 49068 12986 49096 14350
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 50632 13530 50660 14758
rect 50816 14482 50844 16594
rect 51092 16590 51120 16934
rect 51080 16584 51132 16590
rect 51080 16526 51132 16532
rect 51460 16250 51488 17138
rect 53392 16794 53420 18158
rect 53380 16788 53432 16794
rect 53380 16730 53432 16736
rect 53196 16516 53248 16522
rect 53196 16458 53248 16464
rect 52460 16448 52512 16454
rect 52460 16390 52512 16396
rect 51448 16244 51500 16250
rect 51448 16186 51500 16192
rect 51080 16176 51132 16182
rect 51080 16118 51132 16124
rect 50896 14816 50948 14822
rect 50896 14758 50948 14764
rect 50804 14476 50856 14482
rect 50804 14418 50856 14424
rect 50620 13524 50672 13530
rect 50620 13466 50672 13472
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 49056 12980 49108 12986
rect 49056 12922 49108 12928
rect 50816 12850 50844 14418
rect 50908 14414 50936 14758
rect 51092 14618 51120 16118
rect 51540 15904 51592 15910
rect 51540 15846 51592 15852
rect 51552 15706 51580 15846
rect 51540 15700 51592 15706
rect 51540 15642 51592 15648
rect 52472 15638 52500 16390
rect 52920 16176 52972 16182
rect 52920 16118 52972 16124
rect 52552 15904 52604 15910
rect 52552 15846 52604 15852
rect 52460 15632 52512 15638
rect 52460 15574 52512 15580
rect 52472 15502 52500 15574
rect 52564 15570 52592 15846
rect 52932 15706 52960 16118
rect 53208 15978 53236 16458
rect 53288 16108 53340 16114
rect 53288 16050 53340 16056
rect 53472 16108 53524 16114
rect 53472 16050 53524 16056
rect 53196 15972 53248 15978
rect 53196 15914 53248 15920
rect 52920 15700 52972 15706
rect 52920 15642 52972 15648
rect 53104 15632 53156 15638
rect 53104 15574 53156 15580
rect 52552 15564 52604 15570
rect 52552 15506 52604 15512
rect 52460 15496 52512 15502
rect 52460 15438 52512 15444
rect 52564 15026 52592 15506
rect 52552 15020 52604 15026
rect 52552 14962 52604 14968
rect 53116 14958 53144 15574
rect 53300 15502 53328 16050
rect 53484 15910 53512 16050
rect 53472 15904 53524 15910
rect 53472 15846 53524 15852
rect 53380 15632 53432 15638
rect 53380 15574 53432 15580
rect 53392 15502 53420 15574
rect 53288 15496 53340 15502
rect 53288 15438 53340 15444
rect 53380 15496 53432 15502
rect 53380 15438 53432 15444
rect 53300 15366 53328 15438
rect 53288 15360 53340 15366
rect 53288 15302 53340 15308
rect 53300 15026 53328 15302
rect 53576 15162 53604 18226
rect 53840 16448 53892 16454
rect 53840 16390 53892 16396
rect 53852 15502 53880 16390
rect 55588 16040 55640 16046
rect 55588 15982 55640 15988
rect 55404 15904 55456 15910
rect 55404 15846 55456 15852
rect 54024 15564 54076 15570
rect 54024 15506 54076 15512
rect 53840 15496 53892 15502
rect 53840 15438 53892 15444
rect 53564 15156 53616 15162
rect 53564 15098 53616 15104
rect 53288 15020 53340 15026
rect 53288 14962 53340 14968
rect 53104 14952 53156 14958
rect 53104 14894 53156 14900
rect 53196 14952 53248 14958
rect 53196 14894 53248 14900
rect 51080 14612 51132 14618
rect 51080 14554 51132 14560
rect 50896 14408 50948 14414
rect 50896 14350 50948 14356
rect 51908 14272 51960 14278
rect 51908 14214 51960 14220
rect 51264 13320 51316 13326
rect 51264 13262 51316 13268
rect 51172 13184 51224 13190
rect 51172 13126 51224 13132
rect 48688 12844 48740 12850
rect 48688 12786 48740 12792
rect 48872 12844 48924 12850
rect 48872 12786 48924 12792
rect 50804 12844 50856 12850
rect 50804 12786 50856 12792
rect 48596 12436 48648 12442
rect 48596 12378 48648 12384
rect 48700 12374 48728 12786
rect 48688 12368 48740 12374
rect 48688 12310 48740 12316
rect 48320 12232 48372 12238
rect 48320 12174 48372 12180
rect 48688 12232 48740 12238
rect 48688 12174 48740 12180
rect 48780 12232 48832 12238
rect 48780 12174 48832 12180
rect 48332 10810 48360 12174
rect 48700 11898 48728 12174
rect 48412 11892 48464 11898
rect 48412 11834 48464 11840
rect 48688 11892 48740 11898
rect 48688 11834 48740 11840
rect 48424 11150 48452 11834
rect 48792 11762 48820 12174
rect 48780 11756 48832 11762
rect 48780 11698 48832 11704
rect 48596 11688 48648 11694
rect 48596 11630 48648 11636
rect 48608 11286 48636 11630
rect 48884 11558 48912 12786
rect 50816 12458 50844 12786
rect 51080 12640 51132 12646
rect 51080 12582 51132 12588
rect 51092 12458 51120 12582
rect 50816 12430 51120 12458
rect 51184 12442 51212 13126
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 48688 11552 48740 11558
rect 48688 11494 48740 11500
rect 48872 11552 48924 11558
rect 48872 11494 48924 11500
rect 48596 11280 48648 11286
rect 48596 11222 48648 11228
rect 48412 11144 48464 11150
rect 48412 11086 48464 11092
rect 48320 10804 48372 10810
rect 48320 10746 48372 10752
rect 48700 10198 48728 11494
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 48688 10192 48740 10198
rect 48688 10134 48740 10140
rect 51092 10130 51120 12430
rect 51172 12436 51224 12442
rect 51172 12378 51224 12384
rect 51276 12374 51304 13262
rect 51816 13184 51868 13190
rect 51816 13126 51868 13132
rect 51828 12918 51856 13126
rect 51816 12912 51868 12918
rect 51816 12854 51868 12860
rect 51920 12442 51948 14214
rect 52184 14068 52236 14074
rect 52184 14010 52236 14016
rect 52000 13184 52052 13190
rect 52000 13126 52052 13132
rect 51448 12436 51500 12442
rect 51448 12378 51500 12384
rect 51908 12436 51960 12442
rect 51908 12378 51960 12384
rect 51264 12368 51316 12374
rect 51264 12310 51316 12316
rect 51460 12306 51488 12378
rect 52012 12374 52040 13126
rect 52196 12986 52224 14010
rect 53116 13870 53144 14894
rect 53208 14618 53236 14894
rect 53196 14612 53248 14618
rect 53196 14554 53248 14560
rect 53208 14006 53236 14554
rect 53852 14006 53880 15438
rect 54036 14958 54064 15506
rect 55416 15434 55444 15846
rect 55220 15428 55272 15434
rect 55220 15370 55272 15376
rect 55404 15428 55456 15434
rect 55404 15370 55456 15376
rect 55036 15156 55088 15162
rect 55036 15098 55088 15104
rect 55048 14958 55076 15098
rect 55232 15026 55260 15370
rect 55416 15094 55444 15370
rect 55404 15088 55456 15094
rect 55404 15030 55456 15036
rect 55220 15020 55272 15026
rect 55220 14962 55272 14968
rect 54024 14952 54076 14958
rect 54024 14894 54076 14900
rect 55036 14952 55088 14958
rect 55036 14894 55088 14900
rect 54036 14074 54064 14894
rect 55048 14414 55076 14894
rect 55232 14618 55260 14962
rect 55220 14612 55272 14618
rect 55220 14554 55272 14560
rect 55036 14408 55088 14414
rect 55036 14350 55088 14356
rect 54208 14272 54260 14278
rect 54208 14214 54260 14220
rect 54220 14074 54248 14214
rect 54024 14068 54076 14074
rect 54024 14010 54076 14016
rect 54208 14068 54260 14074
rect 54208 14010 54260 14016
rect 53196 14000 53248 14006
rect 53196 13942 53248 13948
rect 53840 14000 53892 14006
rect 53840 13942 53892 13948
rect 54116 13932 54168 13938
rect 54116 13874 54168 13880
rect 53104 13864 53156 13870
rect 53104 13806 53156 13812
rect 53288 13728 53340 13734
rect 53288 13670 53340 13676
rect 53932 13728 53984 13734
rect 53932 13670 53984 13676
rect 53300 13326 53328 13670
rect 53944 13326 53972 13670
rect 53288 13320 53340 13326
rect 53288 13262 53340 13268
rect 53932 13320 53984 13326
rect 53932 13262 53984 13268
rect 54128 13258 54156 13874
rect 54576 13864 54628 13870
rect 54576 13806 54628 13812
rect 54588 13530 54616 13806
rect 54576 13524 54628 13530
rect 54576 13466 54628 13472
rect 55036 13524 55088 13530
rect 55036 13466 55088 13472
rect 54116 13252 54168 13258
rect 54116 13194 54168 13200
rect 52184 12980 52236 12986
rect 52184 12922 52236 12928
rect 52000 12368 52052 12374
rect 52000 12310 52052 12316
rect 51448 12300 51500 12306
rect 51448 12242 51500 12248
rect 51460 11762 51488 12242
rect 51540 12096 51592 12102
rect 51540 12038 51592 12044
rect 51448 11756 51500 11762
rect 51448 11698 51500 11704
rect 51356 11620 51408 11626
rect 51356 11562 51408 11568
rect 51368 11150 51396 11562
rect 51356 11144 51408 11150
rect 51356 11086 51408 11092
rect 51460 11014 51488 11698
rect 51552 11694 51580 12038
rect 52012 11762 52040 12310
rect 52196 12170 52224 12922
rect 54588 12918 54616 13466
rect 54852 13456 54904 13462
rect 54852 13398 54904 13404
rect 54864 13258 54892 13398
rect 54852 13252 54904 13258
rect 54852 13194 54904 13200
rect 54576 12912 54628 12918
rect 54576 12854 54628 12860
rect 54864 12850 54892 13194
rect 55048 12986 55076 13466
rect 55232 13394 55260 14554
rect 55600 14482 55628 15982
rect 55680 15496 55732 15502
rect 55680 15438 55732 15444
rect 55692 14618 55720 15438
rect 55772 15360 55824 15366
rect 55772 15302 55824 15308
rect 55784 15094 55812 15302
rect 55772 15088 55824 15094
rect 55772 15030 55824 15036
rect 56324 14816 56376 14822
rect 56324 14758 56376 14764
rect 55680 14612 55732 14618
rect 55680 14554 55732 14560
rect 55588 14476 55640 14482
rect 55588 14418 55640 14424
rect 55220 13388 55272 13394
rect 55220 13330 55272 13336
rect 55036 12980 55088 12986
rect 55036 12922 55088 12928
rect 55128 12912 55180 12918
rect 55128 12854 55180 12860
rect 54852 12844 54904 12850
rect 54852 12786 54904 12792
rect 54668 12640 54720 12646
rect 54668 12582 54720 12588
rect 52184 12164 52236 12170
rect 52184 12106 52236 12112
rect 53932 12096 53984 12102
rect 53932 12038 53984 12044
rect 53944 11830 53972 12038
rect 53932 11824 53984 11830
rect 53932 11766 53984 11772
rect 52000 11756 52052 11762
rect 52000 11698 52052 11704
rect 54680 11694 54708 12582
rect 55140 12238 55168 12854
rect 55404 12776 55456 12782
rect 55404 12718 55456 12724
rect 55416 12238 55444 12718
rect 55600 12306 55628 14418
rect 56336 13326 56364 14758
rect 56324 13320 56376 13326
rect 56324 13262 56376 13268
rect 56048 13252 56100 13258
rect 56048 13194 56100 13200
rect 56060 12986 56088 13194
rect 56232 13184 56284 13190
rect 56232 13126 56284 13132
rect 56048 12980 56100 12986
rect 56048 12922 56100 12928
rect 56244 12850 56272 13126
rect 56232 12844 56284 12850
rect 56232 12786 56284 12792
rect 56336 12646 56364 13262
rect 56324 12640 56376 12646
rect 56324 12582 56376 12588
rect 55588 12300 55640 12306
rect 55588 12242 55640 12248
rect 55128 12232 55180 12238
rect 55128 12174 55180 12180
rect 55404 12232 55456 12238
rect 55404 12174 55456 12180
rect 55140 11830 55168 12174
rect 55416 11898 55444 12174
rect 55404 11892 55456 11898
rect 55404 11834 55456 11840
rect 55128 11824 55180 11830
rect 55128 11766 55180 11772
rect 51540 11688 51592 11694
rect 51540 11630 51592 11636
rect 54668 11688 54720 11694
rect 54668 11630 54720 11636
rect 51552 11150 51580 11630
rect 55600 11558 55628 12242
rect 55588 11552 55640 11558
rect 55588 11494 55640 11500
rect 51632 11280 51684 11286
rect 51632 11222 51684 11228
rect 51540 11144 51592 11150
rect 51540 11086 51592 11092
rect 51448 11008 51500 11014
rect 51448 10950 51500 10956
rect 51460 10266 51488 10950
rect 51448 10260 51500 10266
rect 51448 10202 51500 10208
rect 48044 10124 48096 10130
rect 48044 10066 48096 10072
rect 51080 10124 51132 10130
rect 51080 10066 51132 10072
rect 51540 10124 51592 10130
rect 51540 10066 51592 10072
rect 48780 9988 48832 9994
rect 48780 9930 48832 9936
rect 47124 9580 47176 9586
rect 47124 9522 47176 9528
rect 47032 9376 47084 9382
rect 47032 9318 47084 9324
rect 46664 9036 46716 9042
rect 46664 8978 46716 8984
rect 46676 8838 46704 8978
rect 47044 8974 47072 9318
rect 47136 8974 47164 9522
rect 48504 9376 48556 9382
rect 48504 9318 48556 9324
rect 47032 8968 47084 8974
rect 47032 8910 47084 8916
rect 47124 8968 47176 8974
rect 47124 8910 47176 8916
rect 46572 8832 46624 8838
rect 46572 8774 46624 8780
rect 46664 8832 46716 8838
rect 46664 8774 46716 8780
rect 46480 8084 46532 8090
rect 46480 8026 46532 8032
rect 45468 7948 45520 7954
rect 45468 7890 45520 7896
rect 45928 7812 45980 7818
rect 45928 7754 45980 7760
rect 46020 7812 46072 7818
rect 46020 7754 46072 7760
rect 45940 7546 45968 7754
rect 45928 7540 45980 7546
rect 45928 7482 45980 7488
rect 45940 7410 45968 7482
rect 46032 7410 46060 7754
rect 46204 7472 46256 7478
rect 46204 7414 46256 7420
rect 44548 7404 44600 7410
rect 44548 7346 44600 7352
rect 44640 7404 44692 7410
rect 44640 7346 44692 7352
rect 45928 7404 45980 7410
rect 45928 7346 45980 7352
rect 46020 7404 46072 7410
rect 46020 7346 46072 7352
rect 44180 6860 44232 6866
rect 44180 6802 44232 6808
rect 44192 6390 44220 6802
rect 44560 6458 44588 7346
rect 45284 7200 45336 7206
rect 45284 7142 45336 7148
rect 45296 6730 45324 7142
rect 45376 6996 45428 7002
rect 45376 6938 45428 6944
rect 45388 6730 45416 6938
rect 45284 6724 45336 6730
rect 45284 6666 45336 6672
rect 45376 6724 45428 6730
rect 45376 6666 45428 6672
rect 45928 6656 45980 6662
rect 45928 6598 45980 6604
rect 44548 6452 44600 6458
rect 44548 6394 44600 6400
rect 45940 6390 45968 6598
rect 46216 6458 46244 7414
rect 47136 6798 47164 8910
rect 48228 8424 48280 8430
rect 48228 8366 48280 8372
rect 47216 7200 47268 7206
rect 47216 7142 47268 7148
rect 47228 6798 47256 7142
rect 48240 6798 48268 8366
rect 46940 6792 46992 6798
rect 46940 6734 46992 6740
rect 47124 6792 47176 6798
rect 47124 6734 47176 6740
rect 47216 6792 47268 6798
rect 47216 6734 47268 6740
rect 48228 6792 48280 6798
rect 48228 6734 48280 6740
rect 46204 6452 46256 6458
rect 46204 6394 46256 6400
rect 46848 6452 46900 6458
rect 46848 6394 46900 6400
rect 44180 6384 44232 6390
rect 44180 6326 44232 6332
rect 45928 6384 45980 6390
rect 46860 6338 46888 6394
rect 45928 6326 45980 6332
rect 43076 6316 43128 6322
rect 43076 6258 43128 6264
rect 43996 6316 44048 6322
rect 43996 6258 44048 6264
rect 44364 6316 44416 6322
rect 44364 6258 44416 6264
rect 43168 6248 43220 6254
rect 43168 6190 43220 6196
rect 42800 5568 42852 5574
rect 42800 5510 42852 5516
rect 42984 5568 43036 5574
rect 42984 5510 43036 5516
rect 42708 5296 42760 5302
rect 42708 5238 42760 5244
rect 42616 5024 42668 5030
rect 42616 4966 42668 4972
rect 42628 3942 42656 4966
rect 42720 4321 42748 5238
rect 42812 4826 42840 5510
rect 43180 5370 43208 6190
rect 43812 6112 43864 6118
rect 43812 6054 43864 6060
rect 43168 5364 43220 5370
rect 43168 5306 43220 5312
rect 42892 5296 42944 5302
rect 42892 5238 42944 5244
rect 42800 4820 42852 4826
rect 42800 4762 42852 4768
rect 42706 4312 42762 4321
rect 42706 4247 42762 4256
rect 42800 4276 42852 4282
rect 42904 4264 42932 5238
rect 42984 4616 43036 4622
rect 42984 4558 43036 4564
rect 43536 4616 43588 4622
rect 43536 4558 43588 4564
rect 42996 4282 43024 4558
rect 43548 4282 43576 4558
rect 42852 4236 42932 4264
rect 42800 4218 42852 4224
rect 42708 4208 42760 4214
rect 42708 4150 42760 4156
rect 42616 3936 42668 3942
rect 42616 3878 42668 3884
rect 42720 3534 42748 4150
rect 42904 4078 42932 4236
rect 42984 4276 43036 4282
rect 42984 4218 43036 4224
rect 43536 4276 43588 4282
rect 43536 4218 43588 4224
rect 42892 4072 42944 4078
rect 42892 4014 42944 4020
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 42720 3058 42748 3470
rect 43824 3126 43852 6054
rect 44008 3670 44036 6258
rect 44376 5302 44404 6258
rect 45376 5636 45428 5642
rect 45376 5578 45428 5584
rect 45388 5302 45416 5578
rect 44364 5296 44416 5302
rect 44364 5238 44416 5244
rect 45376 5296 45428 5302
rect 45376 5238 45428 5244
rect 45468 5024 45520 5030
rect 45468 4966 45520 4972
rect 44916 4616 44968 4622
rect 44916 4558 44968 4564
rect 44928 4321 44956 4558
rect 45376 4480 45428 4486
rect 45376 4422 45428 4428
rect 44914 4312 44970 4321
rect 44914 4247 44970 4256
rect 43996 3664 44048 3670
rect 43996 3606 44048 3612
rect 44088 3188 44140 3194
rect 44088 3130 44140 3136
rect 43812 3120 43864 3126
rect 43812 3062 43864 3068
rect 42708 3052 42760 3058
rect 42708 2994 42760 3000
rect 42616 2848 42668 2854
rect 42616 2790 42668 2796
rect 42432 2440 42484 2446
rect 42432 2382 42484 2388
rect 42064 2372 42116 2378
rect 42064 2314 42116 2320
rect 42076 800 42104 2314
rect 42628 800 42656 2790
rect 43536 2372 43588 2378
rect 43536 2314 43588 2320
rect 43548 800 43576 2314
rect 43812 2304 43864 2310
rect 43812 2246 43864 2252
rect 43824 1494 43852 2246
rect 43812 1488 43864 1494
rect 43812 1430 43864 1436
rect 44100 800 44128 3130
rect 44928 2922 44956 4247
rect 45388 3126 45416 4422
rect 45480 4078 45508 4966
rect 45940 4146 45968 6326
rect 46296 6316 46348 6322
rect 46296 6258 46348 6264
rect 46492 6310 46888 6338
rect 46020 5704 46072 5710
rect 46020 5646 46072 5652
rect 46032 4146 46060 5646
rect 46112 4616 46164 4622
rect 46112 4558 46164 4564
rect 46124 4214 46152 4558
rect 46204 4548 46256 4554
rect 46204 4490 46256 4496
rect 46112 4208 46164 4214
rect 46112 4150 46164 4156
rect 45928 4140 45980 4146
rect 45928 4082 45980 4088
rect 46020 4140 46072 4146
rect 46020 4082 46072 4088
rect 45468 4072 45520 4078
rect 45468 4014 45520 4020
rect 45836 4004 45888 4010
rect 45836 3946 45888 3952
rect 45744 3596 45796 3602
rect 45744 3538 45796 3544
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 44916 2916 44968 2922
rect 44916 2858 44968 2864
rect 45008 2372 45060 2378
rect 45008 2314 45060 2320
rect 45020 800 45048 2314
rect 45480 800 45508 3334
rect 45756 2854 45784 3538
rect 45848 2854 45876 3946
rect 45940 3126 45968 4082
rect 46032 3534 46060 4082
rect 46020 3528 46072 3534
rect 46020 3470 46072 3476
rect 46216 3398 46244 4490
rect 46308 4146 46336 6258
rect 46492 6254 46520 6310
rect 46480 6248 46532 6254
rect 46480 6190 46532 6196
rect 46388 5636 46440 5642
rect 46388 5578 46440 5584
rect 46400 4622 46428 5578
rect 46480 5160 46532 5166
rect 46480 5102 46532 5108
rect 46492 4826 46520 5102
rect 46756 5024 46808 5030
rect 46756 4966 46808 4972
rect 46480 4820 46532 4826
rect 46480 4762 46532 4768
rect 46388 4616 46440 4622
rect 46388 4558 46440 4564
rect 46296 4140 46348 4146
rect 46296 4082 46348 4088
rect 46480 4140 46532 4146
rect 46480 4082 46532 4088
rect 46492 3602 46520 4082
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 46768 3466 46796 4966
rect 46848 4480 46900 4486
rect 46848 4422 46900 4428
rect 46860 4214 46888 4422
rect 46952 4214 46980 6734
rect 48412 6656 48464 6662
rect 48412 6598 48464 6604
rect 48424 6322 48452 6598
rect 48412 6316 48464 6322
rect 48412 6258 48464 6264
rect 47124 5228 47176 5234
rect 47124 5170 47176 5176
rect 47136 4622 47164 5170
rect 48228 5160 48280 5166
rect 48228 5102 48280 5108
rect 48240 4622 48268 5102
rect 47124 4616 47176 4622
rect 47124 4558 47176 4564
rect 47400 4616 47452 4622
rect 47400 4558 47452 4564
rect 48228 4616 48280 4622
rect 48228 4558 48280 4564
rect 46848 4208 46900 4214
rect 46848 4150 46900 4156
rect 46940 4208 46992 4214
rect 46940 4150 46992 4156
rect 47412 4010 47440 4558
rect 48240 4214 48268 4558
rect 48228 4208 48280 4214
rect 48228 4150 48280 4156
rect 47400 4004 47452 4010
rect 47400 3946 47452 3952
rect 46756 3460 46808 3466
rect 46756 3402 46808 3408
rect 46204 3392 46256 3398
rect 46204 3334 46256 3340
rect 45928 3120 45980 3126
rect 45928 3062 45980 3068
rect 46216 3058 46244 3334
rect 48424 3126 48452 6258
rect 48412 3120 48464 3126
rect 48412 3062 48464 3068
rect 46204 3052 46256 3058
rect 46204 2994 46256 3000
rect 47032 2916 47084 2922
rect 47032 2858 47084 2864
rect 45744 2848 45796 2854
rect 45744 2790 45796 2796
rect 45836 2848 45888 2854
rect 45836 2790 45888 2796
rect 46480 2372 46532 2378
rect 46480 2314 46532 2320
rect 45560 2304 45612 2310
rect 45560 2246 45612 2252
rect 45572 1426 45600 2246
rect 45560 1420 45612 1426
rect 45560 1362 45612 1368
rect 46492 800 46520 2314
rect 46756 2304 46808 2310
rect 46756 2246 46808 2252
rect 46768 2038 46796 2246
rect 46756 2032 46808 2038
rect 46756 1974 46808 1980
rect 47044 1442 47072 2858
rect 48516 2446 48544 9318
rect 48596 8900 48648 8906
rect 48596 8842 48648 8848
rect 48608 8634 48636 8842
rect 48596 8628 48648 8634
rect 48596 8570 48648 8576
rect 48792 8498 48820 9930
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 49700 9648 49752 9654
rect 49700 9590 49752 9596
rect 49516 9512 49568 9518
rect 49516 9454 49568 9460
rect 49424 9376 49476 9382
rect 49424 9318 49476 9324
rect 48780 8492 48832 8498
rect 48780 8434 48832 8440
rect 48792 7410 48820 8434
rect 49436 8294 49464 9318
rect 49528 8838 49556 9454
rect 49608 9376 49660 9382
rect 49608 9318 49660 9324
rect 49516 8832 49568 8838
rect 49516 8774 49568 8780
rect 49424 8288 49476 8294
rect 49424 8230 49476 8236
rect 49424 8016 49476 8022
rect 49424 7958 49476 7964
rect 49436 7410 49464 7958
rect 48780 7404 48832 7410
rect 48780 7346 48832 7352
rect 49332 7404 49384 7410
rect 49332 7346 49384 7352
rect 49424 7404 49476 7410
rect 49424 7346 49476 7352
rect 49344 6798 49372 7346
rect 48872 6792 48924 6798
rect 48872 6734 48924 6740
rect 49332 6792 49384 6798
rect 49332 6734 49384 6740
rect 48884 6390 48912 6734
rect 48872 6384 48924 6390
rect 48778 6352 48834 6361
rect 48872 6326 48924 6332
rect 49528 6338 49556 8774
rect 49620 8498 49648 9318
rect 49712 8974 49740 9590
rect 51552 9042 51580 10066
rect 51644 10062 51672 11222
rect 51632 10056 51684 10062
rect 51632 9998 51684 10004
rect 51540 9036 51592 9042
rect 51540 8978 51592 8984
rect 49700 8968 49752 8974
rect 49700 8910 49752 8916
rect 51080 8968 51132 8974
rect 51080 8910 51132 8916
rect 49712 8634 49740 8910
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 51092 8634 51120 8910
rect 49700 8628 49752 8634
rect 49700 8570 49752 8576
rect 51080 8628 51132 8634
rect 51080 8570 51132 8576
rect 49608 8492 49660 8498
rect 49608 8434 49660 8440
rect 49700 8424 49752 8430
rect 49700 8366 49752 8372
rect 49712 8090 49740 8366
rect 49700 8084 49752 8090
rect 49700 8026 49752 8032
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 51552 7410 51580 8978
rect 52736 8832 52788 8838
rect 52736 8774 52788 8780
rect 52920 8832 52972 8838
rect 52920 8774 52972 8780
rect 52460 8492 52512 8498
rect 52460 8434 52512 8440
rect 51540 7404 51592 7410
rect 51540 7346 51592 7352
rect 49608 7336 49660 7342
rect 49608 7278 49660 7284
rect 49884 7336 49936 7342
rect 49884 7278 49936 7284
rect 49620 6458 49648 7278
rect 49700 6656 49752 6662
rect 49700 6598 49752 6604
rect 49608 6452 49660 6458
rect 49608 6394 49660 6400
rect 49528 6322 49648 6338
rect 48700 6296 48778 6304
rect 48700 6276 48780 6296
rect 48596 6180 48648 6186
rect 48700 6168 48728 6276
rect 48832 6287 48834 6296
rect 49424 6316 49476 6322
rect 48780 6258 48832 6264
rect 49528 6316 49660 6322
rect 49528 6310 49608 6316
rect 49424 6258 49476 6264
rect 49608 6258 49660 6264
rect 49436 6202 49464 6258
rect 49436 6186 49556 6202
rect 49436 6180 49568 6186
rect 49436 6174 49516 6180
rect 48648 6140 48728 6168
rect 48596 6122 48648 6128
rect 49516 6122 49568 6128
rect 49528 5642 49556 6122
rect 49516 5636 49568 5642
rect 49516 5578 49568 5584
rect 49620 3058 49648 6258
rect 49712 5234 49740 6598
rect 49790 6352 49846 6361
rect 49790 6287 49792 6296
rect 49844 6287 49846 6296
rect 49792 6258 49844 6264
rect 49896 5370 49924 7278
rect 51540 7200 51592 7206
rect 51540 7142 51592 7148
rect 51552 6866 51580 7142
rect 51540 6860 51592 6866
rect 51540 6802 51592 6808
rect 50160 6792 50212 6798
rect 50160 6734 50212 6740
rect 50068 6724 50120 6730
rect 50068 6666 50120 6672
rect 50080 5846 50108 6666
rect 50172 6458 50200 6734
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 50160 6452 50212 6458
rect 50160 6394 50212 6400
rect 50988 6384 51040 6390
rect 50988 6326 51040 6332
rect 50068 5840 50120 5846
rect 50068 5782 50120 5788
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 51000 5370 51028 6326
rect 49884 5364 49936 5370
rect 49884 5306 49936 5312
rect 50988 5364 51040 5370
rect 50988 5306 51040 5312
rect 49700 5228 49752 5234
rect 49700 5170 49752 5176
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 51000 3058 51028 5306
rect 49608 3052 49660 3058
rect 49608 2994 49660 3000
rect 50988 3052 51040 3058
rect 50988 2994 51040 3000
rect 51552 2990 51580 6802
rect 52184 6384 52236 6390
rect 52182 6352 52184 6361
rect 52236 6352 52238 6361
rect 52182 6287 52238 6296
rect 52196 5710 52224 6287
rect 52368 6180 52420 6186
rect 52368 6122 52420 6128
rect 52380 5710 52408 6122
rect 52472 5778 52500 8434
rect 52748 7886 52776 8774
rect 52932 8498 52960 8774
rect 52920 8492 52972 8498
rect 52920 8434 52972 8440
rect 54852 8424 54904 8430
rect 54852 8366 54904 8372
rect 52736 7880 52788 7886
rect 52736 7822 52788 7828
rect 53012 7880 53064 7886
rect 53012 7822 53064 7828
rect 52552 7744 52604 7750
rect 52552 7686 52604 7692
rect 52564 7478 52592 7686
rect 52552 7472 52604 7478
rect 52552 7414 52604 7420
rect 52748 6866 52776 7822
rect 52736 6860 52788 6866
rect 52736 6802 52788 6808
rect 52920 6792 52972 6798
rect 52920 6734 52972 6740
rect 52736 6316 52788 6322
rect 52736 6258 52788 6264
rect 52460 5772 52512 5778
rect 52460 5714 52512 5720
rect 52184 5704 52236 5710
rect 52184 5646 52236 5652
rect 52368 5704 52420 5710
rect 52368 5646 52420 5652
rect 52472 3126 52500 5714
rect 52748 5574 52776 6258
rect 52932 5914 52960 6734
rect 53024 6458 53052 7822
rect 54864 7546 54892 8366
rect 54852 7540 54904 7546
rect 54852 7482 54904 7488
rect 53104 7404 53156 7410
rect 53104 7346 53156 7352
rect 53012 6452 53064 6458
rect 53012 6394 53064 6400
rect 52920 5908 52972 5914
rect 52920 5850 52972 5856
rect 53116 5710 53144 7346
rect 53288 6656 53340 6662
rect 53288 6598 53340 6604
rect 53300 5710 53328 6598
rect 54864 6390 54892 7482
rect 54852 6384 54904 6390
rect 54852 6326 54904 6332
rect 53104 5704 53156 5710
rect 53104 5646 53156 5652
rect 53288 5704 53340 5710
rect 53288 5646 53340 5652
rect 52736 5568 52788 5574
rect 52736 5510 52788 5516
rect 54392 5568 54444 5574
rect 54392 5510 54444 5516
rect 52460 3120 52512 3126
rect 52460 3062 52512 3068
rect 51540 2984 51592 2990
rect 51540 2926 51592 2932
rect 49884 2848 49936 2854
rect 49884 2790 49936 2796
rect 51356 2848 51408 2854
rect 51356 2790 51408 2796
rect 52828 2848 52880 2854
rect 52828 2790 52880 2796
rect 54300 2848 54352 2854
rect 54300 2790 54352 2796
rect 48504 2440 48556 2446
rect 48504 2382 48556 2388
rect 47952 2372 48004 2378
rect 47952 2314 48004 2320
rect 49424 2372 49476 2378
rect 49424 2314 49476 2320
rect 46952 1414 47072 1442
rect 46952 800 46980 1414
rect 47964 800 47992 2314
rect 48228 2304 48280 2310
rect 48228 2246 48280 2252
rect 48412 2304 48464 2310
rect 48412 2246 48464 2252
rect 48240 1970 48268 2246
rect 48228 1964 48280 1970
rect 48228 1906 48280 1912
rect 48424 800 48452 2246
rect 49436 800 49464 2314
rect 49896 800 49924 2790
rect 50896 2372 50948 2378
rect 50896 2314 50948 2320
rect 50712 2304 50764 2310
rect 50712 2246 50764 2252
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 50724 1766 50752 2246
rect 50712 1760 50764 1766
rect 50712 1702 50764 1708
rect 50908 800 50936 2314
rect 51368 800 51396 2790
rect 52368 2440 52420 2446
rect 52368 2382 52420 2388
rect 51632 2304 51684 2310
rect 51632 2246 51684 2252
rect 51644 1834 51672 2246
rect 51632 1828 51684 1834
rect 51632 1770 51684 1776
rect 52380 800 52408 2382
rect 52840 800 52868 2790
rect 53840 2440 53892 2446
rect 53840 2382 53892 2388
rect 53012 2372 53064 2378
rect 53012 2314 53064 2320
rect 53024 1698 53052 2314
rect 53012 1692 53064 1698
rect 53012 1634 53064 1640
rect 53852 800 53880 2382
rect 54208 2372 54260 2378
rect 54208 2314 54260 2320
rect 54220 1630 54248 2314
rect 54208 1624 54260 1630
rect 54208 1566 54260 1572
rect 54312 800 54340 2790
rect 54404 2514 54432 5510
rect 54864 3194 54892 6326
rect 57152 3664 57204 3670
rect 57152 3606 57204 3612
rect 54852 3188 54904 3194
rect 54852 3130 54904 3136
rect 57164 3126 57192 3606
rect 58164 3528 58216 3534
rect 58164 3470 58216 3476
rect 57152 3120 57204 3126
rect 57152 3062 57204 3068
rect 55772 2848 55824 2854
rect 55772 2790 55824 2796
rect 54392 2508 54444 2514
rect 54392 2450 54444 2456
rect 55220 2440 55272 2446
rect 55220 2382 55272 2388
rect 55232 800 55260 2382
rect 55588 2372 55640 2378
rect 55588 2314 55640 2320
rect 55600 1902 55628 2314
rect 55588 1896 55640 1902
rect 55588 1838 55640 1844
rect 55784 800 55812 2790
rect 56692 2440 56744 2446
rect 56692 2382 56744 2388
rect 56704 800 56732 2382
rect 57060 2372 57112 2378
rect 57060 2314 57112 2320
rect 57072 1562 57100 2314
rect 57244 2304 57296 2310
rect 57244 2246 57296 2252
rect 57060 1556 57112 1562
rect 57060 1498 57112 1504
rect 57256 800 57284 2246
rect 58176 800 58204 3470
rect 59636 2984 59688 2990
rect 59636 2926 59688 2932
rect 58716 2848 58768 2854
rect 58716 2790 58768 2796
rect 58728 800 58756 2790
rect 59648 800 59676 2926
rect 22664 734 22876 762
rect 23110 0 23166 800
rect 23570 0 23626 800
rect 24030 0 24086 800
rect 24582 0 24638 800
rect 25042 0 25098 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28446 0 28502 800
rect 28906 0 28962 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31850 0 31906 800
rect 32310 0 32366 800
rect 32862 0 32918 800
rect 33322 0 33378 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34794 0 34850 800
rect 35254 0 35310 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36726 0 36782 800
rect 37186 0 37242 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39670 0 39726 800
rect 40130 0 40186 800
rect 40590 0 40646 800
rect 41142 0 41198 800
rect 41602 0 41658 800
rect 42062 0 42118 800
rect 42614 0 42670 800
rect 43074 0 43130 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44546 0 44602 800
rect 45006 0 45062 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 47950 0 48006 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49422 0 49478 800
rect 49882 0 49938 800
rect 50342 0 50398 800
rect 50894 0 50950 800
rect 51354 0 51410 800
rect 51814 0 51870 800
rect 52366 0 52422 800
rect 52826 0 52882 800
rect 53286 0 53342 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55770 0 55826 800
rect 56230 0 56286 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59174 0 59230 800
rect 59634 0 59690 800
<< via2 >>
rect 2870 41656 2926 41712
rect 2778 40024 2834 40080
rect 1398 32000 1454 32056
rect 1582 39244 1584 39264
rect 1584 39244 1636 39264
rect 1636 39244 1638 39264
rect 1582 39208 1638 39244
rect 3054 40840 3110 40896
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 1582 38392 1638 38448
rect 1582 37612 1584 37632
rect 1584 37612 1636 37632
rect 1636 37612 1638 37632
rect 1582 37576 1638 37612
rect 1582 36644 1638 36680
rect 1582 36624 1584 36644
rect 1584 36624 1636 36644
rect 1636 36624 1638 36644
rect 1582 35808 1638 35864
rect 1582 34992 1638 35048
rect 1582 33804 1584 33824
rect 1584 33804 1636 33824
rect 1636 33804 1638 33824
rect 1582 33768 1638 33804
rect 1582 32408 1638 32464
rect 1582 31592 1638 31648
rect 1582 31184 1638 31240
rect 1582 29996 1584 30016
rect 1584 29996 1636 30016
rect 1636 29996 1638 30016
rect 1582 29960 1638 29996
rect 1582 27376 1638 27432
rect 1490 27004 1492 27024
rect 1492 27004 1544 27024
rect 1544 27004 1546 27024
rect 1490 26968 1546 27004
rect 1398 25744 1454 25800
rect 1858 34584 1914 34640
rect 1858 33360 1914 33416
rect 1858 30776 1914 30832
rect 1858 29552 1914 29608
rect 1858 28328 1914 28384
rect 1582 24928 1638 24984
rect 1398 24520 1454 24576
rect 1398 23976 1454 24032
rect 1582 23704 1638 23760
rect 1398 23160 1454 23216
rect 1582 22380 1584 22400
rect 1584 22380 1636 22400
rect 1636 22380 1638 22400
rect 1582 22344 1638 22380
rect 1858 21972 1860 21992
rect 1860 21972 1912 21992
rect 1912 21972 1914 21992
rect 1858 21936 1914 21972
rect 1398 21528 1454 21584
rect 1582 21120 1638 21176
rect 1674 20712 1730 20768
rect 1582 19896 1638 19952
rect 1398 19488 1454 19544
rect 1398 18128 1454 18184
rect 1582 18536 1638 18592
rect 1582 16088 1638 16144
rect 1490 15680 1546 15736
rect 1582 14864 1638 14920
rect 1398 14456 1454 14512
rect 2318 34176 2374 34232
rect 1858 16904 1914 16960
rect 2318 26188 2320 26208
rect 2320 26188 2372 26208
rect 2372 26188 2374 26208
rect 2318 26152 2374 26188
rect 2318 25336 2374 25392
rect 2870 32952 2926 33008
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 2962 30368 3018 30424
rect 2870 29144 2926 29200
rect 2226 22752 2282 22808
rect 2870 28736 2926 28792
rect 3054 27784 3110 27840
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 3146 24112 3202 24168
rect 3698 26560 3754 26616
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 5446 24012 5448 24032
rect 5448 24012 5500 24032
rect 5500 24012 5502 24032
rect 5446 23976 5502 24012
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 3882 20304 3938 20360
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 3974 19080 4030 19136
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 2318 17312 2374 17368
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 3422 17720 3478 17776
rect 2870 16496 2926 16552
rect 2318 15272 2374 15328
rect 1582 13504 1638 13560
rect 2778 13912 2834 13968
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1582 13232 1638 13288
rect 1398 13096 1454 13152
rect 1858 11872 1914 11928
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 2778 12688 2834 12744
rect 2870 12280 2926 12336
rect 1582 11056 1638 11112
rect 1858 10648 1914 10704
rect 1582 10240 1638 10296
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 3514 11464 3570 11520
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1582 8472 1638 8528
rect 1398 8064 1454 8120
rect 1490 7248 1546 7304
rect 1398 6432 1454 6488
rect 1582 6060 1584 6080
rect 1584 6060 1636 6080
rect 1636 6060 1638 6080
rect 1582 6024 1638 6060
rect 3054 8916 3056 8936
rect 3056 8916 3108 8936
rect 3108 8916 3110 8936
rect 3054 8880 3110 8916
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 2870 7692 2872 7712
rect 2872 7692 2924 7712
rect 2924 7692 2926 7712
rect 2870 7656 2926 7692
rect 1858 5616 1914 5672
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3514 6840 3570 6896
rect 1398 1808 1454 1864
rect 2686 4392 2742 4448
rect 1858 3848 1914 3904
rect 1490 584 1546 640
rect 2870 4256 2926 4312
rect 3054 2644 3110 2680
rect 3054 2624 3056 2644
rect 3056 2624 3108 2644
rect 3108 2624 3110 2644
rect 2962 1400 3018 1456
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3790 4664 3846 4720
rect 3146 992 3202 1048
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4066 3032 4122 3088
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4066 2216 4122 2272
rect 8390 13252 8446 13288
rect 8390 13232 8392 13252
rect 8392 13232 8444 13252
rect 8444 13232 8446 13252
rect 8666 4392 8722 4448
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 2778 176 2834 232
rect 12530 10648 12586 10704
rect 13082 18672 13138 18728
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 13358 20884 13360 20904
rect 13360 20884 13412 20904
rect 13412 20884 13414 20904
rect 13358 20848 13414 20884
rect 14186 21936 14242 21992
rect 14554 20848 14610 20904
rect 13266 10648 13322 10704
rect 14554 14492 14556 14512
rect 14556 14492 14608 14512
rect 14608 14492 14610 14512
rect 14554 14456 14610 14492
rect 16210 21528 16266 21584
rect 17038 21972 17040 21992
rect 17040 21972 17092 21992
rect 17092 21972 17094 21992
rect 17038 21936 17094 21972
rect 15934 17720 15990 17776
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 16670 16788 16726 16824
rect 16670 16768 16672 16788
rect 16672 16768 16724 16788
rect 16724 16768 16726 16788
rect 17590 21528 17646 21584
rect 18050 21972 18052 21992
rect 18052 21972 18104 21992
rect 18104 21972 18106 21992
rect 18050 21936 18106 21972
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 17590 18944 17646 19000
rect 13910 4120 13966 4176
rect 13450 3168 13506 3224
rect 14462 3304 14518 3360
rect 15014 3168 15070 3224
rect 14738 2916 14794 2952
rect 14738 2896 14740 2916
rect 14740 2896 14792 2916
rect 14792 2896 14794 2916
rect 18142 18808 18198 18864
rect 18234 18420 18290 18456
rect 18234 18400 18236 18420
rect 18236 18400 18288 18420
rect 18288 18400 18290 18420
rect 18142 18128 18198 18184
rect 17774 17740 17830 17776
rect 17774 17720 17776 17740
rect 17776 17720 17828 17740
rect 17828 17720 17830 17740
rect 18510 18944 18566 19000
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 18878 18808 18934 18864
rect 18970 18692 19026 18728
rect 18970 18672 18972 18692
rect 18972 18672 19024 18692
rect 19024 18672 19026 18692
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19338 18420 19394 18456
rect 19338 18400 19340 18420
rect 19340 18400 19392 18420
rect 19392 18400 19394 18420
rect 19338 18284 19394 18320
rect 19338 18264 19340 18284
rect 19340 18264 19392 18284
rect 19392 18264 19394 18284
rect 18510 17992 18566 18048
rect 19062 17992 19118 18048
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 21730 19760 21786 19816
rect 20810 18128 20866 18184
rect 20810 17584 20866 17640
rect 20902 17448 20958 17504
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 20810 16768 20866 16824
rect 17866 14476 17922 14512
rect 17866 14456 17868 14476
rect 17868 14456 17920 14476
rect 17920 14456 17922 14476
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 15566 3476 15568 3496
rect 15568 3476 15620 3496
rect 15620 3476 15622 3496
rect 15566 3440 15622 3476
rect 16118 2760 16174 2816
rect 16486 3476 16488 3496
rect 16488 3476 16540 3496
rect 16540 3476 16542 3496
rect 16486 3440 16542 3476
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 17406 3304 17462 3360
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19338 5616 19394 5672
rect 18050 2896 18106 2952
rect 18786 3884 18788 3904
rect 18788 3884 18840 3904
rect 18840 3884 18842 3904
rect 18786 3848 18842 3884
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19522 3884 19524 3904
rect 19524 3884 19576 3904
rect 19576 3884 19578 3904
rect 19522 3848 19578 3884
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20350 9424 20406 9480
rect 20074 2796 20076 2816
rect 20076 2796 20128 2816
rect 20128 2796 20130 2816
rect 20074 2760 20130 2796
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21270 10648 21326 10704
rect 21546 12144 21602 12200
rect 21914 18128 21970 18184
rect 21822 12008 21878 12064
rect 22190 18300 22192 18320
rect 22192 18300 22244 18320
rect 22244 18300 22246 18320
rect 22190 18264 22246 18300
rect 23846 19796 23848 19816
rect 23848 19796 23900 19816
rect 23900 19796 23902 19816
rect 23846 19760 23902 19796
rect 22098 8880 22154 8936
rect 21730 8200 21786 8256
rect 22742 12144 22798 12200
rect 22926 12144 22982 12200
rect 22926 11228 22928 11248
rect 22928 11228 22980 11248
rect 22980 11228 22982 11248
rect 22926 11192 22982 11228
rect 21914 3576 21970 3632
rect 22650 5616 22706 5672
rect 24398 16904 24454 16960
rect 24398 7928 24454 7984
rect 24490 7812 24546 7848
rect 24490 7792 24492 7812
rect 24492 7792 24544 7812
rect 24544 7792 24546 7812
rect 25042 7792 25098 7848
rect 25686 16788 25742 16824
rect 26422 18128 26478 18184
rect 25686 16768 25688 16788
rect 25688 16768 25740 16788
rect 25740 16768 25742 16788
rect 25778 16396 25780 16416
rect 25780 16396 25832 16416
rect 25832 16396 25834 16416
rect 25778 16360 25834 16396
rect 25594 7948 25650 7984
rect 25594 7928 25596 7948
rect 25596 7928 25648 7948
rect 25648 7928 25650 7948
rect 26054 11212 26110 11248
rect 26054 11192 26056 11212
rect 26056 11192 26108 11212
rect 26108 11192 26110 11212
rect 26330 16360 26386 16416
rect 27158 17584 27214 17640
rect 26514 17448 26570 17504
rect 26974 12008 27030 12064
rect 25410 3576 25466 3632
rect 27894 10668 27950 10704
rect 27894 10648 27896 10668
rect 27896 10648 27948 10668
rect 27948 10648 27950 10668
rect 26882 8880 26938 8936
rect 26330 7792 26386 7848
rect 27802 7928 27858 7984
rect 27710 7284 27712 7304
rect 27712 7284 27764 7304
rect 27764 7284 27766 7304
rect 27710 7248 27766 7284
rect 27802 6996 27858 7032
rect 27802 6976 27804 6996
rect 27804 6976 27856 6996
rect 27856 6976 27858 6996
rect 28262 6976 28318 7032
rect 32034 19896 32090 19952
rect 28722 16360 28778 16416
rect 29274 16768 29330 16824
rect 29274 14864 29330 14920
rect 28630 9460 28632 9480
rect 28632 9460 28684 9480
rect 28684 9460 28686 9480
rect 28630 9424 28686 9460
rect 28906 12180 28908 12200
rect 28908 12180 28960 12200
rect 28960 12180 28962 12200
rect 28906 12144 28962 12180
rect 29274 11056 29330 11112
rect 28722 7928 28778 7984
rect 28998 8236 29000 8256
rect 29000 8236 29052 8256
rect 29052 8236 29054 8256
rect 28998 8200 29054 8236
rect 29182 7248 29238 7304
rect 28446 4120 28502 4176
rect 29826 15036 29828 15056
rect 29828 15036 29880 15056
rect 29880 15036 29882 15056
rect 29826 15000 29882 15036
rect 29458 11636 29460 11656
rect 29460 11636 29512 11656
rect 29512 11636 29514 11656
rect 29458 11600 29514 11636
rect 29918 11076 29974 11112
rect 29918 11056 29920 11076
rect 29920 11056 29972 11076
rect 29972 11056 29974 11076
rect 30378 15000 30434 15056
rect 30930 14864 30986 14920
rect 30654 6876 30656 6896
rect 30656 6876 30708 6896
rect 30708 6876 30710 6896
rect 30654 6840 30710 6876
rect 31298 8336 31354 8392
rect 31114 3576 31170 3632
rect 31298 3476 31300 3496
rect 31300 3476 31352 3496
rect 31352 3476 31354 3496
rect 31298 3440 31354 3476
rect 31574 6160 31630 6216
rect 32126 5244 32128 5264
rect 32128 5244 32180 5264
rect 32180 5244 32182 5264
rect 32126 5208 32182 5244
rect 32126 4564 32128 4584
rect 32128 4564 32180 4584
rect 32180 4564 32182 4584
rect 32126 4528 32182 4564
rect 32126 3052 32182 3088
rect 32126 3032 32128 3052
rect 32128 3032 32180 3052
rect 32180 3032 32182 3052
rect 32310 16940 32312 16960
rect 32312 16940 32364 16960
rect 32364 16940 32366 16960
rect 32310 16904 32366 16940
rect 33230 19896 33286 19952
rect 32402 6024 32458 6080
rect 32494 5752 32550 5808
rect 32494 5480 32550 5536
rect 32770 5888 32826 5944
rect 32494 4392 32550 4448
rect 32126 2488 32182 2544
rect 31942 2352 31998 2408
rect 33138 6060 33140 6080
rect 33140 6060 33192 6080
rect 33192 6060 33194 6080
rect 33138 6024 33194 6060
rect 33046 5888 33102 5944
rect 33046 5788 33048 5808
rect 33048 5788 33100 5808
rect 33100 5788 33102 5808
rect 33046 5752 33102 5788
rect 33046 3712 33102 3768
rect 32770 2080 32826 2136
rect 33598 8880 33654 8936
rect 33322 8336 33378 8392
rect 33322 7964 33324 7984
rect 33324 7964 33376 7984
rect 33376 7964 33378 7984
rect 33322 7928 33378 7964
rect 33322 5516 33324 5536
rect 33324 5516 33376 5536
rect 33376 5516 33378 5536
rect 33322 5480 33378 5516
rect 33598 5208 33654 5264
rect 33322 4120 33378 4176
rect 33322 3304 33378 3360
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34058 7928 34114 7984
rect 34058 3712 34114 3768
rect 34334 3304 34390 3360
rect 34334 3052 34390 3088
rect 34334 3032 34336 3052
rect 34336 3032 34388 3052
rect 34388 3032 34390 3052
rect 34334 2916 34390 2952
rect 34334 2896 34336 2916
rect 34336 2896 34388 2916
rect 34388 2896 34390 2916
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35990 11620 36046 11656
rect 35990 11600 35992 11620
rect 35992 11600 36044 11620
rect 36044 11600 36046 11620
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35070 11228 35072 11248
rect 35072 11228 35124 11248
rect 35124 11228 35126 11248
rect 35070 11192 35126 11228
rect 36174 11192 36230 11248
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34886 7404 34942 7440
rect 34886 7384 34888 7404
rect 34888 7384 34940 7404
rect 34940 7384 34942 7404
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34518 3984 34574 4040
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34702 4256 34758 4312
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 36266 9016 36322 9072
rect 35622 4664 35678 4720
rect 34610 3032 34666 3088
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35070 2508 35126 2544
rect 35070 2488 35072 2508
rect 35072 2488 35124 2508
rect 35124 2488 35126 2508
rect 35162 2352 35218 2408
rect 36358 6196 36360 6216
rect 36360 6196 36412 6216
rect 36412 6196 36414 6216
rect 36358 6160 36414 6196
rect 36634 8472 36690 8528
rect 36634 7384 36690 7440
rect 36634 6840 36690 6896
rect 36082 4120 36138 4176
rect 37002 8900 37058 8936
rect 37002 8880 37004 8900
rect 37004 8880 37056 8900
rect 37056 8880 37058 8900
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 38014 12300 38070 12336
rect 38014 12280 38016 12300
rect 38016 12280 38068 12300
rect 38068 12280 38070 12300
rect 38750 12280 38806 12336
rect 37554 9016 37610 9072
rect 37094 8472 37150 8528
rect 37922 8356 37978 8392
rect 37922 8336 37924 8356
rect 37924 8336 37976 8356
rect 37976 8336 37978 8356
rect 42522 11872 42578 11928
rect 38106 7928 38162 7984
rect 36542 4528 36598 4584
rect 36910 4256 36966 4312
rect 37278 3984 37334 4040
rect 39578 9152 39634 9208
rect 39670 6024 39726 6080
rect 38474 4664 38530 4720
rect 38290 4428 38292 4448
rect 38292 4428 38344 4448
rect 38344 4428 38346 4448
rect 38290 4392 38346 4428
rect 38290 4256 38346 4312
rect 36358 3440 36414 3496
rect 35530 2932 35532 2952
rect 35532 2932 35584 2952
rect 35584 2932 35586 2952
rect 35530 2896 35586 2932
rect 35898 2080 35954 2136
rect 38382 3576 38438 3632
rect 42706 9152 42762 9208
rect 42522 6024 42578 6080
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 46570 11892 46626 11928
rect 46570 11872 46572 11892
rect 46572 11872 46624 11892
rect 46624 11872 46626 11892
rect 45006 9152 45062 9208
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 42706 4256 42762 4312
rect 44914 4256 44970 4312
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 48778 6316 48834 6352
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 48778 6296 48780 6316
rect 48780 6296 48832 6316
rect 48832 6296 48834 6316
rect 49790 6316 49846 6352
rect 49790 6296 49792 6316
rect 49792 6296 49844 6316
rect 49844 6296 49846 6316
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 52182 6332 52184 6352
rect 52184 6332 52236 6352
rect 52236 6332 52238 6352
rect 52182 6296 52238 6332
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 0 41714 800 41744
rect 2865 41714 2931 41717
rect 0 41712 2931 41714
rect 0 41656 2870 41712
rect 2926 41656 2931 41712
rect 0 41654 2931 41656
rect 0 41624 800 41654
rect 2865 41651 2931 41654
rect 0 41216 800 41336
rect 0 40898 800 40928
rect 3049 40898 3115 40901
rect 0 40896 3115 40898
rect 0 40840 3054 40896
rect 3110 40840 3115 40896
rect 0 40838 3115 40840
rect 0 40808 800 40838
rect 3049 40835 3115 40838
rect 0 40400 800 40520
rect 0 40082 800 40112
rect 2773 40082 2839 40085
rect 0 40080 2839 40082
rect 0 40024 2778 40080
rect 2834 40024 2839 40080
rect 0 40022 2839 40024
rect 0 39992 800 40022
rect 2773 40019 2839 40022
rect 4208 39744 4528 39745
rect 0 39584 800 39704
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39266 800 39296
rect 1577 39266 1643 39269
rect 0 39264 1643 39266
rect 0 39208 1582 39264
rect 1638 39208 1643 39264
rect 0 39206 1643 39208
rect 0 39176 800 39206
rect 1577 39203 1643 39206
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 50288 39200 50608 39201
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 39135 50608 39136
rect 0 38768 800 38888
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38450 800 38480
rect 1577 38450 1643 38453
rect 0 38448 1643 38450
rect 0 38392 1582 38448
rect 1638 38392 1643 38448
rect 0 38390 1643 38392
rect 0 38360 800 38390
rect 1577 38387 1643 38390
rect 19568 38112 19888 38113
rect 0 37952 800 38072
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 50288 38112 50608 38113
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 38047 50608 38048
rect 0 37634 800 37664
rect 1577 37634 1643 37637
rect 0 37632 1643 37634
rect 0 37576 1582 37632
rect 1638 37576 1643 37632
rect 0 37574 1643 37576
rect 0 37544 800 37574
rect 1577 37571 1643 37574
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 0 37000 800 37120
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 0 36682 800 36712
rect 1577 36682 1643 36685
rect 0 36680 1643 36682
rect 0 36624 1582 36680
rect 1638 36624 1643 36680
rect 0 36622 1643 36624
rect 0 36592 800 36622
rect 1577 36619 1643 36622
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36184 800 36304
rect 19568 35936 19888 35937
rect 0 35866 800 35896
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 1577 35866 1643 35869
rect 0 35864 1643 35866
rect 0 35808 1582 35864
rect 1638 35808 1643 35864
rect 0 35806 1643 35808
rect 0 35776 800 35806
rect 1577 35803 1643 35806
rect 0 35368 800 35488
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 35050 800 35080
rect 1577 35050 1643 35053
rect 0 35048 1643 35050
rect 0 34992 1582 35048
rect 1638 34992 1643 35048
rect 0 34990 1643 34992
rect 0 34960 800 34990
rect 1577 34987 1643 34990
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 0 34642 800 34672
rect 1853 34642 1919 34645
rect 0 34640 1919 34642
rect 0 34584 1858 34640
rect 1914 34584 1919 34640
rect 0 34582 1919 34584
rect 0 34552 800 34582
rect 1853 34579 1919 34582
rect 4208 34304 4528 34305
rect 0 34234 800 34264
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 2313 34234 2379 34237
rect 0 34232 2379 34234
rect 0 34176 2318 34232
rect 2374 34176 2379 34232
rect 0 34174 2379 34176
rect 0 34144 800 34174
rect 2313 34171 2379 34174
rect 0 33826 800 33856
rect 1577 33826 1643 33829
rect 0 33824 1643 33826
rect 0 33768 1582 33824
rect 1638 33768 1643 33824
rect 0 33766 1643 33768
rect 0 33736 800 33766
rect 1577 33763 1643 33766
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 0 33418 800 33448
rect 1853 33418 1919 33421
rect 0 33416 1919 33418
rect 0 33360 1858 33416
rect 1914 33360 1919 33416
rect 0 33358 1919 33360
rect 0 33328 800 33358
rect 1853 33355 1919 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 33010 800 33040
rect 2865 33010 2931 33013
rect 0 33008 2931 33010
rect 0 32952 2870 33008
rect 2926 32952 2931 33008
rect 0 32950 2931 32952
rect 0 32920 800 32950
rect 2865 32947 2931 32950
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 0 32466 800 32496
rect 1577 32466 1643 32469
rect 0 32464 1643 32466
rect 0 32408 1582 32464
rect 1638 32408 1643 32464
rect 0 32406 1643 32408
rect 0 32376 800 32406
rect 1577 32403 1643 32406
rect 4208 32128 4528 32129
rect 0 32058 800 32088
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 1393 32058 1459 32061
rect 0 32056 1459 32058
rect 0 32000 1398 32056
rect 1454 32000 1459 32056
rect 0 31998 1459 32000
rect 0 31968 800 31998
rect 1393 31995 1459 31998
rect 0 31650 800 31680
rect 1577 31650 1643 31653
rect 0 31648 1643 31650
rect 0 31592 1582 31648
rect 1638 31592 1643 31648
rect 0 31590 1643 31592
rect 0 31560 800 31590
rect 1577 31587 1643 31590
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 0 31242 800 31272
rect 1577 31242 1643 31245
rect 0 31240 1643 31242
rect 0 31184 1582 31240
rect 1638 31184 1643 31240
rect 0 31182 1643 31184
rect 0 31152 800 31182
rect 1577 31179 1643 31182
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30834 800 30864
rect 1853 30834 1919 30837
rect 0 30832 1919 30834
rect 0 30776 1858 30832
rect 1914 30776 1919 30832
rect 0 30774 1919 30776
rect 0 30744 800 30774
rect 1853 30771 1919 30774
rect 19568 30496 19888 30497
rect 0 30426 800 30456
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 2957 30426 3023 30429
rect 0 30424 3023 30426
rect 0 30368 2962 30424
rect 3018 30368 3023 30424
rect 0 30366 3023 30368
rect 0 30336 800 30366
rect 2957 30363 3023 30366
rect 0 30018 800 30048
rect 1577 30018 1643 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 800 29958
rect 1577 29955 1643 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 0 29610 800 29640
rect 1853 29610 1919 29613
rect 0 29608 1919 29610
rect 0 29552 1858 29608
rect 1914 29552 1919 29608
rect 0 29550 1919 29552
rect 0 29520 800 29550
rect 1853 29547 1919 29550
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 0 29202 800 29232
rect 2865 29202 2931 29205
rect 0 29200 2931 29202
rect 0 29144 2870 29200
rect 2926 29144 2931 29200
rect 0 29142 2931 29144
rect 0 29112 800 29142
rect 2865 29139 2931 29142
rect 4208 28864 4528 28865
rect 0 28794 800 28824
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 2865 28794 2931 28797
rect 0 28792 2931 28794
rect 0 28736 2870 28792
rect 2926 28736 2931 28792
rect 0 28734 2931 28736
rect 0 28704 800 28734
rect 2865 28731 2931 28734
rect 0 28386 800 28416
rect 1853 28386 1919 28389
rect 0 28384 1919 28386
rect 0 28328 1858 28384
rect 1914 28328 1919 28384
rect 0 28326 1919 28328
rect 0 28296 800 28326
rect 1853 28323 1919 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 0 27842 800 27872
rect 3049 27842 3115 27845
rect 0 27840 3115 27842
rect 0 27784 3054 27840
rect 3110 27784 3115 27840
rect 0 27782 3115 27784
rect 0 27752 800 27782
rect 3049 27779 3115 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27434 800 27464
rect 1577 27434 1643 27437
rect 0 27432 1643 27434
rect 0 27376 1582 27432
rect 1638 27376 1643 27432
rect 0 27374 1643 27376
rect 0 27344 800 27374
rect 1577 27371 1643 27374
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 0 27026 800 27056
rect 1485 27026 1551 27029
rect 0 27024 1551 27026
rect 0 26968 1490 27024
rect 1546 26968 1551 27024
rect 0 26966 1551 26968
rect 0 26936 800 26966
rect 1485 26963 1551 26966
rect 4208 26688 4528 26689
rect 0 26618 800 26648
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 3693 26618 3759 26621
rect 0 26616 3759 26618
rect 0 26560 3698 26616
rect 3754 26560 3759 26616
rect 0 26558 3759 26560
rect 0 26528 800 26558
rect 3693 26555 3759 26558
rect 0 26210 800 26240
rect 2313 26210 2379 26213
rect 0 26208 2379 26210
rect 0 26152 2318 26208
rect 2374 26152 2379 26208
rect 0 26150 2379 26152
rect 0 26120 800 26150
rect 2313 26147 2379 26150
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 0 25802 800 25832
rect 1393 25802 1459 25805
rect 0 25800 1459 25802
rect 0 25744 1398 25800
rect 1454 25744 1459 25800
rect 0 25742 1459 25744
rect 0 25712 800 25742
rect 1393 25739 1459 25742
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25394 800 25424
rect 2313 25394 2379 25397
rect 0 25392 2379 25394
rect 0 25336 2318 25392
rect 2374 25336 2379 25392
rect 0 25334 2379 25336
rect 0 25304 800 25334
rect 2313 25331 2379 25334
rect 19568 25056 19888 25057
rect 0 24986 800 25016
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 1577 24986 1643 24989
rect 0 24984 1643 24986
rect 0 24928 1582 24984
rect 1638 24928 1643 24984
rect 0 24926 1643 24928
rect 0 24896 800 24926
rect 1577 24923 1643 24926
rect 0 24578 800 24608
rect 1393 24578 1459 24581
rect 0 24576 1459 24578
rect 0 24520 1398 24576
rect 1454 24520 1459 24576
rect 0 24518 1459 24520
rect 0 24488 800 24518
rect 1393 24515 1459 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 0 24170 800 24200
rect 3141 24170 3207 24173
rect 0 24168 3207 24170
rect 0 24112 3146 24168
rect 3202 24112 3207 24168
rect 0 24110 3207 24112
rect 0 24080 800 24110
rect 3141 24107 3207 24110
rect 1393 24034 1459 24037
rect 5441 24034 5507 24037
rect 1393 24032 5507 24034
rect 1393 23976 1398 24032
rect 1454 23976 5446 24032
rect 5502 23976 5507 24032
rect 1393 23974 5507 23976
rect 1393 23971 1459 23974
rect 5441 23971 5507 23974
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 0 23762 800 23792
rect 1577 23762 1643 23765
rect 0 23760 1643 23762
rect 0 23704 1582 23760
rect 1638 23704 1643 23760
rect 0 23702 1643 23704
rect 0 23672 800 23702
rect 1577 23699 1643 23702
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 19568 22880 19888 22881
rect 0 22810 800 22840
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 2221 22810 2287 22813
rect 0 22808 2287 22810
rect 0 22752 2226 22808
rect 2282 22752 2287 22808
rect 0 22750 2287 22752
rect 0 22720 800 22750
rect 2221 22747 2287 22750
rect 0 22402 800 22432
rect 1577 22402 1643 22405
rect 0 22400 1643 22402
rect 0 22344 1582 22400
rect 1638 22344 1643 22400
rect 0 22342 1643 22344
rect 0 22312 800 22342
rect 1577 22339 1643 22342
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21994 800 22024
rect 1853 21994 1919 21997
rect 0 21992 1919 21994
rect 0 21936 1858 21992
rect 1914 21936 1919 21992
rect 0 21934 1919 21936
rect 0 21904 800 21934
rect 1853 21931 1919 21934
rect 14181 21994 14247 21997
rect 17033 21994 17099 21997
rect 18045 21994 18111 21997
rect 14181 21992 18111 21994
rect 14181 21936 14186 21992
rect 14242 21936 17038 21992
rect 17094 21936 18050 21992
rect 18106 21936 18111 21992
rect 14181 21934 18111 21936
rect 14181 21931 14247 21934
rect 17033 21931 17099 21934
rect 18045 21931 18111 21934
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 0 21586 800 21616
rect 1393 21586 1459 21589
rect 0 21584 1459 21586
rect 0 21528 1398 21584
rect 1454 21528 1459 21584
rect 0 21526 1459 21528
rect 0 21496 800 21526
rect 1393 21523 1459 21526
rect 16205 21586 16271 21589
rect 17585 21586 17651 21589
rect 16205 21584 17651 21586
rect 16205 21528 16210 21584
rect 16266 21528 17590 21584
rect 17646 21528 17651 21584
rect 16205 21526 17651 21528
rect 16205 21523 16271 21526
rect 17585 21523 17651 21526
rect 4208 21248 4528 21249
rect 0 21178 800 21208
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 1577 21178 1643 21181
rect 0 21176 1643 21178
rect 0 21120 1582 21176
rect 1638 21120 1643 21176
rect 0 21118 1643 21120
rect 0 21088 800 21118
rect 1577 21115 1643 21118
rect 13353 20906 13419 20909
rect 14549 20906 14615 20909
rect 13353 20904 14615 20906
rect 13353 20848 13358 20904
rect 13414 20848 14554 20904
rect 14610 20848 14615 20904
rect 13353 20846 14615 20848
rect 13353 20843 13419 20846
rect 14549 20843 14615 20846
rect 0 20770 800 20800
rect 1669 20770 1735 20773
rect 0 20768 1735 20770
rect 0 20712 1674 20768
rect 1730 20712 1735 20768
rect 0 20710 1735 20712
rect 0 20680 800 20710
rect 1669 20707 1735 20710
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19954 800 19984
rect 1577 19954 1643 19957
rect 0 19952 1643 19954
rect 0 19896 1582 19952
rect 1638 19896 1643 19952
rect 0 19894 1643 19896
rect 0 19864 800 19894
rect 1577 19891 1643 19894
rect 32029 19954 32095 19957
rect 33225 19954 33291 19957
rect 32029 19952 33291 19954
rect 32029 19896 32034 19952
rect 32090 19896 33230 19952
rect 33286 19896 33291 19952
rect 32029 19894 33291 19896
rect 32029 19891 32095 19894
rect 33225 19891 33291 19894
rect 21725 19818 21791 19821
rect 23841 19818 23907 19821
rect 21725 19816 23907 19818
rect 21725 19760 21730 19816
rect 21786 19760 23846 19816
rect 23902 19760 23907 19816
rect 21725 19758 23907 19760
rect 21725 19755 21791 19758
rect 23841 19755 23907 19758
rect 19568 19616 19888 19617
rect 0 19546 800 19576
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 1393 19546 1459 19549
rect 0 19544 1459 19546
rect 0 19488 1398 19544
rect 1454 19488 1459 19544
rect 0 19486 1459 19488
rect 0 19456 800 19486
rect 1393 19483 1459 19486
rect 0 19138 800 19168
rect 3969 19138 4035 19141
rect 0 19136 4035 19138
rect 0 19080 3974 19136
rect 4030 19080 4035 19136
rect 0 19078 4035 19080
rect 0 19048 800 19078
rect 3969 19075 4035 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 17585 19002 17651 19005
rect 18505 19002 18571 19005
rect 17585 19000 18571 19002
rect 17585 18944 17590 19000
rect 17646 18944 18510 19000
rect 18566 18944 18571 19000
rect 17585 18942 18571 18944
rect 17585 18939 17651 18942
rect 18505 18939 18571 18942
rect 18137 18866 18203 18869
rect 18873 18866 18939 18869
rect 18137 18864 18939 18866
rect 18137 18808 18142 18864
rect 18198 18808 18878 18864
rect 18934 18808 18939 18864
rect 18137 18806 18939 18808
rect 18137 18803 18203 18806
rect 18873 18803 18939 18806
rect 13077 18730 13143 18733
rect 18965 18730 19031 18733
rect 13077 18728 19031 18730
rect 13077 18672 13082 18728
rect 13138 18672 18970 18728
rect 19026 18672 19031 18728
rect 13077 18670 19031 18672
rect 13077 18667 13143 18670
rect 18965 18667 19031 18670
rect 0 18594 800 18624
rect 1577 18594 1643 18597
rect 0 18592 1643 18594
rect 0 18536 1582 18592
rect 1638 18536 1643 18592
rect 0 18534 1643 18536
rect 0 18504 800 18534
rect 1577 18531 1643 18534
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 18229 18458 18295 18461
rect 19333 18458 19399 18461
rect 18229 18456 19399 18458
rect 18229 18400 18234 18456
rect 18290 18400 19338 18456
rect 19394 18400 19399 18456
rect 18229 18398 19399 18400
rect 18229 18395 18295 18398
rect 19333 18395 19399 18398
rect 19333 18322 19399 18325
rect 22185 18322 22251 18325
rect 19333 18320 22251 18322
rect 19333 18264 19338 18320
rect 19394 18264 22190 18320
rect 22246 18264 22251 18320
rect 19333 18262 22251 18264
rect 19333 18259 19399 18262
rect 22185 18259 22251 18262
rect 0 18186 800 18216
rect 1393 18186 1459 18189
rect 0 18184 1459 18186
rect 0 18128 1398 18184
rect 1454 18128 1459 18184
rect 0 18126 1459 18128
rect 0 18096 800 18126
rect 1393 18123 1459 18126
rect 18137 18186 18203 18189
rect 20805 18186 20871 18189
rect 18137 18184 20871 18186
rect 18137 18128 18142 18184
rect 18198 18128 20810 18184
rect 20866 18128 20871 18184
rect 18137 18126 20871 18128
rect 18137 18123 18203 18126
rect 20805 18123 20871 18126
rect 21909 18186 21975 18189
rect 26417 18186 26483 18189
rect 21909 18184 26483 18186
rect 21909 18128 21914 18184
rect 21970 18128 26422 18184
rect 26478 18128 26483 18184
rect 21909 18126 26483 18128
rect 21909 18123 21975 18126
rect 26417 18123 26483 18126
rect 18505 18050 18571 18053
rect 19057 18050 19123 18053
rect 18505 18048 19123 18050
rect 18505 17992 18510 18048
rect 18566 17992 19062 18048
rect 19118 17992 19123 18048
rect 18505 17990 19123 17992
rect 18505 17987 18571 17990
rect 19057 17987 19123 17990
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17808
rect 3417 17778 3483 17781
rect 0 17776 3483 17778
rect 0 17720 3422 17776
rect 3478 17720 3483 17776
rect 0 17718 3483 17720
rect 0 17688 800 17718
rect 3417 17715 3483 17718
rect 15929 17778 15995 17781
rect 17769 17778 17835 17781
rect 15929 17776 17835 17778
rect 15929 17720 15934 17776
rect 15990 17720 17774 17776
rect 17830 17720 17835 17776
rect 15929 17718 17835 17720
rect 15929 17715 15995 17718
rect 17769 17715 17835 17718
rect 20805 17642 20871 17645
rect 27153 17642 27219 17645
rect 20805 17640 27219 17642
rect 20805 17584 20810 17640
rect 20866 17584 27158 17640
rect 27214 17584 27219 17640
rect 20805 17582 27219 17584
rect 20805 17579 20871 17582
rect 27153 17579 27219 17582
rect 20897 17506 20963 17509
rect 26509 17506 26575 17509
rect 20897 17504 26575 17506
rect 20897 17448 20902 17504
rect 20958 17448 26514 17504
rect 26570 17448 26575 17504
rect 20897 17446 26575 17448
rect 20897 17443 20963 17446
rect 26509 17443 26575 17446
rect 19568 17440 19888 17441
rect 0 17370 800 17400
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 2313 17370 2379 17373
rect 0 17368 2379 17370
rect 0 17312 2318 17368
rect 2374 17312 2379 17368
rect 0 17310 2379 17312
rect 0 17280 800 17310
rect 2313 17307 2379 17310
rect 0 16962 800 16992
rect 1853 16962 1919 16965
rect 0 16960 1919 16962
rect 0 16904 1858 16960
rect 1914 16904 1919 16960
rect 0 16902 1919 16904
rect 0 16872 800 16902
rect 1853 16899 1919 16902
rect 24393 16962 24459 16965
rect 32305 16962 32371 16965
rect 24393 16960 32371 16962
rect 24393 16904 24398 16960
rect 24454 16904 32310 16960
rect 32366 16904 32371 16960
rect 24393 16902 32371 16904
rect 24393 16899 24459 16902
rect 32305 16899 32371 16902
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 16665 16826 16731 16829
rect 20805 16826 20871 16829
rect 16665 16824 20871 16826
rect 16665 16768 16670 16824
rect 16726 16768 20810 16824
rect 20866 16768 20871 16824
rect 16665 16766 20871 16768
rect 16665 16763 16731 16766
rect 20805 16763 20871 16766
rect 25681 16826 25747 16829
rect 29269 16826 29335 16829
rect 25681 16824 29335 16826
rect 25681 16768 25686 16824
rect 25742 16768 29274 16824
rect 29330 16768 29335 16824
rect 25681 16766 29335 16768
rect 25681 16763 25747 16766
rect 29269 16763 29335 16766
rect 0 16554 800 16584
rect 2865 16554 2931 16557
rect 0 16552 2931 16554
rect 0 16496 2870 16552
rect 2926 16496 2931 16552
rect 0 16494 2931 16496
rect 0 16464 800 16494
rect 2865 16491 2931 16494
rect 25773 16418 25839 16421
rect 26325 16418 26391 16421
rect 28717 16418 28783 16421
rect 25773 16416 28783 16418
rect 25773 16360 25778 16416
rect 25834 16360 26330 16416
rect 26386 16360 28722 16416
rect 28778 16360 28783 16416
rect 25773 16358 28783 16360
rect 25773 16355 25839 16358
rect 26325 16355 26391 16358
rect 28717 16355 28783 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 16287 50608 16288
rect 0 16146 800 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 4208 15808 4528 15809
rect 0 15738 800 15768
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 1485 15738 1551 15741
rect 0 15736 1551 15738
rect 0 15680 1490 15736
rect 1546 15680 1551 15736
rect 0 15678 1551 15680
rect 0 15648 800 15678
rect 1485 15675 1551 15678
rect 0 15330 800 15360
rect 2313 15330 2379 15333
rect 0 15328 2379 15330
rect 0 15272 2318 15328
rect 2374 15272 2379 15328
rect 0 15270 2379 15272
rect 0 15240 800 15270
rect 2313 15267 2379 15270
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 29821 15058 29887 15061
rect 30373 15058 30439 15061
rect 29821 15056 30439 15058
rect 29821 15000 29826 15056
rect 29882 15000 30378 15056
rect 30434 15000 30439 15056
rect 29821 14998 30439 15000
rect 29821 14995 29887 14998
rect 30373 14995 30439 14998
rect 0 14922 800 14952
rect 1577 14922 1643 14925
rect 0 14920 1643 14922
rect 0 14864 1582 14920
rect 1638 14864 1643 14920
rect 0 14862 1643 14864
rect 0 14832 800 14862
rect 1577 14859 1643 14862
rect 29269 14922 29335 14925
rect 30925 14922 30991 14925
rect 29269 14920 30991 14922
rect 29269 14864 29274 14920
rect 29330 14864 30930 14920
rect 30986 14864 30991 14920
rect 29269 14862 30991 14864
rect 29269 14859 29335 14862
rect 30925 14859 30991 14862
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14514 800 14544
rect 1393 14514 1459 14517
rect 0 14512 1459 14514
rect 0 14456 1398 14512
rect 1454 14456 1459 14512
rect 0 14454 1459 14456
rect 0 14424 800 14454
rect 1393 14451 1459 14454
rect 14549 14514 14615 14517
rect 17861 14514 17927 14517
rect 14549 14512 17927 14514
rect 14549 14456 14554 14512
rect 14610 14456 17866 14512
rect 17922 14456 17927 14512
rect 14549 14454 17927 14456
rect 14549 14451 14615 14454
rect 17861 14451 17927 14454
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 0 13970 800 14000
rect 2773 13970 2839 13973
rect 0 13968 2839 13970
rect 0 13912 2778 13968
rect 2834 13912 2839 13968
rect 0 13910 2839 13912
rect 0 13880 800 13910
rect 2773 13907 2839 13910
rect 4208 13632 4528 13633
rect 0 13562 800 13592
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 1577 13562 1643 13565
rect 0 13560 1643 13562
rect 0 13504 1582 13560
rect 1638 13504 1643 13560
rect 0 13502 1643 13504
rect 0 13472 800 13502
rect 1577 13499 1643 13502
rect 1577 13290 1643 13293
rect 8385 13290 8451 13293
rect 1577 13288 8451 13290
rect 1577 13232 1582 13288
rect 1638 13232 8390 13288
rect 8446 13232 8451 13288
rect 1577 13230 8451 13232
rect 1577 13227 1643 13230
rect 8385 13227 8451 13230
rect 0 13154 800 13184
rect 1393 13154 1459 13157
rect 0 13152 1459 13154
rect 0 13096 1398 13152
rect 1454 13096 1459 13152
rect 0 13094 1459 13096
rect 0 13064 800 13094
rect 1393 13091 1459 13094
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 0 12746 800 12776
rect 2773 12746 2839 12749
rect 0 12744 2839 12746
rect 0 12688 2778 12744
rect 2834 12688 2839 12744
rect 0 12686 2839 12688
rect 0 12656 800 12686
rect 2773 12683 2839 12686
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12368
rect 2865 12338 2931 12341
rect 0 12336 2931 12338
rect 0 12280 2870 12336
rect 2926 12280 2931 12336
rect 0 12278 2931 12280
rect 0 12248 800 12278
rect 2865 12275 2931 12278
rect 38009 12338 38075 12341
rect 38745 12338 38811 12341
rect 38009 12336 38811 12338
rect 38009 12280 38014 12336
rect 38070 12280 38750 12336
rect 38806 12280 38811 12336
rect 38009 12278 38811 12280
rect 38009 12275 38075 12278
rect 38745 12275 38811 12278
rect 21541 12202 21607 12205
rect 22737 12202 22803 12205
rect 21541 12200 22803 12202
rect 21541 12144 21546 12200
rect 21602 12144 22742 12200
rect 22798 12144 22803 12200
rect 21541 12142 22803 12144
rect 21541 12139 21607 12142
rect 22737 12139 22803 12142
rect 22921 12202 22987 12205
rect 28901 12202 28967 12205
rect 22921 12200 28967 12202
rect 22921 12144 22926 12200
rect 22982 12144 28906 12200
rect 28962 12144 28967 12200
rect 22921 12142 28967 12144
rect 22921 12139 22987 12142
rect 28901 12139 28967 12142
rect 21817 12066 21883 12069
rect 26969 12066 27035 12069
rect 21817 12064 27035 12066
rect 21817 12008 21822 12064
rect 21878 12008 26974 12064
rect 27030 12008 27035 12064
rect 21817 12006 27035 12008
rect 21817 12003 21883 12006
rect 26969 12003 27035 12006
rect 19568 12000 19888 12001
rect 0 11930 800 11960
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 1853 11930 1919 11933
rect 0 11928 1919 11930
rect 0 11872 1858 11928
rect 1914 11872 1919 11928
rect 0 11870 1919 11872
rect 0 11840 800 11870
rect 1853 11867 1919 11870
rect 42517 11930 42583 11933
rect 46565 11930 46631 11933
rect 42517 11928 46631 11930
rect 42517 11872 42522 11928
rect 42578 11872 46570 11928
rect 46626 11872 46631 11928
rect 42517 11870 46631 11872
rect 42517 11867 42583 11870
rect 46565 11867 46631 11870
rect 29453 11658 29519 11661
rect 35985 11658 36051 11661
rect 29453 11656 36051 11658
rect 29453 11600 29458 11656
rect 29514 11600 35990 11656
rect 36046 11600 36051 11656
rect 29453 11598 36051 11600
rect 29453 11595 29519 11598
rect 35985 11595 36051 11598
rect 0 11522 800 11552
rect 3509 11522 3575 11525
rect 0 11520 3575 11522
rect 0 11464 3514 11520
rect 3570 11464 3575 11520
rect 0 11462 3575 11464
rect 0 11432 800 11462
rect 3509 11459 3575 11462
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 22921 11250 22987 11253
rect 26049 11250 26115 11253
rect 22921 11248 26115 11250
rect 22921 11192 22926 11248
rect 22982 11192 26054 11248
rect 26110 11192 26115 11248
rect 22921 11190 26115 11192
rect 22921 11187 22987 11190
rect 26049 11187 26115 11190
rect 35065 11250 35131 11253
rect 36169 11250 36235 11253
rect 35065 11248 36235 11250
rect 35065 11192 35070 11248
rect 35126 11192 36174 11248
rect 36230 11192 36235 11248
rect 35065 11190 36235 11192
rect 35065 11187 35131 11190
rect 36169 11187 36235 11190
rect 0 11114 800 11144
rect 1577 11114 1643 11117
rect 0 11112 1643 11114
rect 0 11056 1582 11112
rect 1638 11056 1643 11112
rect 0 11054 1643 11056
rect 0 11024 800 11054
rect 1577 11051 1643 11054
rect 29269 11114 29335 11117
rect 29913 11114 29979 11117
rect 29269 11112 29979 11114
rect 29269 11056 29274 11112
rect 29330 11056 29918 11112
rect 29974 11056 29979 11112
rect 29269 11054 29979 11056
rect 29269 11051 29335 11054
rect 29913 11051 29979 11054
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 0 10706 800 10736
rect 1853 10706 1919 10709
rect 0 10704 1919 10706
rect 0 10648 1858 10704
rect 1914 10648 1919 10704
rect 0 10646 1919 10648
rect 0 10616 800 10646
rect 1853 10643 1919 10646
rect 12525 10706 12591 10709
rect 13261 10706 13327 10709
rect 12525 10704 13327 10706
rect 12525 10648 12530 10704
rect 12586 10648 13266 10704
rect 13322 10648 13327 10704
rect 12525 10646 13327 10648
rect 12525 10643 12591 10646
rect 13261 10643 13327 10646
rect 21265 10706 21331 10709
rect 27889 10706 27955 10709
rect 21265 10704 27955 10706
rect 21265 10648 21270 10704
rect 21326 10648 27894 10704
rect 27950 10648 27955 10704
rect 21265 10646 27955 10648
rect 21265 10643 21331 10646
rect 27889 10643 27955 10646
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 1577 10298 1643 10301
rect 0 10296 1643 10298
rect 0 10240 1582 10296
rect 1638 10240 1643 10296
rect 0 10238 1643 10240
rect 0 10208 800 10238
rect 1577 10235 1643 10238
rect 0 9800 800 9920
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 20345 9482 20411 9485
rect 28625 9482 28691 9485
rect 20345 9480 28691 9482
rect 20345 9424 20350 9480
rect 20406 9424 28630 9480
rect 28686 9424 28691 9480
rect 20345 9422 28691 9424
rect 20345 9419 20411 9422
rect 28625 9419 28691 9422
rect 0 9346 800 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 800 9286
rect 1577 9283 1643 9286
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 39573 9210 39639 9213
rect 42701 9210 42767 9213
rect 45001 9210 45067 9213
rect 39573 9208 45067 9210
rect 39573 9152 39578 9208
rect 39634 9152 42706 9208
rect 42762 9152 45006 9208
rect 45062 9152 45067 9208
rect 39573 9150 45067 9152
rect 39573 9147 39639 9150
rect 42701 9147 42767 9150
rect 45001 9147 45067 9150
rect 36261 9074 36327 9077
rect 37549 9074 37615 9077
rect 36261 9072 37615 9074
rect 36261 9016 36266 9072
rect 36322 9016 37554 9072
rect 37610 9016 37615 9072
rect 36261 9014 37615 9016
rect 36261 9011 36327 9014
rect 37549 9011 37615 9014
rect 0 8938 800 8968
rect 3049 8938 3115 8941
rect 0 8936 3115 8938
rect 0 8880 3054 8936
rect 3110 8880 3115 8936
rect 0 8878 3115 8880
rect 0 8848 800 8878
rect 3049 8875 3115 8878
rect 22093 8938 22159 8941
rect 26877 8938 26943 8941
rect 22093 8936 26943 8938
rect 22093 8880 22098 8936
rect 22154 8880 26882 8936
rect 26938 8880 26943 8936
rect 22093 8878 26943 8880
rect 22093 8875 22159 8878
rect 26877 8875 26943 8878
rect 33593 8938 33659 8941
rect 36997 8938 37063 8941
rect 33593 8936 37063 8938
rect 33593 8880 33598 8936
rect 33654 8880 37002 8936
rect 37058 8880 37063 8936
rect 33593 8878 37063 8880
rect 33593 8875 33659 8878
rect 36997 8875 37063 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 0 8530 800 8560
rect 1577 8530 1643 8533
rect 0 8528 1643 8530
rect 0 8472 1582 8528
rect 1638 8472 1643 8528
rect 0 8470 1643 8472
rect 0 8440 800 8470
rect 1577 8467 1643 8470
rect 36629 8530 36695 8533
rect 37089 8530 37155 8533
rect 36629 8528 37155 8530
rect 36629 8472 36634 8528
rect 36690 8472 37094 8528
rect 37150 8472 37155 8528
rect 36629 8470 37155 8472
rect 36629 8467 36695 8470
rect 37089 8467 37155 8470
rect 31293 8394 31359 8397
rect 33317 8394 33383 8397
rect 37917 8394 37983 8397
rect 31293 8392 37983 8394
rect 31293 8336 31298 8392
rect 31354 8336 33322 8392
rect 33378 8336 37922 8392
rect 37978 8336 37983 8392
rect 31293 8334 37983 8336
rect 31293 8331 31359 8334
rect 33317 8331 33383 8334
rect 37917 8331 37983 8334
rect 21725 8258 21791 8261
rect 28993 8258 29059 8261
rect 21725 8256 29059 8258
rect 21725 8200 21730 8256
rect 21786 8200 28998 8256
rect 29054 8200 29059 8256
rect 21725 8198 29059 8200
rect 21725 8195 21791 8198
rect 28993 8195 29059 8198
rect 4208 8192 4528 8193
rect 0 8122 800 8152
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 1393 8122 1459 8125
rect 0 8120 1459 8122
rect 0 8064 1398 8120
rect 1454 8064 1459 8120
rect 0 8062 1459 8064
rect 0 8032 800 8062
rect 1393 8059 1459 8062
rect 24393 7986 24459 7989
rect 25589 7986 25655 7989
rect 27797 7986 27863 7989
rect 28717 7986 28783 7989
rect 24393 7984 28783 7986
rect 24393 7928 24398 7984
rect 24454 7928 25594 7984
rect 25650 7928 27802 7984
rect 27858 7928 28722 7984
rect 28778 7928 28783 7984
rect 24393 7926 28783 7928
rect 24393 7923 24459 7926
rect 25589 7923 25655 7926
rect 27797 7923 27863 7926
rect 28717 7923 28783 7926
rect 33317 7986 33383 7989
rect 34053 7986 34119 7989
rect 38101 7986 38167 7989
rect 33317 7984 38167 7986
rect 33317 7928 33322 7984
rect 33378 7928 34058 7984
rect 34114 7928 38106 7984
rect 38162 7928 38167 7984
rect 33317 7926 38167 7928
rect 33317 7923 33383 7926
rect 34053 7923 34119 7926
rect 38101 7923 38167 7926
rect 24485 7850 24551 7853
rect 25037 7850 25103 7853
rect 26325 7850 26391 7853
rect 24485 7848 26391 7850
rect 24485 7792 24490 7848
rect 24546 7792 25042 7848
rect 25098 7792 26330 7848
rect 26386 7792 26391 7848
rect 24485 7790 26391 7792
rect 24485 7787 24551 7790
rect 25037 7787 25103 7790
rect 26325 7787 26391 7790
rect 0 7714 800 7744
rect 2865 7714 2931 7717
rect 0 7712 2931 7714
rect 0 7656 2870 7712
rect 2926 7656 2931 7712
rect 0 7654 2931 7656
rect 0 7624 800 7654
rect 2865 7651 2931 7654
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 34881 7442 34947 7445
rect 36629 7442 36695 7445
rect 34881 7440 36695 7442
rect 34881 7384 34886 7440
rect 34942 7384 36634 7440
rect 36690 7384 36695 7440
rect 34881 7382 36695 7384
rect 34881 7379 34947 7382
rect 36629 7379 36695 7382
rect 0 7306 800 7336
rect 1485 7306 1551 7309
rect 0 7304 1551 7306
rect 0 7248 1490 7304
rect 1546 7248 1551 7304
rect 0 7246 1551 7248
rect 0 7216 800 7246
rect 1485 7243 1551 7246
rect 27705 7306 27771 7309
rect 29177 7306 29243 7309
rect 27705 7304 29243 7306
rect 27705 7248 27710 7304
rect 27766 7248 29182 7304
rect 29238 7248 29243 7304
rect 27705 7246 29243 7248
rect 27705 7243 27771 7246
rect 29177 7243 29243 7246
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 27797 7034 27863 7037
rect 28257 7034 28323 7037
rect 27797 7032 28323 7034
rect 27797 6976 27802 7032
rect 27858 6976 28262 7032
rect 28318 6976 28323 7032
rect 27797 6974 28323 6976
rect 27797 6971 27863 6974
rect 28257 6971 28323 6974
rect 0 6898 800 6928
rect 3509 6898 3575 6901
rect 0 6896 3575 6898
rect 0 6840 3514 6896
rect 3570 6840 3575 6896
rect 0 6838 3575 6840
rect 0 6808 800 6838
rect 3509 6835 3575 6838
rect 30649 6898 30715 6901
rect 36629 6898 36695 6901
rect 30649 6896 36695 6898
rect 30649 6840 30654 6896
rect 30710 6840 36634 6896
rect 36690 6840 36695 6896
rect 30649 6838 36695 6840
rect 30649 6835 30715 6838
rect 36629 6835 36695 6838
rect 19568 6560 19888 6561
rect 0 6490 800 6520
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 1393 6490 1459 6493
rect 0 6488 1459 6490
rect 0 6432 1398 6488
rect 1454 6432 1459 6488
rect 0 6430 1459 6432
rect 0 6400 800 6430
rect 1393 6427 1459 6430
rect 48773 6354 48839 6357
rect 49785 6354 49851 6357
rect 52177 6354 52243 6357
rect 48773 6352 52243 6354
rect 48773 6296 48778 6352
rect 48834 6296 49790 6352
rect 49846 6296 52182 6352
rect 52238 6296 52243 6352
rect 48773 6294 52243 6296
rect 48773 6291 48839 6294
rect 49785 6291 49851 6294
rect 52177 6291 52243 6294
rect 31569 6218 31635 6221
rect 36353 6218 36419 6221
rect 31569 6216 36419 6218
rect 31569 6160 31574 6216
rect 31630 6160 36358 6216
rect 36414 6160 36419 6216
rect 31569 6158 36419 6160
rect 31569 6155 31635 6158
rect 36353 6155 36419 6158
rect 0 6082 800 6112
rect 1577 6082 1643 6085
rect 0 6080 1643 6082
rect 0 6024 1582 6080
rect 1638 6024 1643 6080
rect 0 6022 1643 6024
rect 0 5992 800 6022
rect 1577 6019 1643 6022
rect 32397 6082 32463 6085
rect 33133 6082 33199 6085
rect 32397 6080 33199 6082
rect 32397 6024 32402 6080
rect 32458 6024 33138 6080
rect 33194 6024 33199 6080
rect 32397 6022 33199 6024
rect 32397 6019 32463 6022
rect 33133 6019 33199 6022
rect 39665 6082 39731 6085
rect 42517 6082 42583 6085
rect 39665 6080 42583 6082
rect 39665 6024 39670 6080
rect 39726 6024 42522 6080
rect 42578 6024 42583 6080
rect 39665 6022 42583 6024
rect 39665 6019 39731 6022
rect 42517 6019 42583 6022
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 32765 5946 32831 5949
rect 33041 5946 33107 5949
rect 32765 5944 33107 5946
rect 32765 5888 32770 5944
rect 32826 5888 33046 5944
rect 33102 5888 33107 5944
rect 32765 5886 33107 5888
rect 32765 5883 32831 5886
rect 33041 5883 33107 5886
rect 32489 5810 32555 5813
rect 33041 5810 33107 5813
rect 32489 5808 33107 5810
rect 32489 5752 32494 5808
rect 32550 5752 33046 5808
rect 33102 5752 33107 5808
rect 32489 5750 33107 5752
rect 32489 5747 32555 5750
rect 33041 5747 33107 5750
rect 0 5674 800 5704
rect 1853 5674 1919 5677
rect 0 5672 1919 5674
rect 0 5616 1858 5672
rect 1914 5616 1919 5672
rect 0 5614 1919 5616
rect 0 5584 800 5614
rect 1853 5611 1919 5614
rect 19333 5674 19399 5677
rect 22645 5674 22711 5677
rect 19333 5672 22711 5674
rect 19333 5616 19338 5672
rect 19394 5616 22650 5672
rect 22706 5616 22711 5672
rect 19333 5614 22711 5616
rect 19333 5611 19399 5614
rect 22645 5611 22711 5614
rect 32489 5538 32555 5541
rect 33317 5538 33383 5541
rect 32489 5536 33383 5538
rect 32489 5480 32494 5536
rect 32550 5480 33322 5536
rect 33378 5480 33383 5536
rect 32489 5478 33383 5480
rect 32489 5475 32555 5478
rect 33317 5475 33383 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 0 5176 800 5296
rect 32121 5266 32187 5269
rect 33593 5266 33659 5269
rect 32121 5264 33659 5266
rect 32121 5208 32126 5264
rect 32182 5208 33598 5264
rect 33654 5208 33659 5264
rect 32121 5206 33659 5208
rect 32121 5203 32187 5206
rect 33593 5203 33659 5206
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 0 4722 800 4752
rect 3785 4722 3851 4725
rect 0 4720 3851 4722
rect 0 4664 3790 4720
rect 3846 4664 3851 4720
rect 0 4662 3851 4664
rect 0 4632 800 4662
rect 3785 4659 3851 4662
rect 35617 4722 35683 4725
rect 38469 4722 38535 4725
rect 35617 4720 38535 4722
rect 35617 4664 35622 4720
rect 35678 4664 38474 4720
rect 38530 4664 38535 4720
rect 35617 4662 38535 4664
rect 35617 4659 35683 4662
rect 38469 4659 38535 4662
rect 32121 4586 32187 4589
rect 36537 4586 36603 4589
rect 32121 4584 36603 4586
rect 32121 4528 32126 4584
rect 32182 4528 36542 4584
rect 36598 4528 36603 4584
rect 32121 4526 36603 4528
rect 32121 4523 32187 4526
rect 36537 4523 36603 4526
rect 2681 4450 2747 4453
rect 8661 4450 8727 4453
rect 2681 4448 8727 4450
rect 2681 4392 2686 4448
rect 2742 4392 8666 4448
rect 8722 4392 8727 4448
rect 2681 4390 8727 4392
rect 2681 4387 2747 4390
rect 8661 4387 8727 4390
rect 32489 4450 32555 4453
rect 38285 4450 38351 4453
rect 32489 4448 38351 4450
rect 32489 4392 32494 4448
rect 32550 4392 38290 4448
rect 38346 4392 38351 4448
rect 32489 4390 38351 4392
rect 32489 4387 32555 4390
rect 38285 4387 38351 4390
rect 19568 4384 19888 4385
rect 0 4314 800 4344
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 2865 4314 2931 4317
rect 0 4312 2931 4314
rect 0 4256 2870 4312
rect 2926 4256 2931 4312
rect 0 4254 2931 4256
rect 0 4224 800 4254
rect 2865 4251 2931 4254
rect 34697 4314 34763 4317
rect 36905 4314 36971 4317
rect 34697 4312 36971 4314
rect 34697 4256 34702 4312
rect 34758 4256 36910 4312
rect 36966 4256 36971 4312
rect 34697 4254 36971 4256
rect 34697 4251 34763 4254
rect 36905 4251 36971 4254
rect 38285 4314 38351 4317
rect 42701 4314 42767 4317
rect 44909 4314 44975 4317
rect 38285 4312 44975 4314
rect 38285 4256 38290 4312
rect 38346 4256 42706 4312
rect 42762 4256 44914 4312
rect 44970 4256 44975 4312
rect 38285 4254 44975 4256
rect 38285 4251 38351 4254
rect 42701 4251 42767 4254
rect 44909 4251 44975 4254
rect 13905 4178 13971 4181
rect 28441 4178 28507 4181
rect 13905 4176 28507 4178
rect 13905 4120 13910 4176
rect 13966 4120 28446 4176
rect 28502 4120 28507 4176
rect 13905 4118 28507 4120
rect 13905 4115 13971 4118
rect 28441 4115 28507 4118
rect 33317 4178 33383 4181
rect 36077 4178 36143 4181
rect 33317 4176 36143 4178
rect 33317 4120 33322 4176
rect 33378 4120 36082 4176
rect 36138 4120 36143 4176
rect 33317 4118 36143 4120
rect 33317 4115 33383 4118
rect 36077 4115 36143 4118
rect 34513 4042 34579 4045
rect 37273 4042 37339 4045
rect 34513 4040 37339 4042
rect 34513 3984 34518 4040
rect 34574 3984 37278 4040
rect 37334 3984 37339 4040
rect 34513 3982 37339 3984
rect 34513 3979 34579 3982
rect 37273 3979 37339 3982
rect 0 3906 800 3936
rect 1853 3906 1919 3909
rect 0 3904 1919 3906
rect 0 3848 1858 3904
rect 1914 3848 1919 3904
rect 0 3846 1919 3848
rect 0 3816 800 3846
rect 1853 3843 1919 3846
rect 18781 3906 18847 3909
rect 19517 3906 19583 3909
rect 18781 3904 19583 3906
rect 18781 3848 18786 3904
rect 18842 3848 19522 3904
rect 19578 3848 19583 3904
rect 18781 3846 19583 3848
rect 18781 3843 18847 3846
rect 19517 3843 19583 3846
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 33041 3770 33107 3773
rect 34053 3770 34119 3773
rect 33041 3768 34119 3770
rect 33041 3712 33046 3768
rect 33102 3712 34058 3768
rect 34114 3712 34119 3768
rect 33041 3710 34119 3712
rect 33041 3707 33107 3710
rect 34053 3707 34119 3710
rect 21909 3634 21975 3637
rect 25405 3634 25471 3637
rect 21909 3632 25471 3634
rect 21909 3576 21914 3632
rect 21970 3576 25410 3632
rect 25466 3576 25471 3632
rect 21909 3574 25471 3576
rect 21909 3571 21975 3574
rect 25405 3571 25471 3574
rect 31109 3634 31175 3637
rect 38377 3634 38443 3637
rect 31109 3632 38443 3634
rect 31109 3576 31114 3632
rect 31170 3576 38382 3632
rect 38438 3576 38443 3632
rect 31109 3574 38443 3576
rect 31109 3571 31175 3574
rect 38377 3571 38443 3574
rect 0 3408 800 3528
rect 15561 3498 15627 3501
rect 16481 3498 16547 3501
rect 15561 3496 16547 3498
rect 15561 3440 15566 3496
rect 15622 3440 16486 3496
rect 16542 3440 16547 3496
rect 15561 3438 16547 3440
rect 15561 3435 15627 3438
rect 16481 3435 16547 3438
rect 31293 3498 31359 3501
rect 36353 3498 36419 3501
rect 31293 3496 36419 3498
rect 31293 3440 31298 3496
rect 31354 3440 36358 3496
rect 36414 3440 36419 3496
rect 31293 3438 36419 3440
rect 31293 3435 31359 3438
rect 36353 3435 36419 3438
rect 14457 3362 14523 3365
rect 17401 3362 17467 3365
rect 14457 3360 17467 3362
rect 14457 3304 14462 3360
rect 14518 3304 17406 3360
rect 17462 3304 17467 3360
rect 14457 3302 17467 3304
rect 14457 3299 14523 3302
rect 17401 3299 17467 3302
rect 33317 3362 33383 3365
rect 34329 3362 34395 3365
rect 33317 3360 34395 3362
rect 33317 3304 33322 3360
rect 33378 3304 34334 3360
rect 34390 3304 34395 3360
rect 33317 3302 34395 3304
rect 33317 3299 33383 3302
rect 34329 3299 34395 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 13445 3226 13511 3229
rect 15009 3226 15075 3229
rect 13445 3224 15075 3226
rect 13445 3168 13450 3224
rect 13506 3168 15014 3224
rect 15070 3168 15075 3224
rect 13445 3166 15075 3168
rect 13445 3163 13511 3166
rect 15009 3163 15075 3166
rect 0 3090 800 3120
rect 4061 3090 4127 3093
rect 0 3088 4127 3090
rect 0 3032 4066 3088
rect 4122 3032 4127 3088
rect 0 3030 4127 3032
rect 0 3000 800 3030
rect 4061 3027 4127 3030
rect 32121 3090 32187 3093
rect 34329 3090 34395 3093
rect 34605 3090 34671 3093
rect 32121 3088 34671 3090
rect 32121 3032 32126 3088
rect 32182 3032 34334 3088
rect 34390 3032 34610 3088
rect 34666 3032 34671 3088
rect 32121 3030 34671 3032
rect 32121 3027 32187 3030
rect 34329 3027 34395 3030
rect 34605 3027 34671 3030
rect 14733 2954 14799 2957
rect 18045 2954 18111 2957
rect 14733 2952 18111 2954
rect 14733 2896 14738 2952
rect 14794 2896 18050 2952
rect 18106 2896 18111 2952
rect 14733 2894 18111 2896
rect 14733 2891 14799 2894
rect 18045 2891 18111 2894
rect 34329 2954 34395 2957
rect 35525 2954 35591 2957
rect 34329 2952 35591 2954
rect 34329 2896 34334 2952
rect 34390 2896 35530 2952
rect 35586 2896 35591 2952
rect 34329 2894 35591 2896
rect 34329 2891 34395 2894
rect 35525 2891 35591 2894
rect 16113 2818 16179 2821
rect 20069 2818 20135 2821
rect 16113 2816 20135 2818
rect 16113 2760 16118 2816
rect 16174 2760 20074 2816
rect 20130 2760 20135 2816
rect 16113 2758 20135 2760
rect 16113 2755 16179 2758
rect 20069 2755 20135 2758
rect 4208 2752 4528 2753
rect 0 2682 800 2712
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 3049 2682 3115 2685
rect 0 2680 3115 2682
rect 0 2624 3054 2680
rect 3110 2624 3115 2680
rect 0 2622 3115 2624
rect 0 2592 800 2622
rect 3049 2619 3115 2622
rect 32121 2546 32187 2549
rect 35065 2546 35131 2549
rect 32121 2544 35131 2546
rect 32121 2488 32126 2544
rect 32182 2488 35070 2544
rect 35126 2488 35131 2544
rect 32121 2486 35131 2488
rect 32121 2483 32187 2486
rect 35065 2483 35131 2486
rect 31937 2410 32003 2413
rect 35157 2410 35223 2413
rect 31937 2408 35223 2410
rect 31937 2352 31942 2408
rect 31998 2352 35162 2408
rect 35218 2352 35223 2408
rect 31937 2350 35223 2352
rect 31937 2347 32003 2350
rect 35157 2347 35223 2350
rect 0 2274 800 2304
rect 4061 2274 4127 2277
rect 0 2272 4127 2274
rect 0 2216 4066 2272
rect 4122 2216 4127 2272
rect 0 2214 4127 2216
rect 0 2184 800 2214
rect 4061 2211 4127 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
rect 32765 2138 32831 2141
rect 35893 2138 35959 2141
rect 32765 2136 35959 2138
rect 32765 2080 32770 2136
rect 32826 2080 35898 2136
rect 35954 2080 35959 2136
rect 32765 2078 35959 2080
rect 32765 2075 32831 2078
rect 35893 2075 35959 2078
rect 0 1866 800 1896
rect 1393 1866 1459 1869
rect 0 1864 1459 1866
rect 0 1808 1398 1864
rect 1454 1808 1459 1864
rect 0 1806 1459 1808
rect 0 1776 800 1806
rect 1393 1803 1459 1806
rect 0 1458 800 1488
rect 2957 1458 3023 1461
rect 0 1456 3023 1458
rect 0 1400 2962 1456
rect 3018 1400 3023 1456
rect 0 1398 3023 1400
rect 0 1368 800 1398
rect 2957 1395 3023 1398
rect 0 1050 800 1080
rect 3141 1050 3207 1053
rect 0 1048 3207 1050
rect 0 992 3146 1048
rect 3202 992 3207 1048
rect 0 990 3207 992
rect 0 960 800 990
rect 3141 987 3207 990
rect 0 642 800 672
rect 1485 642 1551 645
rect 0 640 1551 642
rect 0 584 1490 640
rect 1546 584 1551 640
rect 0 582 1551 584
rect 0 552 800 582
rect 1485 579 1551 582
rect 0 234 800 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 800 174
rect 2773 171 2839 174
<< via3 >>
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 39744 4528 39760
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 39200 19888 39760
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 39744 35248 39760
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 39200 50608 39760
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__fill_1  FILLER_0_3 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76
timestamp 1644511149
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_123
timestamp 1644511149
transform 1 0 12420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_127
timestamp 1644511149
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1644511149
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1644511149
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_155
timestamp 1644511149
transform 1 0 15364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1644511149
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1644511149
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_183
timestamp 1644511149
transform 1 0 17940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1644511149
transform 1 0 18308 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_214
timestamp 1644511149
transform 1 0 20792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1644511149
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_229
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1644511149
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1644511149
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_285
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_313
timestamp 1644511149
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1644511149
transform 1 0 30544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1644511149
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1644511149
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1644511149
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1644511149
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_375
timestamp 1644511149
transform 1 0 35604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_387
timestamp 1644511149
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1644511149
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1644511149
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_437
timestamp 1644511149
transform 1 0 41308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1644511149
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1644511149
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1644511149
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_485
timestamp 1644511149
transform 1 0 45724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_493
timestamp 1644511149
transform 1 0 46460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1644511149
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_509
timestamp 1644511149
transform 1 0 47932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_514
timestamp 1644511149
transform 1 0 48392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 1644511149
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1644511149
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1644511149
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_553
timestamp 1644511149
transform 1 0 51980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1644511149
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_567
timestamp 1644511149
transform 1 0 53268 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_580
timestamp 1644511149
transform 1 0 54464 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_595
timestamp 1644511149
transform 1 0 55844 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_603
timestamp 1644511149
transform 1 0 56580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_611
timestamp 1644511149
transform 1 0 57316 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1644511149
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1644511149
transform 1 0 58236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1644511149
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_25
timestamp 1644511149
transform 1 0 3404 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_31
timestamp 1644511149
transform 1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1644511149
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_63
timestamp 1644511149
transform 1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1644511149
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 1644511149
transform 1 0 8004 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_79
timestamp 1644511149
transform 1 0 8372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_86
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_116
timestamp 1644511149
transform 1 0 11776 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_124
timestamp 1644511149
transform 1 0 12512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_128
timestamp 1644511149
transform 1 0 12880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1644511149
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_143
timestamp 1644511149
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_155
timestamp 1644511149
transform 1 0 15364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1644511149
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1644511149
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_185
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1644511149
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1644511149
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_269
timestamp 1644511149
transform 1 0 25852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1644511149
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_301 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_313
timestamp 1644511149
transform 1 0 29900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_353
timestamp 1644511149
transform 1 0 33580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp 1644511149
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_411
timestamp 1644511149
transform 1 0 38916 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_419
timestamp 1644511149
transform 1 0 39652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_437
timestamp 1644511149
transform 1 0 41308 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_445
timestamp 1644511149
transform 1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_456
timestamp 1644511149
transform 1 0 43056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_460
timestamp 1644511149
transform 1 0 43424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_477
timestamp 1644511149
transform 1 0 44988 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_499
timestamp 1644511149
transform 1 0 47012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_509
timestamp 1644511149
transform 1 0 47932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1644511149
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_529
timestamp 1644511149
transform 1 0 49772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_535
timestamp 1644511149
transform 1 0 50324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_551
timestamp 1644511149
transform 1 0 51796 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1644511149
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_567
timestamp 1644511149
transform 1 0 53268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_583
timestamp 1644511149
transform 1 0 54740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_599
timestamp 1644511149
transform 1 0 56212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_605
timestamp 1644511149
transform 1 0 56764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_612
timestamp 1644511149
transform 1 0 57408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_621
timestamp 1644511149
transform 1 0 58236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1644511149
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1644511149
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_103
timestamp 1644511149
transform 1 0 10580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_112
timestamp 1644511149
transform 1 0 11408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_158
timestamp 1644511149
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_170
timestamp 1644511149
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_212
timestamp 1644511149
transform 1 0 20608 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_269
timestamp 1644511149
transform 1 0 25852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_296
timestamp 1644511149
transform 1 0 28336 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_317
timestamp 1644511149
transform 1 0 30268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp 1644511149
transform 1 0 30728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_331
timestamp 1644511149
transform 1 0 31556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_343
timestamp 1644511149
transform 1 0 32660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_385
timestamp 1644511149
transform 1 0 36524 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_400
timestamp 1644511149
transform 1 0 37904 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_408
timestamp 1644511149
transform 1 0 38640 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_426
timestamp 1644511149
transform 1 0 40296 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_442
timestamp 1644511149
transform 1 0 41768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_462
timestamp 1644511149
transform 1 0 43608 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1644511149
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_509
timestamp 1644511149
transform 1 0 47932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_521
timestamp 1644511149
transform 1 0 49036 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_529
timestamp 1644511149
transform 1 0 49772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_613
timestamp 1644511149
transform 1 0 57500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1644511149
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_34
timestamp 1644511149
transform 1 0 4232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_41
timestamp 1644511149
transform 1 0 4876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1644511149
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_72
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_101
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1644511149
transform 1 0 12420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1644511149
transform 1 0 13524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1644511149
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_179
timestamp 1644511149
transform 1 0 17572 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_185
timestamp 1644511149
transform 1 0 18124 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_189
timestamp 1644511149
transform 1 0 18492 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_212
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_240
timestamp 1644511149
transform 1 0 23184 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_252
timestamp 1644511149
transform 1 0 24288 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_264
timestamp 1644511149
transform 1 0 25392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_311
timestamp 1644511149
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_323
timestamp 1644511149
transform 1 0 30820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_372
timestamp 1644511149
transform 1 0 35328 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_384
timestamp 1644511149
transform 1 0 36432 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_414
timestamp 1644511149
transform 1 0 39192 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_420
timestamp 1644511149
transform 1 0 39744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_424
timestamp 1644511149
transform 1 0 40112 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_440
timestamp 1644511149
transform 1 0 41584 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_456
timestamp 1644511149
transform 1 0 43056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_465
timestamp 1644511149
transform 1 0 43884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_477
timestamp 1644511149
transform 1 0 44988 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_494
timestamp 1644511149
transform 1 0 46552 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1644511149
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1644511149
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_32
timestamp 1644511149
transform 1 0 4048 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_48
timestamp 1644511149
transform 1 0 5520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_55
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1644511149
transform 1 0 6900 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_71
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_101
timestamp 1644511149
transform 1 0 10396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_113
timestamp 1644511149
transform 1 0 11500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_119
timestamp 1644511149
transform 1 0 12052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 1644511149
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_157
timestamp 1644511149
transform 1 0 15548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_171
timestamp 1644511149
transform 1 0 16836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_183
timestamp 1644511149
transform 1 0 17940 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_204
timestamp 1644511149
transform 1 0 19872 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_211
timestamp 1644511149
transform 1 0 20516 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_226
timestamp 1644511149
transform 1 0 21896 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_238
timestamp 1644511149
transform 1 0 23000 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1644511149
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_259
timestamp 1644511149
transform 1 0 24932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_269
timestamp 1644511149
transform 1 0 25852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_273
timestamp 1644511149
transform 1 0 26220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_279
timestamp 1644511149
transform 1 0 26772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_288
timestamp 1644511149
transform 1 0 27600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_300
timestamp 1644511149
transform 1 0 28704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_343
timestamp 1644511149
transform 1 0 32660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp 1644511149
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_373
timestamp 1644511149
transform 1 0 35420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_383
timestamp 1644511149
transform 1 0 36340 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_391
timestamp 1644511149
transform 1 0 37076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_399
timestamp 1644511149
transform 1 0 37812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_406
timestamp 1644511149
transform 1 0 38456 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_418
timestamp 1644511149
transform 1 0 39560 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_452
timestamp 1644511149
transform 1 0 42688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_462
timestamp 1644511149
transform 1 0 43608 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_474
timestamp 1644511149
transform 1 0 44712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_485
timestamp 1644511149
transform 1 0 45724 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_494
timestamp 1644511149
transform 1 0 46552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_504
timestamp 1644511149
transform 1 0 47472 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_528
timestamp 1644511149
transform 1 0 49680 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1644511149
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_21
timestamp 1644511149
transform 1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1644511149
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_35
timestamp 1644511149
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_42
timestamp 1644511149
transform 1 0 4968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1644511149
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_65
timestamp 1644511149
transform 1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_84
timestamp 1644511149
transform 1 0 8832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_96
timestamp 1644511149
transform 1 0 9936 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_104
timestamp 1644511149
transform 1 0 10672 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1644511149
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_145
timestamp 1644511149
transform 1 0 14444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_153
timestamp 1644511149
transform 1 0 15180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1644511149
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_187
timestamp 1644511149
transform 1 0 18308 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1644511149
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_200
timestamp 1644511149
transform 1 0 19504 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_212
timestamp 1644511149
transform 1 0 20608 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1644511149
transform 1 0 22448 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_244
timestamp 1644511149
transform 1 0 23552 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_256
timestamp 1644511149
transform 1 0 24656 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_264
timestamp 1644511149
transform 1 0 25392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1644511149
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_287
timestamp 1644511149
transform 1 0 27508 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_294
timestamp 1644511149
transform 1 0 28152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_298
timestamp 1644511149
transform 1 0 28520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_323
timestamp 1644511149
transform 1 0 30820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1644511149
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_346
timestamp 1644511149
transform 1 0 32936 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_358
timestamp 1644511149
transform 1 0 34040 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_364
timestamp 1644511149
transform 1 0 34592 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_381
timestamp 1644511149
transform 1 0 36156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1644511149
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1644511149
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_411
timestamp 1644511149
transform 1 0 38916 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_423
timestamp 1644511149
transform 1 0 40020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_431
timestamp 1644511149
transform 1 0 40756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_443
timestamp 1644511149
transform 1 0 41860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_457
timestamp 1644511149
transform 1 0 43148 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_469
timestamp 1644511149
transform 1 0 44252 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_477
timestamp 1644511149
transform 1 0 44988 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_484
timestamp 1644511149
transform 1 0 45632 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_494
timestamp 1644511149
transform 1 0 46552 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1644511149
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1644511149
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_543
timestamp 1644511149
transform 1 0 51060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_555
timestamp 1644511149
transform 1 0 52164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_48
timestamp 1644511149
transform 1 0 5520 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_60
timestamp 1644511149
transform 1 0 6624 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_72
timestamp 1644511149
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1644511149
transform 1 0 9200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_92
timestamp 1644511149
transform 1 0 9568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1644511149
transform 1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_122
timestamp 1644511149
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1644511149
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_160
timestamp 1644511149
transform 1 0 15824 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_172
timestamp 1644511149
transform 1 0 16928 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1644511149
transform 1 0 18032 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_224
timestamp 1644511149
transform 1 0 21712 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_238
timestamp 1644511149
transform 1 0 23000 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1644511149
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_259
timestamp 1644511149
transform 1 0 24932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_268
timestamp 1644511149
transform 1 0 25760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_280
timestamp 1644511149
transform 1 0 26864 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_292
timestamp 1644511149
transform 1 0 27968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1644511149
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_314
timestamp 1644511149
transform 1 0 29992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_326
timestamp 1644511149
transform 1 0 31096 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_338
timestamp 1644511149
transform 1 0 32200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_346
timestamp 1644511149
transform 1 0 32936 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_358
timestamp 1644511149
transform 1 0 34040 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_373
timestamp 1644511149
transform 1 0 35420 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_379
timestamp 1644511149
transform 1 0 35972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_387
timestamp 1644511149
transform 1 0 36708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_399
timestamp 1644511149
transform 1 0 37812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_406
timestamp 1644511149
transform 1 0 38456 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 1644511149
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_437
timestamp 1644511149
transform 1 0 41308 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_449
timestamp 1644511149
transform 1 0 42412 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_461
timestamp 1644511149
transform 1 0 43516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_473
timestamp 1644511149
transform 1 0 44620 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_493
timestamp 1644511149
transform 1 0 46460 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_505
timestamp 1644511149
transform 1 0 47564 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_517
timestamp 1644511149
transform 1 0 48668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_529
timestamp 1644511149
transform 1 0 49772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_560
timestamp 1644511149
transform 1 0 52624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_580
timestamp 1644511149
transform 1 0 54464 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_7
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_20
timestamp 1644511149
transform 1 0 2944 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_32
timestamp 1644511149
transform 1 0 4048 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 1644511149
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1644511149
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_73
timestamp 1644511149
transform 1 0 7820 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_88
timestamp 1644511149
transform 1 0 9200 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_100
timestamp 1644511149
transform 1 0 10304 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_129
timestamp 1644511149
transform 1 0 12972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_146
timestamp 1644511149
transform 1 0 14536 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_152
timestamp 1644511149
transform 1 0 15088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1644511149
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_176
timestamp 1644511149
transform 1 0 17296 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1644511149
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_202
timestamp 1644511149
transform 1 0 19688 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_214
timestamp 1644511149
transform 1 0 20792 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1644511149
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_235
timestamp 1644511149
transform 1 0 22724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_247
timestamp 1644511149
transform 1 0 23828 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_259
timestamp 1644511149
transform 1 0 24932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_271
timestamp 1644511149
transform 1 0 26036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_313
timestamp 1644511149
transform 1 0 29900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_325
timestamp 1644511149
transform 1 0 31004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp 1644511149
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_353
timestamp 1644511149
transform 1 0 33580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_365
timestamp 1644511149
transform 1 0 34684 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_377
timestamp 1644511149
transform 1 0 35788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_381
timestamp 1644511149
transform 1 0 36156 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_387
timestamp 1644511149
transform 1 0 36708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_426
timestamp 1644511149
transform 1 0 40296 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_438
timestamp 1644511149
transform 1 0 41400 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_446
timestamp 1644511149
transform 1 0 42136 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_458
timestamp 1644511149
transform 1 0 43240 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_489
timestamp 1644511149
transform 1 0 46092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1644511149
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_523
timestamp 1644511149
transform 1 0 49220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_534
timestamp 1644511149
transform 1 0 50232 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_546
timestamp 1644511149
transform 1 0 51336 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_558
timestamp 1644511149
transform 1 0 52440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_568
timestamp 1644511149
transform 1 0 53360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_580
timestamp 1644511149
transform 1 0 54464 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_592
timestamp 1644511149
transform 1 0 55568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_604
timestamp 1644511149
transform 1 0 56672 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_13
timestamp 1644511149
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1644511149
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_49
timestamp 1644511149
transform 1 0 5612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_58
timestamp 1644511149
transform 1 0 6440 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_70
timestamp 1644511149
transform 1 0 7544 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1644511149
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_95
timestamp 1644511149
transform 1 0 9844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_107
timestamp 1644511149
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_119
timestamp 1644511149
transform 1 0 12052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_131
timestamp 1644511149
transform 1 0 13156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_147
timestamp 1644511149
transform 1 0 14628 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_155
timestamp 1644511149
transform 1 0 15364 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_168
timestamp 1644511149
transform 1 0 16560 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_179
timestamp 1644511149
transform 1 0 17572 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_191
timestamp 1644511149
transform 1 0 18676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_203
timestamp 1644511149
transform 1 0 19780 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1644511149
transform 1 0 20884 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_227
timestamp 1644511149
transform 1 0 21988 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp 1644511149
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_261
timestamp 1644511149
transform 1 0 25116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_273
timestamp 1644511149
transform 1 0 26220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_285
timestamp 1644511149
transform 1 0 27324 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_295
timestamp 1644511149
transform 1 0 28244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_317
timestamp 1644511149
transform 1 0 30268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_323
timestamp 1644511149
transform 1 0 30820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_335
timestamp 1644511149
transform 1 0 31924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_346
timestamp 1644511149
transform 1 0 32936 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_358
timestamp 1644511149
transform 1 0 34040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_383
timestamp 1644511149
transform 1 0 36340 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_396
timestamp 1644511149
transform 1 0 37536 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_408
timestamp 1644511149
transform 1 0 38640 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_440
timestamp 1644511149
transform 1 0 41584 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_452
timestamp 1644511149
transform 1 0 42688 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_464
timestamp 1644511149
transform 1 0 43792 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_493
timestamp 1644511149
transform 1 0 46460 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_499
timestamp 1644511149
transform 1 0 47012 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_516
timestamp 1644511149
transform 1 0 48576 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_528
timestamp 1644511149
transform 1 0 49680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_564
timestamp 1644511149
transform 1 0 52992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_576
timestamp 1644511149
transform 1 0 54096 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_20
timestamp 1644511149
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_79
timestamp 1644511149
transform 1 0 8372 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_89
timestamp 1644511149
transform 1 0 9292 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_102
timestamp 1644511149
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1644511149
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_118
timestamp 1644511149
transform 1 0 11960 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_124
timestamp 1644511149
transform 1 0 12512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_131
timestamp 1644511149
transform 1 0 13156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_143
timestamp 1644511149
transform 1 0 14260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_151
timestamp 1644511149
transform 1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1644511149
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_176
timestamp 1644511149
transform 1 0 17296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_188
timestamp 1644511149
transform 1 0 18400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_196
timestamp 1644511149
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_202
timestamp 1644511149
transform 1 0 19688 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_206
timestamp 1644511149
transform 1 0 20056 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_213
timestamp 1644511149
transform 1 0 20700 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1644511149
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_233
timestamp 1644511149
transform 1 0 22540 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_241
timestamp 1644511149
transform 1 0 23276 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_255
timestamp 1644511149
transform 1 0 24564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_263
timestamp 1644511149
transform 1 0 25300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_271
timestamp 1644511149
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_289
timestamp 1644511149
transform 1 0 27692 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_296
timestamp 1644511149
transform 1 0 28336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_313
timestamp 1644511149
transform 1 0 29900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_319
timestamp 1644511149
transform 1 0 30452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_327
timestamp 1644511149
transform 1 0 31188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_343
timestamp 1644511149
transform 1 0 32660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_355
timestamp 1644511149
transform 1 0 33764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_376
timestamp 1644511149
transform 1 0 35696 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1644511149
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_397
timestamp 1644511149
transform 1 0 37628 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_415
timestamp 1644511149
transform 1 0 39284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_427
timestamp 1644511149
transform 1 0 40388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_439
timestamp 1644511149
transform 1 0 41492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_457
timestamp 1644511149
transform 1 0 43148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_469
timestamp 1644511149
transform 1 0 44252 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_477
timestamp 1644511149
transform 1 0 44988 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_495
timestamp 1644511149
transform 1 0 46644 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_521
timestamp 1644511149
transform 1 0 49036 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_528
timestamp 1644511149
transform 1 0 49680 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_548
timestamp 1644511149
transform 1 0 51520 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_586
timestamp 1644511149
transform 1 0 55016 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_598
timestamp 1644511149
transform 1 0 56120 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_610
timestamp 1644511149
transform 1 0 57224 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1644511149
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1644511149
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1644511149
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1644511149
transform 1 0 6072 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_66
timestamp 1644511149
transform 1 0 7176 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_74
timestamp 1644511149
transform 1 0 7912 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1644511149
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1644511149
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_104
timestamp 1644511149
transform 1 0 10672 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_112
timestamp 1644511149
transform 1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1644511149
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_146
timestamp 1644511149
transform 1 0 14536 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_161
timestamp 1644511149
transform 1 0 15916 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_173
timestamp 1644511149
transform 1 0 17020 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1644511149
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1644511149
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_203
timestamp 1644511149
transform 1 0 19780 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1644511149
transform 1 0 20884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1644511149
transform 1 0 21988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1644511149
transform 1 0 23092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_259
timestamp 1644511149
transform 1 0 24932 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_268
timestamp 1644511149
transform 1 0 25760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_276
timestamp 1644511149
transform 1 0 26496 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_284
timestamp 1644511149
transform 1 0 27232 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_290
timestamp 1644511149
transform 1 0 27784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1644511149
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_314
timestamp 1644511149
transform 1 0 29992 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_322
timestamp 1644511149
transform 1 0 30728 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_341
timestamp 1644511149
transform 1 0 32476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_349
timestamp 1644511149
transform 1 0 33212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1644511149
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_370
timestamp 1644511149
transform 1 0 35144 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_382
timestamp 1644511149
transform 1 0 36248 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_394
timestamp 1644511149
transform 1 0 37352 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_398
timestamp 1644511149
transform 1 0 37720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_402
timestamp 1644511149
transform 1 0 38088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_410
timestamp 1644511149
transform 1 0 38824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp 1644511149
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_452
timestamp 1644511149
transform 1 0 42688 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_464
timestamp 1644511149
transform 1 0 43792 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_487
timestamp 1644511149
transform 1 0 45908 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_495
timestamp 1644511149
transform 1 0 46644 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_507
timestamp 1644511149
transform 1 0 47748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_519
timestamp 1644511149
transform 1 0 48852 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_565
timestamp 1644511149
transform 1 0 53084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_577
timestamp 1644511149
transform 1 0 54188 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_585
timestamp 1644511149
transform 1 0 54924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_25
timestamp 1644511149
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_37
timestamp 1644511149
transform 1 0 4508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_43
timestamp 1644511149
transform 1 0 5060 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_50
timestamp 1644511149
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_153
timestamp 1644511149
transform 1 0 15180 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1644511149
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_179
timestamp 1644511149
transform 1 0 17572 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_187
timestamp 1644511149
transform 1 0 18308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_233
timestamp 1644511149
transform 1 0 22540 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_245
timestamp 1644511149
transform 1 0 23644 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_253
timestamp 1644511149
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_264
timestamp 1644511149
transform 1 0 25392 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_287
timestamp 1644511149
transform 1 0 27508 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_294
timestamp 1644511149
transform 1 0 28152 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_298
timestamp 1644511149
transform 1 0 28520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_313
timestamp 1644511149
transform 1 0 29900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_326
timestamp 1644511149
transform 1 0 31096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1644511149
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_341
timestamp 1644511149
transform 1 0 32476 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_355
timestamp 1644511149
transform 1 0 33764 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_367
timestamp 1644511149
transform 1 0 34868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_374
timestamp 1644511149
transform 1 0 35512 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1644511149
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_401
timestamp 1644511149
transform 1 0 37996 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_407
timestamp 1644511149
transform 1 0 38548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_413
timestamp 1644511149
transform 1 0 39100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_421
timestamp 1644511149
transform 1 0 39836 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_433
timestamp 1644511149
transform 1 0 40940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_437
timestamp 1644511149
transform 1 0 41308 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_444
timestamp 1644511149
transform 1 0 41952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_457
timestamp 1644511149
transform 1 0 43148 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_469
timestamp 1644511149
transform 1 0 44252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_482
timestamp 1644511149
transform 1 0 45448 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_494
timestamp 1644511149
transform 1 0 46552 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1644511149
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1644511149
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_522
timestamp 1644511149
transform 1 0 49128 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_539
timestamp 1644511149
transform 1 0 50692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_551
timestamp 1644511149
transform 1 0 51796 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_6
timestamp 1644511149
transform 1 0 1656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1644511149
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_90
timestamp 1644511149
transform 1 0 9384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_94
timestamp 1644511149
transform 1 0 9752 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_101
timestamp 1644511149
transform 1 0 10396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_113
timestamp 1644511149
transform 1 0 11500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_125
timestamp 1644511149
transform 1 0 12604 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1644511149
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_147
timestamp 1644511149
transform 1 0 14628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_158
timestamp 1644511149
transform 1 0 15640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_169
timestamp 1644511149
transform 1 0 16652 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_181
timestamp 1644511149
transform 1 0 17756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1644511149
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_203
timestamp 1644511149
transform 1 0 19780 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1644511149
transform 1 0 20884 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_223
timestamp 1644511149
transform 1 0 21620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_229
timestamp 1644511149
transform 1 0 22172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_235
timestamp 1644511149
transform 1 0 22724 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_246
timestamp 1644511149
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_293
timestamp 1644511149
transform 1 0 28060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_300
timestamp 1644511149
transform 1 0 28704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_349
timestamp 1644511149
transform 1 0 33212 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_358
timestamp 1644511149
transform 1 0 34040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_383
timestamp 1644511149
transform 1 0 36340 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_391
timestamp 1644511149
transform 1 0 37076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_405
timestamp 1644511149
transform 1 0 38364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_441
timestamp 1644511149
transform 1 0 41676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_449
timestamp 1644511149
transform 1 0 42412 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_461
timestamp 1644511149
transform 1 0 43516 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_473
timestamp 1644511149
transform 1 0 44620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_485
timestamp 1644511149
transform 1 0 45724 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_494
timestamp 1644511149
transform 1 0 46552 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_506
timestamp 1644511149
transform 1 0 47656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_528
timestamp 1644511149
transform 1 0 49680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_537
timestamp 1644511149
transform 1 0 50508 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_544
timestamp 1644511149
transform 1 0 51152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_564
timestamp 1644511149
transform 1 0 52992 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_576
timestamp 1644511149
transform 1 0 54096 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_7
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_20
timestamp 1644511149
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1644511149
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1644511149
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_74
timestamp 1644511149
transform 1 0 7912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1644511149
transform 1 0 8648 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1644511149
transform 1 0 9752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_100
timestamp 1644511149
transform 1 0 10304 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_121
timestamp 1644511149
transform 1 0 12236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_136
timestamp 1644511149
transform 1 0 13616 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_152
timestamp 1644511149
transform 1 0 15088 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1644511149
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_203
timestamp 1644511149
transform 1 0 19780 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1644511149
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_241
timestamp 1644511149
transform 1 0 23276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_253
timestamp 1644511149
transform 1 0 24380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_266
timestamp 1644511149
transform 1 0 25576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_274
timestamp 1644511149
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_301
timestamp 1644511149
transform 1 0 28796 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_313
timestamp 1644511149
transform 1 0 29900 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_321
timestamp 1644511149
transform 1 0 30636 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1644511149
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_366
timestamp 1644511149
transform 1 0 34776 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_374
timestamp 1644511149
transform 1 0 35512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_379
timestamp 1644511149
transform 1 0 35972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1644511149
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_403
timestamp 1644511149
transform 1 0 38180 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_414
timestamp 1644511149
transform 1 0 39192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_421
timestamp 1644511149
transform 1 0 39836 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_433
timestamp 1644511149
transform 1 0 40940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 1644511149
transform 1 0 42044 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_457
timestamp 1644511149
transform 1 0 43148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_469
timestamp 1644511149
transform 1 0 44252 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_481
timestamp 1644511149
transform 1 0 45356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_500
timestamp 1644511149
transform 1 0 47104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_528
timestamp 1644511149
transform 1 0 49680 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_540
timestamp 1644511149
transform 1 0 50784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_552
timestamp 1644511149
transform 1 0 51888 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1644511149
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_59
timestamp 1644511149
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_74
timestamp 1644511149
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1644511149
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1644511149
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_100
timestamp 1644511149
transform 1 0 10304 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_112
timestamp 1644511149
transform 1 0 11408 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_118
timestamp 1644511149
transform 1 0 11960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1644511149
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_161
timestamp 1644511149
transform 1 0 15916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_169
timestamp 1644511149
transform 1 0 16652 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1644511149
transform 1 0 17480 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1644511149
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_235
timestamp 1644511149
transform 1 0 22724 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp 1644511149
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_285
timestamp 1644511149
transform 1 0 27324 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_302
timestamp 1644511149
transform 1 0 28888 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_340
timestamp 1644511149
transform 1 0 32384 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_352
timestamp 1644511149
transform 1 0 33488 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_384
timestamp 1644511149
transform 1 0 36432 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_393
timestamp 1644511149
transform 1 0 37260 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_400
timestamp 1644511149
transform 1 0 37904 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_408
timestamp 1644511149
transform 1 0 38640 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1644511149
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_452
timestamp 1644511149
transform 1 0 42688 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_464
timestamp 1644511149
transform 1 0 43792 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_485
timestamp 1644511149
transform 1 0 45724 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_493
timestamp 1644511149
transform 1 0 46460 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_511
timestamp 1644511149
transform 1 0 48116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_523
timestamp 1644511149
transform 1 0 49220 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_564
timestamp 1644511149
transform 1 0 52992 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_576
timestamp 1644511149
transform 1 0 54096 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_26
timestamp 1644511149
transform 1 0 3496 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_38
timestamp 1644511149
transform 1 0 4600 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1644511149
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_63
timestamp 1644511149
transform 1 0 6900 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_71
timestamp 1644511149
transform 1 0 7636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_83
timestamp 1644511149
transform 1 0 8740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_87
timestamp 1644511149
transform 1 0 9108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_104
timestamp 1644511149
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp 1644511149
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_140
timestamp 1644511149
transform 1 0 13984 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1644511149
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_156
timestamp 1644511149
transform 1 0 15456 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1644511149
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_176
timestamp 1644511149
transform 1 0 17296 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_184
timestamp 1644511149
transform 1 0 18032 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_201
timestamp 1644511149
transform 1 0 19596 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_213
timestamp 1644511149
transform 1 0 20700 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_229
timestamp 1644511149
transform 1 0 22172 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_235
timestamp 1644511149
transform 1 0 22724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_247
timestamp 1644511149
transform 1 0 23828 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_255
timestamp 1644511149
transform 1 0 24564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_259
timestamp 1644511149
transform 1 0 24932 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_271
timestamp 1644511149
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_289
timestamp 1644511149
transform 1 0 27692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_294
timestamp 1644511149
transform 1 0 28152 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_306
timestamp 1644511149
transform 1 0 29256 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_318
timestamp 1644511149
transform 1 0 30360 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_324
timestamp 1644511149
transform 1 0 30912 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1644511149
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_409
timestamp 1644511149
transform 1 0 38732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_419
timestamp 1644511149
transform 1 0 39652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_432
timestamp 1644511149
transform 1 0 40848 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_444
timestamp 1644511149
transform 1 0 41952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_526
timestamp 1644511149
transform 1 0 49496 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_538
timestamp 1644511149
transform 1 0 50600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_550
timestamp 1644511149
transform 1 0 51704 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_558
timestamp 1644511149
transform 1 0 52440 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1644511149
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1644511149
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_48
timestamp 1644511149
transform 1 0 5520 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_60
timestamp 1644511149
transform 1 0 6624 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_72
timestamp 1644511149
transform 1 0 7728 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1644511149
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_100
timestamp 1644511149
transform 1 0 10304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_112
timestamp 1644511149
transform 1 0 11408 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_124
timestamp 1644511149
transform 1 0 12512 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp 1644511149
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1644511149
transform 1 0 14352 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_156
timestamp 1644511149
transform 1 0 15456 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_164
timestamp 1644511149
transform 1 0 16192 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_175
timestamp 1644511149
transform 1 0 17204 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_186
timestamp 1644511149
transform 1 0 18216 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1644511149
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_217
timestamp 1644511149
transform 1 0 21068 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_223
timestamp 1644511149
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_237
timestamp 1644511149
transform 1 0 22908 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_274
timestamp 1644511149
transform 1 0 26312 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_286
timestamp 1644511149
transform 1 0 27416 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_299
timestamp 1644511149
transform 1 0 28612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_317
timestamp 1644511149
transform 1 0 30268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_329
timestamp 1644511149
transform 1 0 31372 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_341
timestamp 1644511149
transform 1 0 32476 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_353
timestamp 1644511149
transform 1 0 33580 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1644511149
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_372
timestamp 1644511149
transform 1 0 35328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_383
timestamp 1644511149
transform 1 0 36340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_390
timestamp 1644511149
transform 1 0 36984 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_402
timestamp 1644511149
transform 1 0 38088 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_414
timestamp 1644511149
transform 1 0 39192 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_429
timestamp 1644511149
transform 1 0 40572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_435
timestamp 1644511149
transform 1 0 41124 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_447
timestamp 1644511149
transform 1 0 42228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_459
timestamp 1644511149
transform 1 0 43332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_471
timestamp 1644511149
transform 1 0 44436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_505
timestamp 1644511149
transform 1 0 47564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_509
timestamp 1644511149
transform 1 0 47932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_518
timestamp 1644511149
transform 1 0 48760 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_530
timestamp 1644511149
transform 1 0 49864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_550
timestamp 1644511149
transform 1 0 51704 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_562
timestamp 1644511149
transform 1 0 52808 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_574
timestamp 1644511149
transform 1 0 53912 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_586
timestamp 1644511149
transform 1 0 55016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1644511149
transform 1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_20
timestamp 1644511149
transform 1 0 2944 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_47
timestamp 1644511149
transform 1 0 5428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1644511149
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_65
timestamp 1644511149
transform 1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_72
timestamp 1644511149
transform 1 0 7728 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_78
timestamp 1644511149
transform 1 0 8280 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_89
timestamp 1644511149
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1644511149
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1644511149
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1644511149
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_133
timestamp 1644511149
transform 1 0 13340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_145
timestamp 1644511149
transform 1 0 14444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1644511149
transform 1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_189
timestamp 1644511149
transform 1 0 18492 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_198
timestamp 1644511149
transform 1 0 19320 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_210
timestamp 1644511149
transform 1 0 20424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1644511149
transform 1 0 22448 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1644511149
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_253
timestamp 1644511149
transform 1 0 24380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_265
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1644511149
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_300
timestamp 1644511149
transform 1 0 28704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_311
timestamp 1644511149
transform 1 0 29716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_323
timestamp 1644511149
transform 1 0 30820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_345
timestamp 1644511149
transform 1 0 32844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_357
timestamp 1644511149
transform 1 0 33948 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_379
timestamp 1644511149
transform 1 0 35972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_387
timestamp 1644511149
transform 1 0 36708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_455
timestamp 1644511149
transform 1 0 42964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_475
timestamp 1644511149
transform 1 0 44804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_496
timestamp 1644511149
transform 1 0 46736 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_512
timestamp 1644511149
transform 1 0 48208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_523
timestamp 1644511149
transform 1 0 49220 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_535
timestamp 1644511149
transform 1 0 50324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_551
timestamp 1644511149
transform 1 0 51796 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_578
timestamp 1644511149
transform 1 0 54280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_598
timestamp 1644511149
transform 1 0 56120 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_610
timestamp 1644511149
transform 1 0 57224 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1644511149
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1644511149
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_57
timestamp 1644511149
transform 1 0 6348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_63
timestamp 1644511149
transform 1 0 6900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 1644511149
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1644511149
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_95
timestamp 1644511149
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_116
timestamp 1644511149
transform 1 0 11776 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_124
timestamp 1644511149
transform 1 0 12512 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_130
timestamp 1644511149
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1644511149
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_147
timestamp 1644511149
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_158
timestamp 1644511149
transform 1 0 15640 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_167
timestamp 1644511149
transform 1 0 16468 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_185
timestamp 1644511149
transform 1 0 18124 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1644511149
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1644511149
transform 1 0 20884 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_222
timestamp 1644511149
transform 1 0 21528 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_229
timestamp 1644511149
transform 1 0 22172 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1644511149
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1644511149
transform 1 0 24840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_267
timestamp 1644511149
transform 1 0 25668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_287
timestamp 1644511149
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_302
timestamp 1644511149
transform 1 0 28888 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_326
timestamp 1644511149
transform 1 0 31096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_335
timestamp 1644511149
transform 1 0 31924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_347
timestamp 1644511149
transform 1 0 33028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_359
timestamp 1644511149
transform 1 0 34132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_372
timestamp 1644511149
transform 1 0 35328 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_383
timestamp 1644511149
transform 1 0 36340 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_395
timestamp 1644511149
transform 1 0 37444 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_403
timestamp 1644511149
transform 1 0 38180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_412
timestamp 1644511149
transform 1 0 39008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_424
timestamp 1644511149
transform 1 0 40112 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_436
timestamp 1644511149
transform 1 0 41216 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_442
timestamp 1644511149
transform 1 0 41768 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_449
timestamp 1644511149
transform 1 0 42412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_461
timestamp 1644511149
transform 1 0 43516 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_507
timestamp 1644511149
transform 1 0 47748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_517
timestamp 1644511149
transform 1 0 48668 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_529
timestamp 1644511149
transform 1 0 49772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_537
timestamp 1644511149
transform 1 0 50508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_554
timestamp 1644511149
transform 1 0 52072 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_566
timestamp 1644511149
transform 1 0 53176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_578
timestamp 1644511149
transform 1 0 54280 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_586
timestamp 1644511149
transform 1 0 55016 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_593
timestamp 1644511149
transform 1 0 55660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_605
timestamp 1644511149
transform 1 0 56764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_617
timestamp 1644511149
transform 1 0 57868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_13
timestamp 1644511149
transform 1 0 2300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_21
timestamp 1644511149
transform 1 0 3036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1644511149
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_38
timestamp 1644511149
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1644511149
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_65
timestamp 1644511149
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_73
timestamp 1644511149
transform 1 0 7820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1644511149
transform 1 0 8648 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_94
timestamp 1644511149
transform 1 0 9752 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1644511149
transform 1 0 10304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1644511149
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_119
timestamp 1644511149
transform 1 0 12052 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_131
timestamp 1644511149
transform 1 0 13156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_139
timestamp 1644511149
transform 1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_148
timestamp 1644511149
transform 1 0 14720 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1644511149
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_173
timestamp 1644511149
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_190
timestamp 1644511149
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_200
timestamp 1644511149
transform 1 0 19504 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_212
timestamp 1644511149
transform 1 0 20608 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1644511149
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_244
timestamp 1644511149
transform 1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_252
timestamp 1644511149
transform 1 0 24288 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_260
timestamp 1644511149
transform 1 0 25024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_267
timestamp 1644511149
transform 1 0 25668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_326
timestamp 1644511149
transform 1 0 31096 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1644511149
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_354
timestamp 1644511149
transform 1 0 33672 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_366
timestamp 1644511149
transform 1 0 34776 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_372
timestamp 1644511149
transform 1 0 35328 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_379
timestamp 1644511149
transform 1 0 35972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_401
timestamp 1644511149
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_418
timestamp 1644511149
transform 1 0 39560 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_426
timestamp 1644511149
transform 1 0 40296 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_432
timestamp 1644511149
transform 1 0 40848 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_440
timestamp 1644511149
transform 1 0 41584 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 1644511149
transform 1 0 41952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_456
timestamp 1644511149
transform 1 0 43056 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_464
timestamp 1644511149
transform 1 0 43792 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_476
timestamp 1644511149
transform 1 0 44896 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_491
timestamp 1644511149
transform 1 0 46276 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_520
timestamp 1644511149
transform 1 0 48944 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_532
timestamp 1644511149
transform 1 0 50048 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_556
timestamp 1644511149
transform 1 0 52256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_592
timestamp 1644511149
transform 1 0 55568 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_596
timestamp 1644511149
transform 1 0 55936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_600
timestamp 1644511149
transform 1 0 56304 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_612
timestamp 1644511149
transform 1 0 57408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_7
timestamp 1644511149
transform 1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_14
timestamp 1644511149
transform 1 0 2392 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1644511149
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_45
timestamp 1644511149
transform 1 0 5244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_57
timestamp 1644511149
transform 1 0 6348 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_72
timestamp 1644511149
transform 1 0 7728 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1644511149
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_103
timestamp 1644511149
transform 1 0 10580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_111
timestamp 1644511149
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_122
timestamp 1644511149
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1644511149
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_157
timestamp 1644511149
transform 1 0 15548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_169
timestamp 1644511149
transform 1 0 16652 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_181
timestamp 1644511149
transform 1 0 17756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1644511149
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_211
timestamp 1644511149
transform 1 0 20516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_215
timestamp 1644511149
transform 1 0 20884 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_220
timestamp 1644511149
transform 1 0 21344 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_230
timestamp 1644511149
transform 1 0 22264 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_236
timestamp 1644511149
transform 1 0 22816 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_240
timestamp 1644511149
transform 1 0 23184 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1644511149
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_263
timestamp 1644511149
transform 1 0 25300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_267
timestamp 1644511149
transform 1 0 25668 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_273
timestamp 1644511149
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_280
timestamp 1644511149
transform 1 0 26864 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_292
timestamp 1644511149
transform 1 0 27968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_298
timestamp 1644511149
transform 1 0 28520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1644511149
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_317
timestamp 1644511149
transform 1 0 30268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_322
timestamp 1644511149
transform 1 0 30728 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_330
timestamp 1644511149
transform 1 0 31464 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_335
timestamp 1644511149
transform 1 0 31924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_347
timestamp 1644511149
transform 1 0 33028 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_358
timestamp 1644511149
transform 1 0 34040 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_387
timestamp 1644511149
transform 1 0 36708 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_395
timestamp 1644511149
transform 1 0 37444 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_439
timestamp 1644511149
transform 1 0 41492 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_447
timestamp 1644511149
transform 1 0 42228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_456
timestamp 1644511149
transform 1 0 43056 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_468
timestamp 1644511149
transform 1 0 44160 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_485
timestamp 1644511149
transform 1 0 45724 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_504
timestamp 1644511149
transform 1 0 47472 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_512
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_518
timestamp 1644511149
transform 1 0 48760 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_530
timestamp 1644511149
transform 1 0 49864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_539
timestamp 1644511149
transform 1 0 50692 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_547
timestamp 1644511149
transform 1 0 51428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_554
timestamp 1644511149
transform 1 0 52072 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_566
timestamp 1644511149
transform 1 0 53176 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_570
timestamp 1644511149
transform 1 0 53544 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_578
timestamp 1644511149
transform 1 0 54280 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_584
timestamp 1644511149
transform 1 0 54832 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_596
timestamp 1644511149
transform 1 0 55936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_616
timestamp 1644511149
transform 1 0 57776 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_624
timestamp 1644511149
transform 1 0 58512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_7
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_19
timestamp 1644511149
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1644511149
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_43
timestamp 1644511149
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_97
timestamp 1644511149
transform 1 0 10028 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1644511149
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_146
timestamp 1644511149
transform 1 0 14536 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1644511149
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1644511149
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_176
timestamp 1644511149
transform 1 0 17296 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_187
timestamp 1644511149
transform 1 0 18308 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1644511149
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_242
timestamp 1644511149
transform 1 0 23368 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_258
timestamp 1644511149
transform 1 0 24840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_266
timestamp 1644511149
transform 1 0 25576 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1644511149
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_365
timestamp 1644511149
transform 1 0 34684 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_371
timestamp 1644511149
transform 1 0 35236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_376
timestamp 1644511149
transform 1 0 35696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_401
timestamp 1644511149
transform 1 0 37996 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_410
timestamp 1644511149
transform 1 0 38824 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_422
timestamp 1644511149
transform 1 0 39928 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_426
timestamp 1644511149
transform 1 0 40296 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_437
timestamp 1644511149
transform 1 0 41308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1644511149
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_467
timestamp 1644511149
transform 1 0 44068 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_479
timestamp 1644511149
transform 1 0 45172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_483
timestamp 1644511149
transform 1 0 45540 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_489
timestamp 1644511149
transform 1 0 46092 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_501
timestamp 1644511149
transform 1 0 47196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_512
timestamp 1644511149
transform 1 0 48208 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_524
timestamp 1644511149
transform 1 0 49312 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_536
timestamp 1644511149
transform 1 0 50416 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_548
timestamp 1644511149
transform 1 0 51520 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_568
timestamp 1644511149
transform 1 0 53360 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_572
timestamp 1644511149
transform 1 0 53728 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_580
timestamp 1644511149
transform 1 0 54464 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_592
timestamp 1644511149
transform 1 0 55568 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_604
timestamp 1644511149
transform 1 0 56672 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1644511149
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_59
timestamp 1644511149
transform 1 0 6532 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_66
timestamp 1644511149
transform 1 0 7176 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1644511149
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_90
timestamp 1644511149
transform 1 0 9384 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_102
timestamp 1644511149
transform 1 0 10488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_114
timestamp 1644511149
transform 1 0 11592 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_126
timestamp 1644511149
transform 1 0 12696 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1644511149
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_147
timestamp 1644511149
transform 1 0 14628 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_159
timestamp 1644511149
transform 1 0 15732 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_172
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_183
timestamp 1644511149
transform 1 0 17940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_269
timestamp 1644511149
transform 1 0 25852 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_275
timestamp 1644511149
transform 1 0 26404 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_287
timestamp 1644511149
transform 1 0 27508 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_293
timestamp 1644511149
transform 1 0 28060 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1644511149
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_325
timestamp 1644511149
transform 1 0 31004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_337
timestamp 1644511149
transform 1 0 32108 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_349
timestamp 1644511149
transform 1 0 33212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1644511149
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_383
timestamp 1644511149
transform 1 0 36340 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_390
timestamp 1644511149
transform 1 0 36984 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_398
timestamp 1644511149
transform 1 0 37720 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_416
timestamp 1644511149
transform 1 0 39376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_453
timestamp 1644511149
transform 1 0 42780 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_465
timestamp 1644511149
transform 1 0 43884 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1644511149
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_508
timestamp 1644511149
transform 1 0 47840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_517
timestamp 1644511149
transform 1 0 48668 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_524
timestamp 1644511149
transform 1 0 49312 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_539
timestamp 1644511149
transform 1 0 50692 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_556
timestamp 1644511149
transform 1 0 52256 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_568
timestamp 1644511149
transform 1 0 53360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_580
timestamp 1644511149
transform 1 0 54464 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_593
timestamp 1644511149
transform 1 0 55660 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_605
timestamp 1644511149
transform 1 0 56764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_617
timestamp 1644511149
transform 1 0 57868 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_14
timestamp 1644511149
transform 1 0 2392 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_26
timestamp 1644511149
transform 1 0 3496 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_34
timestamp 1644511149
transform 1 0 4232 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_46
timestamp 1644511149
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1644511149
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_65
timestamp 1644511149
transform 1 0 7084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_75
timestamp 1644511149
transform 1 0 8004 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_87
timestamp 1644511149
transform 1 0 9108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_99
timestamp 1644511149
transform 1 0 10212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_122
timestamp 1644511149
transform 1 0 12328 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1644511149
transform 1 0 13524 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1644511149
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1644511149
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1644511149
transform 1 0 17480 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_201
timestamp 1644511149
transform 1 0 19596 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_213
timestamp 1644511149
transform 1 0 20700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1644511149
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1644511149
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_239
timestamp 1644511149
transform 1 0 23092 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_246
timestamp 1644511149
transform 1 0 23736 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_250
timestamp 1644511149
transform 1 0 24104 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1644511149
transform 1 0 24748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_284
timestamp 1644511149
transform 1 0 27232 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_296
timestamp 1644511149
transform 1 0 28336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_300
timestamp 1644511149
transform 1 0 28704 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_307
timestamp 1644511149
transform 1 0 29348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_318
timestamp 1644511149
transform 1 0 30360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_325
timestamp 1644511149
transform 1 0 31004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1644511149
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_353
timestamp 1644511149
transform 1 0 33580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_365
timestamp 1644511149
transform 1 0 34684 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_377
timestamp 1644511149
transform 1 0 35788 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 1644511149
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_414
timestamp 1644511149
transform 1 0 39192 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_426
timestamp 1644511149
transform 1 0 40296 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_434
timestamp 1644511149
transform 1 0 41032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_478
timestamp 1644511149
transform 1 0 45080 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_490
timestamp 1644511149
transform 1 0 46184 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_502
timestamp 1644511149
transform 1 0 47288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_521
timestamp 1644511149
transform 1 0 49036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_537
timestamp 1644511149
transform 1 0 50508 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_544
timestamp 1644511149
transform 1 0 51152 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_556
timestamp 1644511149
transform 1 0 52256 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_568
timestamp 1644511149
transform 1 0 53360 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_580
timestamp 1644511149
transform 1 0 54464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_591
timestamp 1644511149
transform 1 0 55476 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_595
timestamp 1644511149
transform 1 0 55844 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_612
timestamp 1644511149
transform 1 0 57408 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_14
timestamp 1644511149
transform 1 0 2392 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1644511149
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_48
timestamp 1644511149
transform 1 0 5520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_56
timestamp 1644511149
transform 1 0 6256 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1644511149
transform 1 0 7360 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1644511149
transform 1 0 11224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_118
timestamp 1644511149
transform 1 0 11960 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_130
timestamp 1644511149
transform 1 0 13064 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1644511149
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_161
timestamp 1644511149
transform 1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_173
timestamp 1644511149
transform 1 0 17020 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_184
timestamp 1644511149
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_205
timestamp 1644511149
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_223
timestamp 1644511149
transform 1 0 21620 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_235
timestamp 1644511149
transform 1 0 22724 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_240
timestamp 1644511149
transform 1 0 23184 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_259
timestamp 1644511149
transform 1 0 24932 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_267
timestamp 1644511149
transform 1 0 25668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_287
timestamp 1644511149
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1644511149
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_314
timestamp 1644511149
transform 1 0 29992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_326
timestamp 1644511149
transform 1 0 31096 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_338
timestamp 1644511149
transform 1 0 32200 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_349
timestamp 1644511149
transform 1 0 33212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_361
timestamp 1644511149
transform 1 0 34316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_449
timestamp 1644511149
transform 1 0 42412 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_458
timestamp 1644511149
transform 1 0 43240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_468
timestamp 1644511149
transform 1 0 44160 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_507
timestamp 1644511149
transform 1 0 47748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_511
timestamp 1644511149
transform 1 0 48116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_523
timestamp 1644511149
transform 1 0 49220 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_553
timestamp 1644511149
transform 1 0 51980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_559
timestamp 1644511149
transform 1 0 52532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_570
timestamp 1644511149
transform 1 0 53544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_584
timestamp 1644511149
transform 1 0 54832 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_596
timestamp 1644511149
transform 1 0 55936 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_608
timestamp 1644511149
transform 1 0 57040 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_620
timestamp 1644511149
transform 1 0 58144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_624
timestamp 1644511149
transform 1 0 58512 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_19
timestamp 1644511149
transform 1 0 2852 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_31
timestamp 1644511149
transform 1 0 3956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_38
timestamp 1644511149
transform 1 0 4600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1644511149
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_77
timestamp 1644511149
transform 1 0 8188 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_89
timestamp 1644511149
transform 1 0 9292 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1644511149
transform 1 0 11960 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_157
timestamp 1644511149
transform 1 0 15548 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1644511149
transform 1 0 17572 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_190
timestamp 1644511149
transform 1 0 18584 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_202
timestamp 1644511149
transform 1 0 19688 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_214
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1644511149
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_231
timestamp 1644511149
transform 1 0 22356 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_239
timestamp 1644511149
transform 1 0 23092 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_256
timestamp 1644511149
transform 1 0 24656 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_268
timestamp 1644511149
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_301
timestamp 1644511149
transform 1 0 28796 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_309
timestamp 1644511149
transform 1 0 29532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_318
timestamp 1644511149
transform 1 0 30360 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_330
timestamp 1644511149
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_341
timestamp 1644511149
transform 1 0 32476 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_358
timestamp 1644511149
transform 1 0 34040 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_370
timestamp 1644511149
transform 1 0 35144 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_388
timestamp 1644511149
transform 1 0 36800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_430
timestamp 1644511149
transform 1 0 40664 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_442
timestamp 1644511149
transform 1 0 41768 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_465
timestamp 1644511149
transform 1 0 43884 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_477
timestamp 1644511149
transform 1 0 44988 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_489
timestamp 1644511149
transform 1 0 46092 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_509
timestamp 1644511149
transform 1 0 47932 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_521
timestamp 1644511149
transform 1 0 49036 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_533
timestamp 1644511149
transform 1 0 50140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_545
timestamp 1644511149
transform 1 0 51244 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_551
timestamp 1644511149
transform 1 0 51796 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_565
timestamp 1644511149
transform 1 0 53084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_570
timestamp 1644511149
transform 1 0 53544 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_578
timestamp 1644511149
transform 1 0 54280 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_590
timestamp 1644511149
transform 1 0 55384 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_602
timestamp 1644511149
transform 1 0 56488 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_614
timestamp 1644511149
transform 1 0 57592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1644511149
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_64
timestamp 1644511149
transform 1 0 6992 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_76
timestamp 1644511149
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1644511149
transform 1 0 10764 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_110
timestamp 1644511149
transform 1 0 11224 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_118
timestamp 1644511149
transform 1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1644511149
transform 1 0 14720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_156
timestamp 1644511149
transform 1 0 15456 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1644511149
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_168
timestamp 1644511149
transform 1 0 16560 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_176
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1644511149
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_205
timestamp 1644511149
transform 1 0 19964 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_224
timestamp 1644511149
transform 1 0 21712 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_236
timestamp 1644511149
transform 1 0 22816 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_258
timestamp 1644511149
transform 1 0 24840 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_262
timestamp 1644511149
transform 1 0 25208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_270
timestamp 1644511149
transform 1 0 25944 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_282
timestamp 1644511149
transform 1 0 27048 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_294
timestamp 1644511149
transform 1 0 28152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_369
timestamp 1644511149
transform 1 0 35052 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_373
timestamp 1644511149
transform 1 0 35420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_385
timestamp 1644511149
transform 1 0 36524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_392
timestamp 1644511149
transform 1 0 37168 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_412
timestamp 1644511149
transform 1 0 39008 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_429
timestamp 1644511149
transform 1 0 40572 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_438
timestamp 1644511149
transform 1 0 41400 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_454
timestamp 1644511149
transform 1 0 42872 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_466
timestamp 1644511149
transform 1 0 43976 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_474
timestamp 1644511149
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_481
timestamp 1644511149
transform 1 0 45356 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_490
timestamp 1644511149
transform 1 0 46184 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_507
timestamp 1644511149
transform 1 0 47748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_524
timestamp 1644511149
transform 1 0 49312 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_539
timestamp 1644511149
transform 1 0 50692 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_556
timestamp 1644511149
transform 1 0 52256 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_584
timestamp 1644511149
transform 1 0 54832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_13
timestamp 1644511149
transform 1 0 2300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_20
timestamp 1644511149
transform 1 0 2944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_28
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_76
timestamp 1644511149
transform 1 0 8096 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_88
timestamp 1644511149
transform 1 0 9200 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_100
timestamp 1644511149
transform 1 0 10304 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_133
timestamp 1644511149
transform 1 0 13340 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1644511149
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_176
timestamp 1644511149
transform 1 0 17296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_187
timestamp 1644511149
transform 1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_198
timestamp 1644511149
transform 1 0 19320 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_210
timestamp 1644511149
transform 1 0 20424 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1644511149
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_269
timestamp 1644511149
transform 1 0 25852 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_313
timestamp 1644511149
transform 1 0 29900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_327
timestamp 1644511149
transform 1 0 31188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_341
timestamp 1644511149
transform 1 0 32476 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_358
timestamp 1644511149
transform 1 0 34040 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_370
timestamp 1644511149
transform 1 0 35144 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_382
timestamp 1644511149
transform 1 0 36248 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1644511149
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_452
timestamp 1644511149
transform 1 0 42688 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_464
timestamp 1644511149
transform 1 0 43792 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_471
timestamp 1644511149
transform 1 0 44436 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_483
timestamp 1644511149
transform 1 0 45540 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_495
timestamp 1644511149
transform 1 0 46644 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_548
timestamp 1644511149
transform 1 0 51520 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_45
timestamp 1644511149
transform 1 0 5244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1644511149
transform 1 0 7176 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1644511149
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_102
timestamp 1644511149
transform 1 0 10488 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_114
timestamp 1644511149
transform 1 0 11592 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_126
timestamp 1644511149
transform 1 0 12696 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1644511149
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_151
timestamp 1644511149
transform 1 0 14996 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_159
timestamp 1644511149
transform 1 0 15732 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_166
timestamp 1644511149
transform 1 0 16376 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_174
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_185
timestamp 1644511149
transform 1 0 18124 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1644511149
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_229
timestamp 1644511149
transform 1 0 22172 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_241
timestamp 1644511149
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1644511149
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_259
timestamp 1644511149
transform 1 0 24932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_268
timestamp 1644511149
transform 1 0 25760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_288
timestamp 1644511149
transform 1 0 27600 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_300
timestamp 1644511149
transform 1 0 28704 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_317
timestamp 1644511149
transform 1 0 30268 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_325
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_336
timestamp 1644511149
transform 1 0 32016 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_348
timestamp 1644511149
transform 1 0 33120 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1644511149
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_393
timestamp 1644511149
transform 1 0 37260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_404
timestamp 1644511149
transform 1 0 38272 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1644511149
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_429
timestamp 1644511149
transform 1 0 40572 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_447
timestamp 1644511149
transform 1 0 42228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1644511149
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_502
timestamp 1644511149
transform 1 0 47288 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_509
timestamp 1644511149
transform 1 0 47932 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_521
timestamp 1644511149
transform 1 0 49036 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_529
timestamp 1644511149
transform 1 0 49772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_26
timestamp 1644511149
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1644511149
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1644511149
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_62
timestamp 1644511149
transform 1 0 6808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1644511149
transform 1 0 8648 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1644511149
transform 1 0 9752 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1644511149
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_131
timestamp 1644511149
transform 1 0 13156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_139
timestamp 1644511149
transform 1 0 13892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_157
timestamp 1644511149
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1644511149
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_182
timestamp 1644511149
transform 1 0 17848 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_204
timestamp 1644511149
transform 1 0 19872 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1644511149
transform 1 0 20608 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_231
timestamp 1644511149
transform 1 0 22356 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_239
timestamp 1644511149
transform 1 0 23092 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_256
timestamp 1644511149
transform 1 0 24656 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_268
timestamp 1644511149
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_289
timestamp 1644511149
transform 1 0 27692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_301
timestamp 1644511149
transform 1 0 28796 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_307
timestamp 1644511149
transform 1 0 29348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_316
timestamp 1644511149
transform 1 0 30176 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_350
timestamp 1644511149
transform 1 0 33304 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_363
timestamp 1644511149
transform 1 0 34500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_371
timestamp 1644511149
transform 1 0 35236 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_377
timestamp 1644511149
transform 1 0 35788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1644511149
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_403
timestamp 1644511149
transform 1 0 38180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_415
timestamp 1644511149
transform 1 0 39284 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_427
timestamp 1644511149
transform 1 0 40388 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_439
timestamp 1644511149
transform 1 0 41492 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_468
timestamp 1644511149
transform 1 0 44160 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_480
timestamp 1644511149
transform 1 0 45264 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_492
timestamp 1644511149
transform 1 0 46368 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_521
timestamp 1644511149
transform 1 0 49036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_533
timestamp 1644511149
transform 1 0 50140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_545
timestamp 1644511149
transform 1 0 51244 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_557
timestamp 1644511149
transform 1 0 52348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_567
timestamp 1644511149
transform 1 0 53268 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_571
timestamp 1644511149
transform 1 0 53636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_591
timestamp 1644511149
transform 1 0 55476 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_603
timestamp 1644511149
transform 1 0 56580 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1644511149
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_32
timestamp 1644511149
transform 1 0 4048 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_40
timestamp 1644511149
transform 1 0 4784 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_50
timestamp 1644511149
transform 1 0 5704 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_62
timestamp 1644511149
transform 1 0 6808 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_66
timestamp 1644511149
transform 1 0 7176 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1644511149
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1644511149
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_98
timestamp 1644511149
transform 1 0 10120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1644511149
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_128
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1644511149
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_161
timestamp 1644511149
transform 1 0 15916 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_169
timestamp 1644511149
transform 1 0 16652 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1644511149
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1644511149
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_288
timestamp 1644511149
transform 1 0 27600 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_300
timestamp 1644511149
transform 1 0 28704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_319
timestamp 1644511149
transform 1 0 30452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_331
timestamp 1644511149
transform 1 0 31556 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_339
timestamp 1644511149
transform 1 0 32292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_351
timestamp 1644511149
transform 1 0 33396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_385
timestamp 1644511149
transform 1 0 36524 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_396
timestamp 1644511149
transform 1 0 37536 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_406
timestamp 1644511149
transform 1 0 38456 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_414
timestamp 1644511149
transform 1 0 39192 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_437
timestamp 1644511149
transform 1 0 41308 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_449
timestamp 1644511149
transform 1 0 42412 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_455
timestamp 1644511149
transform 1 0 42964 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1644511149
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_505
timestamp 1644511149
transform 1 0 47564 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_517
timestamp 1644511149
transform 1 0 48668 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_529
timestamp 1644511149
transform 1 0 49772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_7
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_32
timestamp 1644511149
transform 1 0 4048 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_89
timestamp 1644511149
transform 1 0 9292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_131
timestamp 1644511149
transform 1 0 13156 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_136
timestamp 1644511149
transform 1 0 13616 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_147
timestamp 1644511149
transform 1 0 14628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_158
timestamp 1644511149
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1644511149
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_183
timestamp 1644511149
transform 1 0 17940 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_194
timestamp 1644511149
transform 1 0 18952 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_206
timestamp 1644511149
transform 1 0 20056 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1644511149
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_230
timestamp 1644511149
transform 1 0 22264 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_242
timestamp 1644511149
transform 1 0 23368 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_250
timestamp 1644511149
transform 1 0 24104 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_255
timestamp 1644511149
transform 1 0 24564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_267
timestamp 1644511149
transform 1 0 25668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_288
timestamp 1644511149
transform 1 0 27600 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_295
timestamp 1644511149
transform 1 0 28244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_309
timestamp 1644511149
transform 1 0 29532 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_321
timestamp 1644511149
transform 1 0 30636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1644511149
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_345
timestamp 1644511149
transform 1 0 32844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_357
timestamp 1644511149
transform 1 0 33948 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_369
timestamp 1644511149
transform 1 0 35052 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_381
timestamp 1644511149
transform 1 0 36156 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1644511149
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_409
timestamp 1644511149
transform 1 0 38732 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_421
timestamp 1644511149
transform 1 0 39836 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_433
timestamp 1644511149
transform 1 0 40940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1644511149
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_468
timestamp 1644511149
transform 1 0 44160 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_480
timestamp 1644511149
transform 1 0 45264 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_492
timestamp 1644511149
transform 1 0 46368 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1644511149
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1644511149
transform 1 0 5152 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1644511149
transform 1 0 6256 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_68
timestamp 1644511149
transform 1 0 7360 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_72
timestamp 1644511149
transform 1 0 7728 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1644511149
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_102
timestamp 1644511149
transform 1 0 10488 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_114
timestamp 1644511149
transform 1 0 11592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1644511149
transform 1 0 12604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1644511149
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1644511149
transform 1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_161
timestamp 1644511149
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_175
timestamp 1644511149
transform 1 0 17204 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_219
timestamp 1644511149
transform 1 0 21252 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_223
timestamp 1644511149
transform 1 0 21620 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_230
timestamp 1644511149
transform 1 0 22264 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_261
timestamp 1644511149
transform 1 0 25116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_273
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_292
timestamp 1644511149
transform 1 0 27968 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_298
timestamp 1644511149
transform 1 0 28520 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_303
timestamp 1644511149
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_316
timestamp 1644511149
transform 1 0 30176 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_328
timestamp 1644511149
transform 1 0 31280 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_332
timestamp 1644511149
transform 1 0 31648 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_341
timestamp 1644511149
transform 1 0 32476 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_353
timestamp 1644511149
transform 1 0 33580 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1644511149
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_392
timestamp 1644511149
transform 1 0 37168 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_402
timestamp 1644511149
transform 1 0 38088 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_414
timestamp 1644511149
transform 1 0 39192 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_7
timestamp 1644511149
transform 1 0 1748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_24
timestamp 1644511149
transform 1 0 3312 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_31
timestamp 1644511149
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_43
timestamp 1644511149
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_142
timestamp 1644511149
transform 1 0 14168 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_154
timestamp 1644511149
transform 1 0 15272 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1644511149
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_175
timestamp 1644511149
transform 1 0 17204 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_186
timestamp 1644511149
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_197
timestamp 1644511149
transform 1 0 19228 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_203
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_254
timestamp 1644511149
transform 1 0 24472 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_260
timestamp 1644511149
transform 1 0 25024 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_268
timestamp 1644511149
transform 1 0 25760 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_299
timestamp 1644511149
transform 1 0 28612 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_348
timestamp 1644511149
transform 1 0 33120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_359
timestamp 1644511149
transform 1 0 34132 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_368
timestamp 1644511149
transform 1 0 34960 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_380
timestamp 1644511149
transform 1 0 36064 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_410
timestamp 1644511149
transform 1 0 38824 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_422
timestamp 1644511149
transform 1 0 39928 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_434
timestamp 1644511149
transform 1 0 41032 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_446
timestamp 1644511149
transform 1 0 42136 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_11
timestamp 1644511149
transform 1 0 2116 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1644511149
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_72
timestamp 1644511149
transform 1 0 7728 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_104
timestamp 1644511149
transform 1 0 10672 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_120
timestamp 1644511149
transform 1 0 12144 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_128
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_148
timestamp 1644511149
transform 1 0 14720 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_159
timestamp 1644511149
transform 1 0 15732 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_171
timestamp 1644511149
transform 1 0 16836 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_179
timestamp 1644511149
transform 1 0 17572 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_188
timestamp 1644511149
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_204
timestamp 1644511149
transform 1 0 19872 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_216
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_228
timestamp 1644511149
transform 1 0 22080 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_240
timestamp 1644511149
transform 1 0 23184 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_297
timestamp 1644511149
transform 1 0 28428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_355
timestamp 1644511149
transform 1 0 33764 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_369
timestamp 1644511149
transform 1 0 35052 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_386
timestamp 1644511149
transform 1 0 36616 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_398
timestamp 1644511149
transform 1 0 37720 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_410
timestamp 1644511149
transform 1 0 38824 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_418
timestamp 1644511149
transform 1 0 39560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_33
timestamp 1644511149
transform 1 0 4140 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_46
timestamp 1644511149
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1644511149
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_65
timestamp 1644511149
transform 1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_73
timestamp 1644511149
transform 1 0 7820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_85
timestamp 1644511149
transform 1 0 8924 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp 1644511149
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_144
timestamp 1644511149
transform 1 0 14352 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1644511149
transform 1 0 15456 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_192
timestamp 1644511149
transform 1 0 18768 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_204
timestamp 1644511149
transform 1 0 19872 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1644511149
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_231
timestamp 1644511149
transform 1 0 22356 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_243
timestamp 1644511149
transform 1 0 23460 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_262
timestamp 1644511149
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_266
timestamp 1644511149
transform 1 0 25576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_287
timestamp 1644511149
transform 1 0 27508 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_304
timestamp 1644511149
transform 1 0 29072 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_311
timestamp 1644511149
transform 1 0 29716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_323
timestamp 1644511149
transform 1 0 30820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_342
timestamp 1644511149
transform 1 0 32568 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_354
timestamp 1644511149
transform 1 0 33672 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_366
timestamp 1644511149
transform 1 0 34776 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_372
timestamp 1644511149
transform 1 0 35328 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_384
timestamp 1644511149
transform 1 0 36432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_11
timestamp 1644511149
transform 1 0 2116 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1644511149
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1644511149
transform 1 0 4048 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1644511149
transform 1 0 5152 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1644511149
transform 1 0 6256 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1644511149
transform 1 0 7360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_166
timestamp 1644511149
transform 1 0 16376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_188
timestamp 1644511149
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_259
timestamp 1644511149
transform 1 0 24932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_268
timestamp 1644511149
transform 1 0 25760 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_280
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_292
timestamp 1644511149
transform 1 0 27968 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_312
timestamp 1644511149
transform 1 0 29808 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_320
timestamp 1644511149
transform 1 0 30544 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_330
timestamp 1644511149
transform 1 0 31464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_339
timestamp 1644511149
transform 1 0 32292 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_343
timestamp 1644511149
transform 1 0 32660 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_351
timestamp 1644511149
transform 1 0 33396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_25
timestamp 1644511149
transform 1 0 3404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1644511149
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1644511149
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_90
timestamp 1644511149
transform 1 0 9384 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_102
timestamp 1644511149
transform 1 0 10488 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1644511149
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1644511149
transform 1 0 14628 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_159
timestamp 1644511149
transform 1 0 15732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_177
timestamp 1644511149
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_186
timestamp 1644511149
transform 1 0 18216 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_198
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_210
timestamp 1644511149
transform 1 0 20424 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_255
timestamp 1644511149
transform 1 0 24564 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_262
timestamp 1644511149
transform 1 0 25208 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 1644511149
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_289
timestamp 1644511149
transform 1 0 27692 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_298
timestamp 1644511149
transform 1 0 28520 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_310
timestamp 1644511149
transform 1 0 29624 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1644511149
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_345
timestamp 1644511149
transform 1 0 32844 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_363
timestamp 1644511149
transform 1 0 34500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_375
timestamp 1644511149
transform 1 0 35604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_387
timestamp 1644511149
transform 1 0 36708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_6
timestamp 1644511149
transform 1 0 1656 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_13
timestamp 1644511149
transform 1 0 2300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1644511149
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_61
timestamp 1644511149
transform 1 0 6716 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1644511149
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_101
timestamp 1644511149
transform 1 0 10396 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_106
timestamp 1644511149
transform 1 0 10856 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_118
timestamp 1644511149
transform 1 0 11960 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_130
timestamp 1644511149
transform 1 0 13064 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1644511149
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_157
timestamp 1644511149
transform 1 0 15548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_169
timestamp 1644511149
transform 1 0 16652 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_173
timestamp 1644511149
transform 1 0 17020 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_181
timestamp 1644511149
transform 1 0 17756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1644511149
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_269
timestamp 1644511149
transform 1 0 25852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_281
timestamp 1644511149
transform 1 0 26956 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_287
timestamp 1644511149
transform 1 0 27508 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_353
timestamp 1644511149
transform 1 0 33580 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1644511149
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_13
timestamp 1644511149
transform 1 0 2300 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_17
timestamp 1644511149
transform 1 0 2668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_30
timestamp 1644511149
transform 1 0 3864 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_38
timestamp 1644511149
transform 1 0 4600 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_50
timestamp 1644511149
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_85
timestamp 1644511149
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_97
timestamp 1644511149
transform 1 0 10028 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_103
timestamp 1644511149
transform 1 0 10580 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1644511149
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_130
timestamp 1644511149
transform 1 0 13064 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_142
timestamp 1644511149
transform 1 0 14168 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1644511149
transform 1 0 15272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_7
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_11
timestamp 1644511149
transform 1 0 2116 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1644511149
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_45
timestamp 1644511149
transform 1 0 5244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_57
timestamp 1644511149
transform 1 0 6348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_69
timestamp 1644511149
transform 1 0 7452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 1644511149
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1644511149
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_149
timestamp 1644511149
transform 1 0 14812 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_155
timestamp 1644511149
transform 1 0 15364 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_172
timestamp 1644511149
transform 1 0 16928 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_184
timestamp 1644511149
transform 1 0 18032 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_9
timestamp 1644511149
transform 1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_16
timestamp 1644511149
transform 1 0 2576 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_23
timestamp 1644511149
transform 1 0 3220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_36
timestamp 1644511149
transform 1 0 4416 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_48
timestamp 1644511149
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_91
timestamp 1644511149
transform 1 0 9476 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_103
timestamp 1644511149
transform 1 0 10580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_119
timestamp 1644511149
transform 1 0 12052 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_123
timestamp 1644511149
transform 1 0 12420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_133
timestamp 1644511149
transform 1 0 13340 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_145
timestamp 1644511149
transform 1 0 14444 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_157
timestamp 1644511149
transform 1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_165
timestamp 1644511149
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_185
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_197
timestamp 1644511149
transform 1 0 19228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_209
timestamp 1644511149
transform 1 0 20332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1644511149
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_7
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1644511149
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_49
timestamp 1644511149
transform 1 0 5612 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_68
timestamp 1644511149
transform 1 0 7360 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1644511149
transform 1 0 8280 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_93
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_107
timestamp 1644511149
transform 1 0 10948 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_131
timestamp 1644511149
transform 1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_171
timestamp 1644511149
transform 1 0 16836 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_178
timestamp 1644511149
transform 1 0 17480 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1644511149
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_7
timestamp 1644511149
transform 1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_14
timestamp 1644511149
transform 1 0 2392 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_20
timestamp 1644511149
transform 1 0 2944 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_30
timestamp 1644511149
transform 1 0 3864 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_34
timestamp 1644511149
transform 1 0 4232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_65
timestamp 1644511149
transform 1 0 7084 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_84
timestamp 1644511149
transform 1 0 8832 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1644511149
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_121
timestamp 1644511149
transform 1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_140
timestamp 1644511149
transform 1 0 13984 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_160
timestamp 1644511149
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_175
timestamp 1644511149
transform 1 0 17204 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_182
timestamp 1644511149
transform 1 0 17848 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_194
timestamp 1644511149
transform 1 0 18952 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_206
timestamp 1644511149
transform 1 0 20056 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_218
timestamp 1644511149
transform 1 0 21160 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_7
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1644511149
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_45
timestamp 1644511149
transform 1 0 5244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_57
timestamp 1644511149
transform 1 0 6348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_69
timestamp 1644511149
transform 1 0 7452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1644511149
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_170
timestamp 1644511149
transform 1 0 16744 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_190
timestamp 1644511149
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_9
timestamp 1644511149
transform 1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_22
timestamp 1644511149
transform 1 0 3128 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_29
timestamp 1644511149
transform 1 0 3772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_41
timestamp 1644511149
transform 1 0 4876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1644511149
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_73
timestamp 1644511149
transform 1 0 7820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_85
timestamp 1644511149
transform 1 0 8924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_97
timestamp 1644511149
transform 1 0 10028 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_101
timestamp 1644511149
transform 1 0 10396 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_175
timestamp 1644511149
transform 1 0 17204 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_187
timestamp 1644511149
transform 1 0 18308 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_199
timestamp 1644511149
transform 1 0 19412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_211
timestamp 1644511149
transform 1 0 20516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1644511149
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_7
timestamp 1644511149
transform 1 0 1748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1644511149
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_70
timestamp 1644511149
transform 1 0 7544 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1644511149
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_127
timestamp 1644511149
transform 1 0 12788 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 1644511149
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_569
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1644511149
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1644511149
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_613
timestamp 1644511149
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_7
timestamp 1644511149
transform 1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_11
timestamp 1644511149
transform 1 0 2116 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_22
timestamp 1644511149
transform 1 0 3128 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_30
timestamp 1644511149
transform 1 0 3864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1644511149
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_63
timestamp 1644511149
transform 1 0 6900 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_75
timestamp 1644511149
transform 1 0 8004 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_87
timestamp 1644511149
transform 1 0 9108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_91
timestamp 1644511149
transform 1 0 9476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1644511149
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_121
timestamp 1644511149
transform 1 0 12236 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_139
timestamp 1644511149
transform 1 0 13892 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_153
timestamp 1644511149
transform 1 0 15180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_165
timestamp 1644511149
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_179
timestamp 1644511149
transform 1 0 17572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_191
timestamp 1644511149
transform 1 0 18676 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_203
timestamp 1644511149
transform 1 0 19780 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_215
timestamp 1644511149
transform 1 0 20884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1644511149
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_13
timestamp 1644511149
transform 1 0 2300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_25
timestamp 1644511149
transform 1 0 3404 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_39
timestamp 1644511149
transform 1 0 4692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_51
timestamp 1644511149
transform 1 0 5796 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_72
timestamp 1644511149
transform 1 0 7728 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_101
timestamp 1644511149
transform 1 0 10396 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_108
timestamp 1644511149
transform 1 0 11040 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_120
timestamp 1644511149
transform 1 0 12144 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_132
timestamp 1644511149
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_157
timestamp 1644511149
transform 1 0 15548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_185
timestamp 1644511149
transform 1 0 18124 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1644511149
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_545
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_557
timestamp 1644511149
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_569
timestamp 1644511149
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1644511149
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_601
timestamp 1644511149
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_613
timestamp 1644511149
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_13
timestamp 1644511149
transform 1 0 2300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_21
timestamp 1644511149
transform 1 0 3036 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_28
timestamp 1644511149
transform 1 0 3680 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_35
timestamp 1644511149
transform 1 0 4324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1644511149
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_61
timestamp 1644511149
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_78
timestamp 1644511149
transform 1 0 8280 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_90
timestamp 1644511149
transform 1 0 9384 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_102
timestamp 1644511149
transform 1 0 10488 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1644511149
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1644511149
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1644511149
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1644511149
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1644511149
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_7
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1644511149
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_33
timestamp 1644511149
transform 1 0 4140 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_43
timestamp 1644511149
transform 1 0 5060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_55
timestamp 1644511149
transform 1 0 6164 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_68
timestamp 1644511149
transform 1 0 7360 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_75
timestamp 1644511149
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1644511149
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_557
timestamp 1644511149
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_7
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_22
timestamp 1644511149
transform 1 0 3128 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_34
timestamp 1644511149
transform 1 0 4232 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1644511149
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1644511149
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_7
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_14
timestamp 1644511149
transform 1 0 2392 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1644511149
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_37
timestamp 1644511149
transform 1 0 4508 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_13
timestamp 1644511149
transform 1 0 2300 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_25
timestamp 1644511149
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_37
timestamp 1644511149
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_49
timestamp 1644511149
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_6
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_18
timestamp 1644511149
transform 1 0 2760 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1644511149
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1644511149
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1644511149
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_19
timestamp 1644511149
transform 1 0 2852 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_31
timestamp 1644511149
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_43
timestamp 1644511149
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_19
timestamp 1644511149
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_513
timestamp 1644511149
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1644511149
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_20
timestamp 1644511149
transform 1 0 2944 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_32
timestamp 1644511149
transform 1 0 4048 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_44
timestamp 1644511149
transform 1 0 5152 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1644511149
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1644511149
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1644511149
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_597
timestamp 1644511149
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1644511149
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_7
timestamp 1644511149
transform 1 0 1748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 1644511149
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_513
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1644511149
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1644511149
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_7
timestamp 1644511149
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_14
timestamp 1644511149
transform 1 0 2392 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_26
timestamp 1644511149
transform 1 0 3496 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_38
timestamp 1644511149
transform 1 0 4600 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1644511149
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_517
timestamp 1644511149
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_529
timestamp 1644511149
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_541
timestamp 1644511149
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1644511149
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_11
timestamp 1644511149
transform 1 0 2116 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_23
timestamp 1644511149
transform 1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_513
timestamp 1644511149
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_529
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_541
timestamp 1644511149
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1644511149
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_7
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1644511149
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1644511149
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_7
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_31
timestamp 1644511149
transform 1 0 3956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_43
timestamp 1644511149
transform 1 0 5060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1644511149
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1644511149
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_545
timestamp 1644511149
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_557
timestamp 1644511149
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_569
timestamp 1644511149
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1644511149
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1644511149
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_601
timestamp 1644511149
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_613
timestamp 1644511149
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_7
timestamp 1644511149
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_19
timestamp 1644511149
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_31
timestamp 1644511149
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_43
timestamp 1644511149
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_517
timestamp 1644511149
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_529
timestamp 1644511149
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_541
timestamp 1644511149
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1644511149
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1644511149
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_561
timestamp 1644511149
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_573
timestamp 1644511149
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_585
timestamp 1644511149
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_597
timestamp 1644511149
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1644511149
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1644511149
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1644511149
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_7
timestamp 1644511149
transform 1 0 1748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_19
timestamp 1644511149
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_501
timestamp 1644511149
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_513
timestamp 1644511149
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1644511149
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1644511149
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_533
timestamp 1644511149
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_545
timestamp 1644511149
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_557
timestamp 1644511149
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_569
timestamp 1644511149
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1644511149
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1644511149
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_589
timestamp 1644511149
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_601
timestamp 1644511149
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_613
timestamp 1644511149
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_7
timestamp 1644511149
transform 1 0 1748 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_19
timestamp 1644511149
transform 1 0 2852 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_31
timestamp 1644511149
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_43
timestamp 1644511149
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_372
timestamp 1644511149
transform 1 0 35328 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_384
timestamp 1644511149
transform 1 0 36432 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_517
timestamp 1644511149
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_529
timestamp 1644511149
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_541
timestamp 1644511149
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1644511149
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1644511149
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_561
timestamp 1644511149
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_573
timestamp 1644511149
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_585
timestamp 1644511149
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_597
timestamp 1644511149
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1644511149
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1644511149
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1644511149
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_7
timestamp 1644511149
transform 1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_23
timestamp 1644511149
transform 1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_33
timestamp 1644511149
transform 1 0 4140 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_37
timestamp 1644511149
transform 1 0 4508 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_49
timestamp 1644511149
transform 1 0 5612 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_55
timestamp 1644511149
transform 1 0 6164 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_57
timestamp 1644511149
transform 1 0 6348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_69
timestamp 1644511149
transform 1 0 7452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_81
timestamp 1644511149
transform 1 0 8556 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_113
timestamp 1644511149
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_125
timestamp 1644511149
transform 1 0 12604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_137
timestamp 1644511149
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_169
timestamp 1644511149
transform 1 0 16652 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_181
timestamp 1644511149
transform 1 0 17756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_193
timestamp 1644511149
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_200
timestamp 1644511149
transform 1 0 19504 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_212
timestamp 1644511149
transform 1 0 20608 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_225
timestamp 1644511149
transform 1 0 21804 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_237
timestamp 1644511149
transform 1 0 22908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_249
timestamp 1644511149
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_285
timestamp 1644511149
transform 1 0 27324 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_297
timestamp 1644511149
transform 1 0 28428 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_305
timestamp 1644511149
transform 1 0 29164 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_337
timestamp 1644511149
transform 1 0 32108 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_349
timestamp 1644511149
transform 1 0 33212 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_359
timestamp 1644511149
transform 1 0 34132 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_393
timestamp 1644511149
transform 1 0 37260 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_405
timestamp 1644511149
transform 1 0 38364 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_417
timestamp 1644511149
transform 1 0 39468 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_439
timestamp 1644511149
transform 1 0 41492 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_447
timestamp 1644511149
transform 1 0 42228 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_449
timestamp 1644511149
transform 1 0 42412 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_461
timestamp 1644511149
transform 1 0 43516 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_473
timestamp 1644511149
transform 1 0 44620 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_501
timestamp 1644511149
transform 1 0 47196 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_505
timestamp 1644511149
transform 1 0 47564 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_517
timestamp 1644511149
transform 1 0 48668 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_521
timestamp 1644511149
transform 1 0 49036 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_529
timestamp 1644511149
transform 1 0 49772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_533
timestamp 1644511149
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_545
timestamp 1644511149
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_557
timestamp 1644511149
transform 1 0 52348 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_561
timestamp 1644511149
transform 1 0 52716 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_573
timestamp 1644511149
transform 1 0 53820 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_585
timestamp 1644511149
transform 1 0 54924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_589
timestamp 1644511149
transform 1 0 55292 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_597
timestamp 1644511149
transform 1 0 56028 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_603
timestamp 1644511149
transform 1 0 56580 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_615
timestamp 1644511149
transform 1 0 57684 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_617
timestamp 1644511149
transform 1 0 57868 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_1
timestamp 1644511149
transform -1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_2
timestamp 1644511149
transform 1 0 12052 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_3
timestamp 1644511149
transform 1 0 12236 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_4
timestamp 1644511149
transform 1 0 24564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_5
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_6
timestamp 1644511149
transform 1 0 23000 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_7
timestamp 1644511149
transform -1 0 23184 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_8
timestamp 1644511149
transform 1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_9
timestamp 1644511149
transform -1 0 43516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_10
timestamp 1644511149
transform -1 0 4508 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_11
timestamp 1644511149
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_12
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_13
timestamp 1644511149
transform 1 0 14720 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_14
timestamp 1644511149
transform 1 0 23184 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_15
timestamp 1644511149
transform 1 0 23920 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_16
timestamp 1644511149
transform 1 0 25024 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_17
timestamp 1644511149
transform 1 0 25116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_18
timestamp 1644511149
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_19
timestamp 1644511149
transform 1 0 24840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_20
timestamp 1644511149
transform 1 0 28336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_21
timestamp 1644511149
transform 1 0 19872 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_22
timestamp 1644511149
transform 1 0 21712 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 32016 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 42320 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 47472 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 52624 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 57776 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0677_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0678_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0679_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0680_
timestamp 1644511149
transform 1 0 15180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0681_
timestamp 1644511149
transform 1 0 15272 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0682_
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0683_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4416 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0684_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0685_
timestamp 1644511149
transform 1 0 3496 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0686_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0687_
timestamp 1644511149
transform 1 0 42596 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0688_
timestamp 1644511149
transform 1 0 43884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _0689_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35696 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 1644511149
transform 1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0692_
timestamp 1644511149
transform 1 0 10948 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0693_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0694_
timestamp 1644511149
transform 1 0 8372 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0695_
timestamp 1644511149
transform 1 0 8188 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0696_
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1644511149
transform 1 0 10580 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0698_
timestamp 1644511149
transform 1 0 11408 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0699_
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0700_
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0701_
timestamp 1644511149
transform 1 0 11592 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0702_
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0703_
timestamp 1644511149
transform 1 0 11776 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0704_
timestamp 1644511149
transform 1 0 13248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0705_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6716 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0706_
timestamp 1644511149
transform 1 0 3772 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0707_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7360 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0708_
timestamp 1644511149
transform 1 0 4876 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_2  _0709_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9016 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0710_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6440 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0711_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8096 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0712_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7268 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0713_
timestamp 1644511149
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0714_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1644511149
transform 1 0 47656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0716_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_4  _0717_
timestamp 1644511149
transform 1 0 48576 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0718_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0719_
timestamp 1644511149
transform 1 0 35052 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0720_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0721_
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_2  _0722_
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0723_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0724_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0725_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_4  _0726_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6900 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__a2111o_1  _0727_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6900 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0728_
timestamp 1644511149
transform 1 0 10120 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0729_
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0730_
timestamp 1644511149
transform 1 0 12604 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0731_
timestamp 1644511149
transform 1 0 27876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0732_
timestamp 1644511149
transform 1 0 7176 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0733_
timestamp 1644511149
transform 1 0 10396 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0734_
timestamp 1644511149
transform 1 0 10580 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_4  _0735_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10212 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0736_
timestamp 1644511149
transform 1 0 22632 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0737_
timestamp 1644511149
transform 1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0738_
timestamp 1644511149
transform 1 0 21896 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0739_
timestamp 1644511149
transform 1 0 36340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0740_
timestamp 1644511149
transform 1 0 35328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0741_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31004 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0742_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30912 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1644511149
transform 1 0 8096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0744_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0745_
timestamp 1644511149
transform 1 0 23460 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0746_
timestamp 1644511149
transform 1 0 25392 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0747_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0748_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0749_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29072 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0750_
timestamp 1644511149
transform 1 0 23920 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0751_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0752_
timestamp 1644511149
transform 1 0 28152 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 1644511149
transform 1 0 28612 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0754_
timestamp 1644511149
transform 1 0 20240 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0755_
timestamp 1644511149
transform 1 0 19044 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0756_
timestamp 1644511149
transform 1 0 30176 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0757_
timestamp 1644511149
transform 1 0 24932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0758_
timestamp 1644511149
transform 1 0 24656 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0759_
timestamp 1644511149
transform 1 0 24748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0760_
timestamp 1644511149
transform 1 0 19228 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0761_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1644511149
transform 1 0 18400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0763_
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0764_
timestamp 1644511149
transform 1 0 18216 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0765_
timestamp 1644511149
transform 1 0 20240 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0766_
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0767_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0768_
timestamp 1644511149
transform 1 0 22080 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0769_
timestamp 1644511149
transform 1 0 21252 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0770_
timestamp 1644511149
transform 1 0 21068 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0771_
timestamp 1644511149
transform 1 0 23368 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1644511149
transform 1 0 23368 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0773_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0774_
timestamp 1644511149
transform 1 0 30360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0775_
timestamp 1644511149
transform 1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0776_
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0777_
timestamp 1644511149
transform 1 0 21160 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0778_
timestamp 1644511149
transform 1 0 22448 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0779_
timestamp 1644511149
transform 1 0 21068 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0780_
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0781_
timestamp 1644511149
transform 1 0 23552 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0782_
timestamp 1644511149
transform 1 0 22264 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0783_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0784_
timestamp 1644511149
transform 1 0 23000 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0785_
timestamp 1644511149
transform 1 0 23920 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0786_
timestamp 1644511149
transform 1 0 24656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0787_
timestamp 1644511149
transform 1 0 22080 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0788_
timestamp 1644511149
transform 1 0 28152 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0789_
timestamp 1644511149
transform 1 0 25208 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0790_
timestamp 1644511149
transform 1 0 25668 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0791_
timestamp 1644511149
transform 1 0 24380 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0792_
timestamp 1644511149
transform 1 0 25760 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0793_
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0794_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1644511149
transform 1 0 25944 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0796_
timestamp 1644511149
transform 1 0 24288 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0797_
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0798_
timestamp 1644511149
transform 1 0 28796 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0799_
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0800_
timestamp 1644511149
transform 1 0 30728 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0801_
timestamp 1644511149
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0802_
timestamp 1644511149
transform 1 0 22908 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0803_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0804_
timestamp 1644511149
transform 1 0 29716 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0805_
timestamp 1644511149
transform 1 0 28244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0806_
timestamp 1644511149
transform 1 0 32568 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0807_
timestamp 1644511149
transform 1 0 21896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0808_
timestamp 1644511149
transform 1 0 37628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0809_
timestamp 1644511149
transform 1 0 32844 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0810_
timestamp 1644511149
transform 1 0 28428 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0811_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0812_
timestamp 1644511149
transform 1 0 28152 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0813_
timestamp 1644511149
transform 1 0 27048 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0814_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0815_
timestamp 1644511149
transform 1 0 25300 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0816_
timestamp 1644511149
transform 1 0 25944 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0817_
timestamp 1644511149
transform 1 0 28612 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0818_
timestamp 1644511149
transform 1 0 27968 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0819_
timestamp 1644511149
transform 1 0 27140 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0820_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0821_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0822_
timestamp 1644511149
transform 1 0 28704 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0823_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28612 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0825_
timestamp 1644511149
transform 1 0 26128 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0826_
timestamp 1644511149
transform 1 0 24748 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0827_
timestamp 1644511149
transform 1 0 24748 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0828_
timestamp 1644511149
transform 1 0 27876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1644511149
transform 1 0 29440 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0830_
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0831_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0832_
timestamp 1644511149
transform 1 0 25300 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0833_
timestamp 1644511149
transform 1 0 27968 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0834_
timestamp 1644511149
transform 1 0 31832 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0835_
timestamp 1644511149
transform 1 0 32292 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0836_
timestamp 1644511149
transform 1 0 21804 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0837_
timestamp 1644511149
transform 1 0 30820 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0838_
timestamp 1644511149
transform 1 0 32752 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0839_
timestamp 1644511149
transform 1 0 25944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0840_
timestamp 1644511149
transform 1 0 25760 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0841_
timestamp 1644511149
transform 1 0 33028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0842_
timestamp 1644511149
transform 1 0 23368 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0843_
timestamp 1644511149
transform 1 0 33488 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0844_
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0845_
timestamp 1644511149
transform 1 0 33304 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0846_
timestamp 1644511149
transform 1 0 34500 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0847_
timestamp 1644511149
transform 1 0 35052 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0848_
timestamp 1644511149
transform 1 0 37812 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0849_
timestamp 1644511149
transform 1 0 36616 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0851_
timestamp 1644511149
transform 1 0 36432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0852_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37536 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0853_
timestamp 1644511149
transform 1 0 25208 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0854_
timestamp 1644511149
transform 1 0 37168 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0855_
timestamp 1644511149
transform 1 0 37076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0856_
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _0857_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38824 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0858_
timestamp 1644511149
transform 1 0 37904 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0859_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0860_
timestamp 1644511149
transform 1 0 37628 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1644511149
transform 1 0 48484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0862_
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0863_
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0864_
timestamp 1644511149
transform 1 0 53268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _0865_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47840 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0866_
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0867_
timestamp 1644511149
transform 1 0 46276 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0868_
timestamp 1644511149
transform 1 0 47564 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0869_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 51428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0870_
timestamp 1644511149
transform 1 0 51336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0871_
timestamp 1644511149
transform 1 0 51612 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0872_
timestamp 1644511149
transform 1 0 50600 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0873_
timestamp 1644511149
transform 1 0 50784 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0874_
timestamp 1644511149
transform 1 0 51796 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0875_
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0876_
timestamp 1644511149
transform 1 0 53912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0877_
timestamp 1644511149
transform 1 0 54372 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0878_
timestamp 1644511149
transform 1 0 55016 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0879_
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0880_
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0881_
timestamp 1644511149
transform 1 0 55016 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0882_
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0883_
timestamp 1644511149
transform 1 0 55660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0884_
timestamp 1644511149
transform 1 0 53912 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0885_
timestamp 1644511149
transform 1 0 53912 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0886_
timestamp 1644511149
transform 1 0 53176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0887_
timestamp 1644511149
transform 1 0 52164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0888_
timestamp 1644511149
transform 1 0 52900 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0889_
timestamp 1644511149
transform 1 0 51336 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0890_
timestamp 1644511149
transform 1 0 51244 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0891_
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0892_
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0893_
timestamp 1644511149
transform 1 0 49864 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0894_
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 1644511149
transform 1 0 48208 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0896_
timestamp 1644511149
transform 1 0 49036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0897_
timestamp 1644511149
transform 1 0 47380 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0898_
timestamp 1644511149
transform 1 0 47840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0899_
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0900_
timestamp 1644511149
transform 1 0 45632 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1644511149
transform 1 0 46000 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0902_
timestamp 1644511149
transform 1 0 36156 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0903_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35328 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0904_
timestamp 1644511149
transform 1 0 36340 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 35144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0907_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36524 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0908_
timestamp 1644511149
transform 1 0 35236 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0909_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0910_
timestamp 1644511149
transform 1 0 30820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0911_
timestamp 1644511149
transform 1 0 30636 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0912_
timestamp 1644511149
transform 1 0 14168 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0913_
timestamp 1644511149
transform 1 0 24472 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0914_
timestamp 1644511149
transform 1 0 22724 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0915_
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0916_
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0917_
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0918_
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _0919_
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0920_
timestamp 1644511149
transform 1 0 20976 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0921_
timestamp 1644511149
transform 1 0 18768 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0922_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0923_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0924_
timestamp 1644511149
transform 1 0 19964 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1644511149
transform 1 0 18952 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0926_
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0927_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0928_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0929_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0930_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _0931_
timestamp 1644511149
transform 1 0 33304 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0932_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0933_
timestamp 1644511149
transform 1 0 24748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0934_
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0935_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0936_
timestamp 1644511149
transform 1 0 20792 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0937_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1644511149
transform 1 0 24656 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0939_
timestamp 1644511149
transform 1 0 24196 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0940_
timestamp 1644511149
transform 1 0 23368 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0941_
timestamp 1644511149
transform 1 0 13064 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0942_
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0943_
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0944_
timestamp 1644511149
transform 1 0 14628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0945_
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0946_
timestamp 1644511149
transform 1 0 42596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1644511149
transform 1 0 41032 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0949_
timestamp 1644511149
transform 1 0 38548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0950_
timestamp 1644511149
transform 1 0 34960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0951_
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0952_
timestamp 1644511149
transform 1 0 35604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0953_
timestamp 1644511149
transform 1 0 42412 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0954_
timestamp 1644511149
transform 1 0 36708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0955_
timestamp 1644511149
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0956_
timestamp 1644511149
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0957_
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0958_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39100 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0959_
timestamp 1644511149
transform 1 0 38824 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0960_
timestamp 1644511149
transform 1 0 38916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0961_
timestamp 1644511149
transform 1 0 37628 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0962_
timestamp 1644511149
transform 1 0 38732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1644511149
transform 1 0 36156 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0964_
timestamp 1644511149
transform 1 0 36340 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0965_
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a32o_1  _0966_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0967_
timestamp 1644511149
transform 1 0 45908 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0968_
timestamp 1644511149
transform 1 0 49220 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0969_
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0970_
timestamp 1644511149
transform 1 0 48576 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0971_
timestamp 1644511149
transform 1 0 36340 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0972_
timestamp 1644511149
transform 1 0 36708 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0973_
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0974_
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0975_
timestamp 1644511149
transform 1 0 38088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0976_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 49588 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0977_
timestamp 1644511149
transform 1 0 6624 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0978_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7544 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0979_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7728 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0980_
timestamp 1644511149
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _0981_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12420 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  _0982_
timestamp 1644511149
transform 1 0 27784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0983_
timestamp 1644511149
transform 1 0 37444 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0984_
timestamp 1644511149
transform 1 0 28152 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0985_
timestamp 1644511149
transform 1 0 27784 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0986_
timestamp 1644511149
transform 1 0 49128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0987_
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0988_
timestamp 1644511149
transform 1 0 45264 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0989_
timestamp 1644511149
transform 1 0 46184 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0990_
timestamp 1644511149
transform 1 0 46000 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0991_
timestamp 1644511149
transform 1 0 48576 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0992_
timestamp 1644511149
transform 1 0 27324 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0993_
timestamp 1644511149
transform 1 0 49128 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0994_
timestamp 1644511149
transform 1 0 50232 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0995_
timestamp 1644511149
transform 1 0 44712 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0996_
timestamp 1644511149
transform 1 0 30084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0997_
timestamp 1644511149
transform 1 0 41216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0998_
timestamp 1644511149
transform 1 0 50600 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0999_
timestamp 1644511149
transform 1 0 51980 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1000_
timestamp 1644511149
transform 1 0 27784 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1001_
timestamp 1644511149
transform 1 0 52440 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1002_
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1644511149
transform 1 0 28428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1004_
timestamp 1644511149
transform 1 0 27600 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1005_
timestamp 1644511149
transform 1 0 52532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1006_
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1007_
timestamp 1644511149
transform 1 0 41952 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1008_
timestamp 1644511149
transform 1 0 25668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1009_
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1010_
timestamp 1644511149
transform 1 0 41400 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1011_
timestamp 1644511149
transform 1 0 31188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1012_
timestamp 1644511149
transform 1 0 42688 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1013_
timestamp 1644511149
transform 1 0 30452 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1014_
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1015_
timestamp 1644511149
transform 1 0 42688 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1016_
timestamp 1644511149
transform 1 0 38088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1017_
timestamp 1644511149
transform 1 0 45908 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1018_
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1019_
timestamp 1644511149
transform 1 0 40572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1020_
timestamp 1644511149
transform 1 0 46000 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1021_
timestamp 1644511149
transform 1 0 40112 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1022_
timestamp 1644511149
transform 1 0 25300 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1023_
timestamp 1644511149
transform 1 0 39744 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1024_
timestamp 1644511149
transform 1 0 42596 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1025_
timestamp 1644511149
transform 1 0 38548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1026_
timestamp 1644511149
transform 1 0 41676 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1027_
timestamp 1644511149
transform 1 0 42136 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1028_
timestamp 1644511149
transform 1 0 43976 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1029_
timestamp 1644511149
transform 1 0 44344 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1030_
timestamp 1644511149
transform 1 0 45908 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1031_
timestamp 1644511149
transform 1 0 28704 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1032_
timestamp 1644511149
transform 1 0 46920 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1033_
timestamp 1644511149
transform 1 0 43424 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1034_
timestamp 1644511149
transform 1 0 42780 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1035_
timestamp 1644511149
transform 1 0 43056 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1036_
timestamp 1644511149
transform 1 0 32016 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1037_
timestamp 1644511149
transform 1 0 24104 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1038_
timestamp 1644511149
transform 1 0 29900 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1039_
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1040_
timestamp 1644511149
transform 1 0 26312 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1041_
timestamp 1644511149
transform 1 0 25024 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1042_
timestamp 1644511149
transform 1 0 25300 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1043_
timestamp 1644511149
transform 1 0 36064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1044_
timestamp 1644511149
transform 1 0 27140 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1045_
timestamp 1644511149
transform 1 0 26128 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1046_
timestamp 1644511149
transform 1 0 25484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1047_
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1048_
timestamp 1644511149
transform 1 0 27232 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1049_
timestamp 1644511149
transform 1 0 27600 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1050_
timestamp 1644511149
transform 1 0 29440 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1051_
timestamp 1644511149
transform 1 0 28336 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1052_
timestamp 1644511149
transform 1 0 28612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1053_
timestamp 1644511149
transform 1 0 32292 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1054_
timestamp 1644511149
transform 1 0 32292 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1055_
timestamp 1644511149
transform 1 0 32292 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1056_
timestamp 1644511149
transform 1 0 28704 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1057_
timestamp 1644511149
transform 1 0 32476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1058_
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1059_
timestamp 1644511149
transform 1 0 35052 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1060_
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 1644511149
transform 1 0 33304 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1062_
timestamp 1644511149
transform 1 0 33304 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1063_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38640 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1064_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36800 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1065_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36432 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1066_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34868 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1067_
timestamp 1644511149
transform 1 0 36248 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1068_
timestamp 1644511149
transform 1 0 36708 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1069_
timestamp 1644511149
transform 1 0 39560 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1070_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38456 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1071_
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1644511149
transform 1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1073_
timestamp 1644511149
transform 1 0 37812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1074_
timestamp 1644511149
transform 1 0 37076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1075_
timestamp 1644511149
transform 1 0 35696 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1076_
timestamp 1644511149
transform 1 0 31096 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1077_
timestamp 1644511149
transform 1 0 30452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1078_
timestamp 1644511149
transform 1 0 34500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1079_
timestamp 1644511149
transform 1 0 35604 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1080_
timestamp 1644511149
transform 1 0 35512 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1081_
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1082_
timestamp 1644511149
transform 1 0 33396 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1083_
timestamp 1644511149
transform 1 0 36340 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1084_
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1085_
timestamp 1644511149
transform 1 0 9752 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_1  _1086_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35696 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1087_
timestamp 1644511149
transform 1 0 38364 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _1089_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42412 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1090_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40664 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1091_
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a2111oi_2  _1092_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41768 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _1093_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1644511149
transform 1 0 40388 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1095_
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1096_
timestamp 1644511149
transform 1 0 43424 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1097_
timestamp 1644511149
transform 1 0 42504 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1098_
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1099_
timestamp 1644511149
transform 1 0 38456 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1100_
timestamp 1644511149
transform 1 0 42780 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1101_
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1102_
timestamp 1644511149
transform 1 0 38548 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1103_
timestamp 1644511149
transform 1 0 40756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _1104_
timestamp 1644511149
transform 1 0 40204 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1105_
timestamp 1644511149
transform 1 0 36064 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1644511149
transform 1 0 53360 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1644511149
transform 1 0 43608 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1108_
timestamp 1644511149
transform 1 0 41400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1109_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42504 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _1110_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43608 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1111_
timestamp 1644511149
transform 1 0 45724 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1112_
timestamp 1644511149
transform 1 0 40204 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1113_
timestamp 1644511149
transform 1 0 46368 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1114_
timestamp 1644511149
transform 1 0 46552 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1115_
timestamp 1644511149
transform 1 0 47656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1644511149
transform 1 0 46644 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1117_
timestamp 1644511149
transform 1 0 47656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1118_
timestamp 1644511149
transform 1 0 46828 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1119_
timestamp 1644511149
transform 1 0 47288 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1120_
timestamp 1644511149
transform 1 0 43884 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1121_
timestamp 1644511149
transform 1 0 44068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1122_
timestamp 1644511149
transform 1 0 43700 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1123_
timestamp 1644511149
transform 1 0 43884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1124_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42596 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1126_
timestamp 1644511149
transform 1 0 6992 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1127_
timestamp 1644511149
transform 1 0 12880 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1128_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1129_
timestamp 1644511149
transform 1 0 31464 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1130_
timestamp 1644511149
transform 1 0 31648 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1131_
timestamp 1644511149
transform 1 0 9844 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1132_
timestamp 1644511149
transform 1 0 9844 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1133_
timestamp 1644511149
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1134_
timestamp 1644511149
transform 1 0 10948 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1135_
timestamp 1644511149
transform 1 0 14076 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _1136_
timestamp 1644511149
transform 1 0 12144 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  _1137_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16008 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1138_
timestamp 1644511149
transform 1 0 15824 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_4  _1139_
timestamp 1644511149
transform 1 0 6900 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__o21a_4  _1140_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4_4  _1141_
timestamp 1644511149
transform 1 0 12052 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_1  _1142_
timestamp 1644511149
transform 1 0 12880 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1143_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1144_
timestamp 1644511149
transform 1 0 14720 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1145_
timestamp 1644511149
transform 1 0 16008 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1146_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1147_
timestamp 1644511149
transform 1 0 12696 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1148_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1149_
timestamp 1644511149
transform 1 0 10028 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1150_
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1151_
timestamp 1644511149
transform 1 0 11684 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1152_
timestamp 1644511149
transform 1 0 11776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1153_
timestamp 1644511149
transform 1 0 10580 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1154_
timestamp 1644511149
transform 1 0 10488 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1155_
timestamp 1644511149
transform 1 0 5520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1156_
timestamp 1644511149
transform 1 0 14444 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1157_
timestamp 1644511149
transform 1 0 15916 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1158_
timestamp 1644511149
transform 1 0 14996 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1159_
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1160_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1161_
timestamp 1644511149
transform 1 0 14904 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1162_
timestamp 1644511149
transform 1 0 13156 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1163_
timestamp 1644511149
transform 1 0 15088 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1164_
timestamp 1644511149
transform 1 0 15548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1165_
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1166_
timestamp 1644511149
transform 1 0 16928 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1167_
timestamp 1644511149
transform 1 0 15272 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1168_
timestamp 1644511149
transform 1 0 15180 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1169_
timestamp 1644511149
transform 1 0 4784 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1170_
timestamp 1644511149
transform 1 0 15640 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1171_
timestamp 1644511149
transform 1 0 14628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1172_
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1173_
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1174_
timestamp 1644511149
transform 1 0 5888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1175_
timestamp 1644511149
transform 1 0 14628 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1176_
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1177_
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1178_
timestamp 1644511149
transform 1 0 15272 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1179_
timestamp 1644511149
transform 1 0 5244 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1180_
timestamp 1644511149
transform 1 0 16008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1181_
timestamp 1644511149
transform 1 0 16008 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1182_
timestamp 1644511149
transform 1 0 14996 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1183_
timestamp 1644511149
transform 1 0 5152 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1184_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1185_
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1186_
timestamp 1644511149
transform 1 0 15456 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1187_
timestamp 1644511149
transform 1 0 4876 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1188_
timestamp 1644511149
transform 1 0 5612 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1189_
timestamp 1644511149
transform 1 0 24656 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1190_
timestamp 1644511149
transform 1 0 22816 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1191_
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1192_
timestamp 1644511149
transform 1 0 17204 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1193_
timestamp 1644511149
transform 1 0 16836 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1194_
timestamp 1644511149
transform 1 0 16836 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1195_
timestamp 1644511149
transform 1 0 15548 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1196_
timestamp 1644511149
transform 1 0 4048 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1197_
timestamp 1644511149
transform 1 0 16100 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1198_
timestamp 1644511149
transform 1 0 21988 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1199_
timestamp 1644511149
transform 1 0 17572 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1200_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1201_
timestamp 1644511149
transform 1 0 2300 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1202_
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1203_
timestamp 1644511149
transform 1 0 14168 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1204_
timestamp 1644511149
transform 1 0 25576 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1205_
timestamp 1644511149
transform 1 0 24748 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1206_
timestamp 1644511149
transform 1 0 14996 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1207_
timestamp 1644511149
transform 1 0 15824 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1208_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1209_
timestamp 1644511149
transform 1 0 17296 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1210_
timestamp 1644511149
transform 1 0 16836 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1211_
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1212_
timestamp 1644511149
transform 1 0 24748 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1213_
timestamp 1644511149
transform 1 0 17664 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1214_
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1215_
timestamp 1644511149
transform 1 0 3772 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1216_
timestamp 1644511149
transform 1 0 24656 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1217_
timestamp 1644511149
transform 1 0 17848 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1218_
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1219_
timestamp 1644511149
transform 1 0 2300 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1220_
timestamp 1644511149
transform 1 0 13340 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1221_
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1222_
timestamp 1644511149
transform 1 0 29716 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1223_
timestamp 1644511149
transform 1 0 29624 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1224_
timestamp 1644511149
transform 1 0 17664 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1225_
timestamp 1644511149
transform 1 0 17664 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1226_
timestamp 1644511149
transform 1 0 17204 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1227_
timestamp 1644511149
transform 1 0 16652 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1228_
timestamp 1644511149
transform 1 0 7820 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1229_
timestamp 1644511149
transform 1 0 17020 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1230_
timestamp 1644511149
transform 1 0 31004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1231_
timestamp 1644511149
transform 1 0 17940 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1232_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1233_
timestamp 1644511149
transform 1 0 7268 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1234_
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1235_
timestamp 1644511149
transform 1 0 16836 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1236_
timestamp 1644511149
transform 1 0 18216 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1237_
timestamp 1644511149
transform 1 0 17204 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1238_
timestamp 1644511149
transform 1 0 10120 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1239_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1240_
timestamp 1644511149
transform 1 0 18676 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1241_
timestamp 1644511149
transform 1 0 18124 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1242_
timestamp 1644511149
transform 1 0 14076 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1243_
timestamp 1644511149
transform 1 0 29440 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1244_
timestamp 1644511149
transform 1 0 19228 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1245_
timestamp 1644511149
transform 1 0 18308 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1246_
timestamp 1644511149
transform 1 0 15640 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1247_
timestamp 1644511149
transform 1 0 14444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1248_
timestamp 1644511149
transform 1 0 30728 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _1249_
timestamp 1644511149
transform 1 0 12788 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1250_
timestamp 1644511149
transform 1 0 32384 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1251_
timestamp 1644511149
transform 1 0 31096 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1252_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1253_
timestamp 1644511149
transform 1 0 13248 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1254_
timestamp 1644511149
transform 1 0 13984 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1255_
timestamp 1644511149
transform 1 0 17572 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1256_
timestamp 1644511149
transform 1 0 18584 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1257_
timestamp 1644511149
transform 1 0 17296 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1258_
timestamp 1644511149
transform 1 0 17756 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1259_
timestamp 1644511149
transform 1 0 16928 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1260_
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1261_
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1262_
timestamp 1644511149
transform 1 0 18124 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1263_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1264_
timestamp 1644511149
transform 1 0 17296 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1265_
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1266_
timestamp 1644511149
transform 1 0 14996 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1267_
timestamp 1644511149
transform 1 0 17756 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1268_
timestamp 1644511149
transform 1 0 17572 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1269_
timestamp 1644511149
transform 1 0 17020 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1270_
timestamp 1644511149
transform 1 0 32384 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1271_
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1272_
timestamp 1644511149
transform 1 0 17112 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1273_
timestamp 1644511149
transform 1 0 14628 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _1274_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32568 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1275_
timestamp 1644511149
transform 1 0 17112 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1276_
timestamp 1644511149
transform 1 0 15732 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1277_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1278_
timestamp 1644511149
transform 1 0 11684 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_2  _1279_
timestamp 1644511149
transform 1 0 33212 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1280_
timestamp 1644511149
transform 1 0 15456 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1281_
timestamp 1644511149
transform 1 0 15088 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1282_
timestamp 1644511149
transform 1 0 10488 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _1283_
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1284_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1285_
timestamp 1644511149
transform 1 0 13984 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1286_
timestamp 1644511149
transform 1 0 12880 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _1287_
timestamp 1644511149
transform 1 0 33672 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1288_
timestamp 1644511149
transform 1 0 14168 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1289_
timestamp 1644511149
transform 1 0 14996 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1290_
timestamp 1644511149
transform 1 0 10488 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1291_
timestamp 1644511149
transform 1 0 15456 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1292_
timestamp 1644511149
transform 1 0 12512 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1293_
timestamp 1644511149
transform 1 0 12420 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1294_
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1295_
timestamp 1644511149
transform 1 0 10672 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1296_
timestamp 1644511149
transform 1 0 10212 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1297_
timestamp 1644511149
transform 1 0 11316 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1298_
timestamp 1644511149
transform 1 0 8740 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1299_
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1300_
timestamp 1644511149
transform 1 0 9292 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1301_
timestamp 1644511149
transform 1 0 11224 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1302_
timestamp 1644511149
transform 1 0 8648 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1303_
timestamp 1644511149
transform 1 0 9844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1304_
timestamp 1644511149
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1305_
timestamp 1644511149
transform 1 0 8648 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1306_
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1307_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_4  _1308_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1309_
timestamp 1644511149
transform 1 0 3864 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1310_
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1311_
timestamp 1644511149
transform 1 0 3404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1312_
timestamp 1644511149
transform 1 0 2116 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1313_
timestamp 1644511149
transform 1 0 2668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1314_
timestamp 1644511149
transform 1 0 2116 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1315_
timestamp 1644511149
transform 1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1316_
timestamp 1644511149
transform 1 0 2116 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1317_
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1318_
timestamp 1644511149
transform 1 0 2116 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1319_
timestamp 1644511149
transform 1 0 3404 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1320_
timestamp 1644511149
transform 1 0 6440 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1321_
timestamp 1644511149
transform 1 0 4508 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1322_
timestamp 1644511149
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1323_
timestamp 1644511149
transform 1 0 6532 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1324_
timestamp 1644511149
transform 1 0 6716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1325_
timestamp 1644511149
transform 1 0 6624 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1327_
timestamp 1644511149
transform 1 0 6348 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1328_
timestamp 1644511149
transform 1 0 6900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1329_
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1330_
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1331_
timestamp 1644511149
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1332_
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1333_
timestamp 1644511149
transform 1 0 2576 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1334_
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1335_
timestamp 1644511149
transform 1 0 2668 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1336_
timestamp 1644511149
transform 1 0 3036 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1337_
timestamp 1644511149
transform 1 0 2392 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1338_
timestamp 1644511149
transform 1 0 2208 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1339_
timestamp 1644511149
transform 1 0 2300 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1340_
timestamp 1644511149
transform 1 0 2576 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1341_
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1342_
timestamp 1644511149
transform 1 0 4324 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1343_
timestamp 1644511149
transform 1 0 3036 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1344_
timestamp 1644511149
transform 1 0 3036 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1345_
timestamp 1644511149
transform 1 0 2300 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1346_
timestamp 1644511149
transform 1 0 2208 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1347_
timestamp 1644511149
transform 1 0 3864 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1348_
timestamp 1644511149
transform 1 0 4048 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1349_
timestamp 1644511149
transform 1 0 2300 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1350_
timestamp 1644511149
transform 1 0 3404 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1351_
timestamp 1644511149
transform 1 0 4232 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1352_
timestamp 1644511149
transform 1 0 4600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1353_
timestamp 1644511149
transform 1 0 7728 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1354_
timestamp 1644511149
transform 1 0 6900 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1355_
timestamp 1644511149
transform 1 0 7728 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1356_
timestamp 1644511149
transform 1 0 6716 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1357_
timestamp 1644511149
transform 1 0 6624 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1358_
timestamp 1644511149
transform 1 0 41676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1359_
timestamp 1644511149
transform 1 0 7820 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _1360_
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1361_
timestamp 1644511149
transform 1 0 9660 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1362_
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1363_
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1364_
timestamp 1644511149
transform 1 0 12328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1365_
timestamp 1644511149
transform 1 0 9660 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1366_
timestamp 1644511149
transform 1 0 9844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1367_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1368_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1369_
timestamp 1644511149
transform 1 0 18676 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1370_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1371_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1372_
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1373_
timestamp 1644511149
transform 1 0 24748 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1644511149
transform 1 0 26036 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1375_
timestamp 1644511149
transform 1 0 25944 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1644511149
transform 1 0 32568 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1644511149
transform 1 0 26128 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1644511149
transform 1 0 26496 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1644511149
transform 1 0 27600 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1644511149
transform 1 0 27600 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1644511149
transform 1 0 30176 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1644511149
transform 1 0 33028 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1644511149
transform 1 0 35144 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1644511149
transform 1 0 37352 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1387_
timestamp 1644511149
transform 1 0 47932 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1644511149
transform 1 0 51520 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1644511149
transform 1 0 50784 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1644511149
transform 1 0 54648 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1644511149
transform 1 0 56304 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1644511149
transform 1 0 55936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1644511149
transform 1 0 53360 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1644511149
transform 1 0 50784 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1644511149
transform 1 0 50784 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1644511149
transform 1 0 46000 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1644511149
transform 1 0 37536 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1644511149
transform 1 0 35328 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1644511149
transform 1 0 22080 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1644511149
transform 1 0 13064 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1644511149
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1644511149
transform 1 0 27416 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1644511149
transform 1 0 18124 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1644511149
transform 1 0 18308 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1644511149
transform 1 0 19412 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1644511149
transform 1 0 17112 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1644511149
transform 1 0 20148 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1644511149
transform 1 0 20240 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1644511149
transform 1 0 23184 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1644511149
transform 1 0 20700 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1644511149
transform 1 0 23184 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1644511149
transform 1 0 19872 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1644511149
transform 1 0 22448 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1644511149
transform 1 0 19964 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1644511149
transform 1 0 20424 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1644511149
transform 1 0 23000 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1422_
timestamp 1644511149
transform 1 0 12696 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1423_
timestamp 1644511149
transform 1 0 11408 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1424_
timestamp 1644511149
transform 1 0 11684 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1425_
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1426_
timestamp 1644511149
transform 1 0 45632 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1427_
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1428_
timestamp 1644511149
transform 1 0 49588 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1429_
timestamp 1644511149
transform 1 0 47104 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1430_
timestamp 1644511149
transform 1 0 50048 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1431_
timestamp 1644511149
transform 1 0 51520 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1432_
timestamp 1644511149
transform 1 0 52992 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1433_
timestamp 1644511149
transform 1 0 53452 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1434_
timestamp 1644511149
transform 1 0 41216 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1435_
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1436_
timestamp 1644511149
transform 1 0 46460 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1437_
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1438_
timestamp 1644511149
transform 1 0 42136 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1439_
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1440_
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1441_
timestamp 1644511149
transform 1 0 45540 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1442_
timestamp 1644511149
transform 1 0 23644 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1443_
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1444_
timestamp 1644511149
transform 1 0 26220 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1445_
timestamp 1644511149
transform 1 0 27324 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1446_
timestamp 1644511149
transform 1 0 28244 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1447_
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1448_
timestamp 1644511149
transform 1 0 31004 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1449_
timestamp 1644511149
transform 1 0 33304 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1450_
timestamp 1644511149
transform 1 0 34776 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1451_
timestamp 1644511149
transform 1 0 37720 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1452_
timestamp 1644511149
transform 1 0 39744 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1453_
timestamp 1644511149
transform 1 0 37352 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1454_
timestamp 1644511149
transform 1 0 30176 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1455_
timestamp 1644511149
transform 1 0 34408 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1456_
timestamp 1644511149
transform 1 0 34684 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1457_
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1458_
timestamp 1644511149
transform 1 0 34500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1459_
timestamp 1644511149
transform 1 0 43332 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1460_
timestamp 1644511149
transform 1 0 37904 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1461_
timestamp 1644511149
transform 1 0 45172 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1462_
timestamp 1644511149
transform 1 0 9200 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1463_
timestamp 1644511149
transform 1 0 38088 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1464_
timestamp 1644511149
transform 1 0 41216 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1465_
timestamp 1644511149
transform 1 0 54004 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1466_
timestamp 1644511149
transform 1 0 43608 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1467_
timestamp 1644511149
transform 1 0 47840 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1468_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1469_
timestamp 1644511149
transform 1 0 43056 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1470_
timestamp 1644511149
transform 1 0 40756 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1471_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1472_
timestamp 1644511149
transform 1 0 9568 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1473_
timestamp 1644511149
transform 1 0 4048 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1474_
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1475_
timestamp 1644511149
transform 1 0 4600 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1476_
timestamp 1644511149
transform 1 0 4508 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1477_
timestamp 1644511149
transform 1 0 4048 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1478_
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1479_
timestamp 1644511149
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1480_
timestamp 1644511149
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1481_
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1482_
timestamp 1644511149
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1483_
timestamp 1644511149
transform 1 0 7084 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1484_
timestamp 1644511149
transform 1 0 6256 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1485_
timestamp 1644511149
transform 1 0 9476 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1486_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1487_
timestamp 1644511149
transform 1 0 15456 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1488_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1489_
timestamp 1644511149
transform 1 0 17112 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1490_
timestamp 1644511149
transform 1 0 16652 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1491_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1492_
timestamp 1644511149
transform 1 0 15272 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1493_
timestamp 1644511149
transform 1 0 9568 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1494_
timestamp 1644511149
transform 1 0 12420 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1495_
timestamp 1644511149
transform 1 0 9660 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1496_
timestamp 1644511149
transform 1 0 12512 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1497_
timestamp 1644511149
transform 1 0 14352 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1498_
timestamp 1644511149
transform 1 0 9568 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1499_
timestamp 1644511149
transform 1 0 5888 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1500_
timestamp 1644511149
transform 1 0 7360 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1501_
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1502_
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1503_
timestamp 1644511149
transform 1 0 6992 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1504_
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1505_
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1506_
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1507_
timestamp 1644511149
transform 1 0 1840 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1508_
timestamp 1644511149
transform 1 0 1932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1509_
timestamp 1644511149
transform 1 0 2024 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1510_
timestamp 1644511149
transform 1 0 1840 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1511_
timestamp 1644511149
transform 1 0 4048 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1512_
timestamp 1644511149
transform 1 0 6716 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1513_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1514_
timestamp 1644511149
transform 1 0 7176 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1515_
timestamp 1644511149
transform 1 0 4416 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1516_
timestamp 1644511149
transform 1 0 2576 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1517_
timestamp 1644511149
transform 1 0 2668 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1518_
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1519_
timestamp 1644511149
transform 1 0 1840 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1520_
timestamp 1644511149
transform 1 0 3772 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1521_
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1522_
timestamp 1644511149
transform 1 0 1840 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1523_
timestamp 1644511149
transform 1 0 4140 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1524_
timestamp 1644511149
transform 1 0 1840 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1525_
timestamp 1644511149
transform 1 0 4416 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1526_
timestamp 1644511149
transform 1 0 6808 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1527_
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1528_
timestamp 1644511149
transform 1 0 42596 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1529_
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1530_
timestamp 1644511149
transform 1 0 7360 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1531_
timestamp 1644511149
transform 1 0 10856 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1532_
timestamp 1644511149
transform 1 0 12144 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1533_
timestamp 1644511149
transform 1 0 9568 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1534__183 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1535__184
timestamp 1644511149
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1536__185
timestamp 1644511149
transform 1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1537__186
timestamp 1644511149
transform 1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1538__187
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1539__179
timestamp 1644511149
transform 1 0 41216 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1540__180
timestamp 1644511149
transform 1 0 48760 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1541__181
timestamp 1644511149
transform 1 0 4600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1542__182
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1543_
timestamp 1644511149
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1544_
timestamp 1644511149
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 33764 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 34868 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 36340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1644511149
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1644511149
transform 1 0 45356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1644511149
transform 1 0 46552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1644511149
transform 1 0 48024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1644511149
transform 1 0 50508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1644511149
transform 1 0 51428 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input21
timestamp 1644511149
transform 1 0 53912 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input22
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input23
timestamp 1644511149
transform 1 0 56764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input25
timestamp 1644511149
transform 1 0 57684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 56856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 21160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 28060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 3220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 3680 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 2944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 3496 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 2852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 2760 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 2668 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 2116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 3312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1644511149
transform 1 0 2668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  input56 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1472 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1644511149
transform 1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input58
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input61
timestamp 1644511149
transform 1 0 1564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1644511149
transform 1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input63
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input64
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input66
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input67
timestamp 1644511149
transform 1 0 1748 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input68
timestamp 1644511149
transform 1 0 1748 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input69
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1644511149
transform 1 0 1748 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input72
timestamp 1644511149
transform 1 0 1748 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1644511149
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input77
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input81
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input82
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1644511149
transform 1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 26956 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 56212 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform 1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1644511149
transform 1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1644511149
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1644511149
transform 1 0 30912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1644511149
transform 1 0 33396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1644511149
transform 1 0 36248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1644511149
transform 1 0 36156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1644511149
transform 1 0 38548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1644511149
transform 1 0 38272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1644511149
transform 1 0 41400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1644511149
transform 1 0 41216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1644511149
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1644511149
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1644511149
transform 1 0 45540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1644511149
transform 1 0 48300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1644511149
transform 1 0 48760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1644511149
transform 1 0 49956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1644511149
transform 1 0 51428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1644511149
transform 1 0 52900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1644511149
transform 1 0 54372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1644511149
transform 1 0 55844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1644511149
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1644511149
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1644511149
transform 1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1644511149
transform 1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1644511149
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1644511149
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1644511149
transform 1 0 2668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1644511149
transform 1 0 2116 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1644511149
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1644511149
transform 1 0 2852 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform 1 0 2668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1644511149
transform 1 0 2116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1644511149
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
<< labels >>
rlabel metal2 s 3698 41200 3754 42000 6 flash_csb
port 0 nsew signal tristate
rlabel metal2 s 11150 41200 11206 42000 6 flash_io0_read
port 1 nsew signal input
rlabel metal2 s 18694 41200 18750 42000 6 flash_io0_we
port 2 nsew signal tristate
rlabel metal2 s 26146 41200 26202 42000 6 flash_io0_write
port 3 nsew signal tristate
rlabel metal2 s 33690 41200 33746 42000 6 flash_io1_read
port 4 nsew signal input
rlabel metal2 s 41142 41200 41198 42000 6 flash_io1_we
port 5 nsew signal tristate
rlabel metal2 s 48686 41200 48742 42000 6 flash_io1_write
port 6 nsew signal tristate
rlabel metal2 s 56138 41200 56194 42000 6 flash_sck
port 7 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 sram_addr0[0]
port 8 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 sram_addr0[1]
port 9 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 sram_addr0[2]
port 10 nsew signal tristate
rlabel metal2 s 11334 0 11390 800 6 sram_addr0[3]
port 11 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 sram_addr0[4]
port 12 nsew signal tristate
rlabel metal2 s 16762 0 16818 800 6 sram_addr0[5]
port 13 nsew signal tristate
rlabel metal2 s 19154 0 19210 800 6 sram_addr0[6]
port 14 nsew signal tristate
rlabel metal2 s 21638 0 21694 800 6 sram_addr0[7]
port 15 nsew signal tristate
rlabel metal2 s 24030 0 24086 800 6 sram_addr0[8]
port 16 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 sram_addr1[0]
port 17 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 sram_addr1[1]
port 18 nsew signal tristate
rlabel metal2 s 8942 0 8998 800 6 sram_addr1[2]
port 19 nsew signal tristate
rlabel metal2 s 11886 0 11942 800 6 sram_addr1[3]
port 20 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 sram_addr1[4]
port 21 nsew signal tristate
rlabel metal2 s 17222 0 17278 800 6 sram_addr1[5]
port 22 nsew signal tristate
rlabel metal2 s 19706 0 19762 800 6 sram_addr1[6]
port 23 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 sram_addr1[7]
port 24 nsew signal tristate
rlabel metal2 s 24582 0 24638 800 6 sram_addr1[8]
port 25 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 sram_clk0
port 26 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 sram_clk1
port 27 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 sram_csb0
port 28 nsew signal tristate
rlabel metal2 s 1582 0 1638 800 6 sram_csb1
port 29 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 sram_din0[0]
port 30 nsew signal tristate
rlabel metal2 s 27986 0 28042 800 6 sram_din0[10]
port 31 nsew signal tristate
rlabel metal2 s 29458 0 29514 800 6 sram_din0[11]
port 32 nsew signal tristate
rlabel metal2 s 30838 0 30894 800 6 sram_din0[12]
port 33 nsew signal tristate
rlabel metal2 s 32310 0 32366 800 6 sram_din0[13]
port 34 nsew signal tristate
rlabel metal2 s 33782 0 33838 800 6 sram_din0[14]
port 35 nsew signal tristate
rlabel metal2 s 35254 0 35310 800 6 sram_din0[15]
port 36 nsew signal tristate
rlabel metal2 s 36726 0 36782 800 6 sram_din0[16]
port 37 nsew signal tristate
rlabel metal2 s 38198 0 38254 800 6 sram_din0[17]
port 38 nsew signal tristate
rlabel metal2 s 39670 0 39726 800 6 sram_din0[18]
port 39 nsew signal tristate
rlabel metal2 s 41142 0 41198 800 6 sram_din0[19]
port 40 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 sram_din0[1]
port 41 nsew signal tristate
rlabel metal2 s 42614 0 42670 800 6 sram_din0[20]
port 42 nsew signal tristate
rlabel metal2 s 44086 0 44142 800 6 sram_din0[21]
port 43 nsew signal tristate
rlabel metal2 s 45466 0 45522 800 6 sram_din0[22]
port 44 nsew signal tristate
rlabel metal2 s 46938 0 46994 800 6 sram_din0[23]
port 45 nsew signal tristate
rlabel metal2 s 48410 0 48466 800 6 sram_din0[24]
port 46 nsew signal tristate
rlabel metal2 s 49882 0 49938 800 6 sram_din0[25]
port 47 nsew signal tristate
rlabel metal2 s 51354 0 51410 800 6 sram_din0[26]
port 48 nsew signal tristate
rlabel metal2 s 52826 0 52882 800 6 sram_din0[27]
port 49 nsew signal tristate
rlabel metal2 s 54298 0 54354 800 6 sram_din0[28]
port 50 nsew signal tristate
rlabel metal2 s 55770 0 55826 800 6 sram_din0[29]
port 51 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 sram_din0[2]
port 52 nsew signal tristate
rlabel metal2 s 57242 0 57298 800 6 sram_din0[30]
port 53 nsew signal tristate
rlabel metal2 s 58714 0 58770 800 6 sram_din0[31]
port 54 nsew signal tristate
rlabel metal2 s 12346 0 12402 800 6 sram_din0[3]
port 55 nsew signal tristate
rlabel metal2 s 15290 0 15346 800 6 sram_din0[4]
port 56 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 sram_din0[5]
port 57 nsew signal tristate
rlabel metal2 s 20166 0 20222 800 6 sram_din0[6]
port 58 nsew signal tristate
rlabel metal2 s 22558 0 22614 800 6 sram_din0[7]
port 59 nsew signal tristate
rlabel metal2 s 25042 0 25098 800 6 sram_din0[8]
port 60 nsew signal tristate
rlabel metal2 s 26514 0 26570 800 6 sram_din0[9]
port 61 nsew signal tristate
rlabel metal2 s 4066 0 4122 800 6 sram_dout0[0]
port 62 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 sram_dout0[10]
port 63 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 sram_dout0[11]
port 64 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 sram_dout0[12]
port 65 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 sram_dout0[13]
port 66 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 sram_dout0[14]
port 67 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 sram_dout0[15]
port 68 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 sram_dout0[16]
port 69 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 sram_dout0[17]
port 70 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 sram_dout0[18]
port 71 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 sram_dout0[19]
port 72 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 sram_dout0[1]
port 73 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 sram_dout0[20]
port 74 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 sram_dout0[21]
port 75 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 sram_dout0[22]
port 76 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 sram_dout0[23]
port 77 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 sram_dout0[24]
port 78 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 sram_dout0[25]
port 79 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 sram_dout0[26]
port 80 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 sram_dout0[27]
port 81 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 sram_dout0[28]
port 82 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 sram_dout0[29]
port 83 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 sram_dout0[2]
port 84 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 sram_dout0[30]
port 85 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 sram_dout0[31]
port 86 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 sram_dout0[3]
port 87 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 sram_dout0[4]
port 88 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 sram_dout0[5]
port 89 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 sram_dout0[6]
port 90 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 sram_dout0[7]
port 91 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 sram_dout0[8]
port 92 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 sram_dout0[9]
port 93 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 sram_dout1[0]
port 94 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 sram_dout1[10]
port 95 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 sram_dout1[11]
port 96 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 sram_dout1[12]
port 97 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 sram_dout1[13]
port 98 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 sram_dout1[14]
port 99 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 sram_dout1[15]
port 100 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 sram_dout1[16]
port 101 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 sram_dout1[17]
port 102 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 sram_dout1[18]
port 103 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 sram_dout1[19]
port 104 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 sram_dout1[1]
port 105 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 sram_dout1[20]
port 106 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 sram_dout1[21]
port 107 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 sram_dout1[22]
port 108 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 sram_dout1[23]
port 109 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 sram_dout1[24]
port 110 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 sram_dout1[25]
port 111 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 sram_dout1[26]
port 112 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 sram_dout1[27]
port 113 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 sram_dout1[28]
port 114 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 sram_dout1[29]
port 115 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 sram_dout1[2]
port 116 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 sram_dout1[30]
port 117 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 sram_dout1[31]
port 118 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 sram_dout1[3]
port 119 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 sram_dout1[4]
port 120 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 sram_dout1[5]
port 121 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 sram_dout1[6]
port 122 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 sram_dout1[7]
port 123 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 sram_dout1[8]
port 124 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 sram_dout1[9]
port 125 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 sram_web0
port 126 nsew signal tristate
rlabel metal2 s 5078 0 5134 800 6 sram_wmask0[0]
port 127 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 sram_wmask0[1]
port 128 nsew signal tristate
rlabel metal2 s 10874 0 10930 800 6 sram_wmask0[2]
port 129 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 sram_wmask0[3]
port 130 nsew signal tristate
rlabel metal4 s 4208 2128 4528 39760 6 vccd1
port 131 nsew power input
rlabel metal4 s 34928 2128 35248 39760 6 vccd1
port 131 nsew power input
rlabel metal4 s 19568 2128 19888 39760 6 vssd1
port 132 nsew ground input
rlabel metal4 s 50288 2128 50608 39760 6 vssd1
port 132 nsew ground input
rlabel metal3 s 0 144 800 264 6 wb_ack_o
port 133 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 wb_adr_i[0]
port 134 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 wb_adr_i[10]
port 135 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_adr_i[11]
port 136 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wb_adr_i[12]
port 137 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 wb_adr_i[13]
port 138 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 wb_adr_i[14]
port 139 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 wb_adr_i[15]
port 140 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 wb_adr_i[16]
port 141 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wb_adr_i[17]
port 142 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 wb_adr_i[18]
port 143 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 wb_adr_i[19]
port 144 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wb_adr_i[1]
port 145 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wb_adr_i[20]
port 146 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 wb_adr_i[21]
port 147 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wb_adr_i[22]
port 148 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wb_adr_i[23]
port 149 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wb_adr_i[2]
port 150 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 wb_adr_i[3]
port 151 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 wb_adr_i[4]
port 152 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 wb_adr_i[5]
port 153 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 wb_adr_i[6]
port 154 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 wb_adr_i[7]
port 155 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 wb_adr_i[8]
port 156 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 wb_adr_i[9]
port 157 nsew signal input
rlabel metal3 s 0 552 800 672 6 wb_clk_i
port 158 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wb_cyc_i
port 159 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 wb_data_i[0]
port 160 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wb_data_i[10]
port 161 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wb_data_i[11]
port 162 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wb_data_i[12]
port 163 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wb_data_i[13]
port 164 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wb_data_i[14]
port 165 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 wb_data_i[15]
port 166 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wb_data_i[16]
port 167 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 wb_data_i[17]
port 168 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 wb_data_i[18]
port 169 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 wb_data_i[19]
port 170 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 wb_data_i[1]
port 171 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 wb_data_i[20]
port 172 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 wb_data_i[21]
port 173 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 wb_data_i[22]
port 174 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 wb_data_i[23]
port 175 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wb_data_i[24]
port 176 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 wb_data_i[25]
port 177 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 wb_data_i[26]
port 178 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 wb_data_i[27]
port 179 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 wb_data_i[28]
port 180 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 wb_data_i[29]
port 181 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 wb_data_i[2]
port 182 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 wb_data_i[30]
port 183 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 wb_data_i[31]
port 184 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 wb_data_i[3]
port 185 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 wb_data_i[4]
port 186 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 wb_data_i[5]
port 187 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 wb_data_i[6]
port 188 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 wb_data_i[7]
port 189 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wb_data_i[8]
port 190 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 wb_data_i[9]
port 191 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 wb_data_o[0]
port 192 nsew signal tristate
rlabel metal3 s 0 18504 800 18624 6 wb_data_o[10]
port 193 nsew signal tristate
rlabel metal3 s 0 19864 800 19984 6 wb_data_o[11]
port 194 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 wb_data_o[12]
port 195 nsew signal tristate
rlabel metal3 s 0 22312 800 22432 6 wb_data_o[13]
port 196 nsew signal tristate
rlabel metal3 s 0 23672 800 23792 6 wb_data_o[14]
port 197 nsew signal tristate
rlabel metal3 s 0 24896 800 25016 6 wb_data_o[15]
port 198 nsew signal tristate
rlabel metal3 s 0 26120 800 26240 6 wb_data_o[16]
port 199 nsew signal tristate
rlabel metal3 s 0 27344 800 27464 6 wb_data_o[17]
port 200 nsew signal tristate
rlabel metal3 s 0 28704 800 28824 6 wb_data_o[18]
port 201 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 wb_data_o[19]
port 202 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 wb_data_o[1]
port 203 nsew signal tristate
rlabel metal3 s 0 31152 800 31272 6 wb_data_o[20]
port 204 nsew signal tristate
rlabel metal3 s 0 32376 800 32496 6 wb_data_o[21]
port 205 nsew signal tristate
rlabel metal3 s 0 33736 800 33856 6 wb_data_o[22]
port 206 nsew signal tristate
rlabel metal3 s 0 34960 800 35080 6 wb_data_o[23]
port 207 nsew signal tristate
rlabel metal3 s 0 35776 800 35896 6 wb_data_o[24]
port 208 nsew signal tristate
rlabel metal3 s 0 36592 800 36712 6 wb_data_o[25]
port 209 nsew signal tristate
rlabel metal3 s 0 37544 800 37664 6 wb_data_o[26]
port 210 nsew signal tristate
rlabel metal3 s 0 38360 800 38480 6 wb_data_o[27]
port 211 nsew signal tristate
rlabel metal3 s 0 39176 800 39296 6 wb_data_o[28]
port 212 nsew signal tristate
rlabel metal3 s 0 39992 800 40112 6 wb_data_o[29]
port 213 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 wb_data_o[2]
port 214 nsew signal tristate
rlabel metal3 s 0 40808 800 40928 6 wb_data_o[30]
port 215 nsew signal tristate
rlabel metal3 s 0 41624 800 41744 6 wb_data_o[31]
port 216 nsew signal tristate
rlabel metal3 s 0 9256 800 9376 6 wb_data_o[3]
port 217 nsew signal tristate
rlabel metal3 s 0 11024 800 11144 6 wb_data_o[4]
port 218 nsew signal tristate
rlabel metal3 s 0 12248 800 12368 6 wb_data_o[5]
port 219 nsew signal tristate
rlabel metal3 s 0 13472 800 13592 6 wb_data_o[6]
port 220 nsew signal tristate
rlabel metal3 s 0 14832 800 14952 6 wb_data_o[7]
port 221 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 wb_data_o[8]
port 222 nsew signal tristate
rlabel metal3 s 0 17280 800 17400 6 wb_data_o[9]
port 223 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 wb_error_o
port 224 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 wb_rst_i
port 225 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 wb_sel_i[0]
port 226 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 wb_sel_i[1]
port 227 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 wb_sel_i[2]
port 228 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wb_sel_i[3]
port 229 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wb_stall_o
port 230 nsew signal tristate
rlabel metal3 s 0 2592 800 2712 6 wb_stb_i
port 231 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 wb_we_i
port 232 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 42000
<< end >>
