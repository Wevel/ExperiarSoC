magic
tech sky130A
magscale 1 2
timestamp 1683761239
<< obsli1 >>
rect 1104 2159 68816 97393
<< obsm1 >>
rect 934 892 69814 97424
<< metal2 >>
rect 4894 0 4950 800
rect 5446 0 5502 800
rect 5998 0 6054 800
rect 6550 0 6606 800
rect 7102 0 7158 800
rect 7654 0 7710 800
rect 8206 0 8262 800
rect 8758 0 8814 800
rect 9310 0 9366 800
rect 9862 0 9918 800
rect 10414 0 10470 800
rect 10966 0 11022 800
rect 11518 0 11574 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15382 0 15438 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17590 0 17646 800
rect 18142 0 18198 800
rect 18694 0 18750 800
rect 19246 0 19302 800
rect 19798 0 19854 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21454 0 21510 800
rect 22006 0 22062 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23662 0 23718 800
rect 24214 0 24270 800
rect 24766 0 24822 800
rect 25318 0 25374 800
rect 25870 0 25926 800
rect 26422 0 26478 800
rect 26974 0 27030 800
rect 27526 0 27582 800
rect 28078 0 28134 800
rect 28630 0 28686 800
rect 29182 0 29238 800
rect 29734 0 29790 800
rect 30286 0 30342 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31942 0 31998 800
rect 32494 0 32550 800
rect 33046 0 33102 800
rect 33598 0 33654 800
rect 34150 0 34206 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36358 0 36414 800
rect 36910 0 36966 800
rect 37462 0 37518 800
rect 38014 0 38070 800
rect 38566 0 38622 800
rect 39118 0 39174 800
rect 39670 0 39726 800
rect 40222 0 40278 800
rect 40774 0 40830 800
rect 41326 0 41382 800
rect 41878 0 41934 800
rect 42430 0 42486 800
rect 42982 0 43038 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44638 0 44694 800
rect 45190 0 45246 800
rect 45742 0 45798 800
rect 46294 0 46350 800
rect 46846 0 46902 800
rect 47398 0 47454 800
rect 47950 0 48006 800
rect 48502 0 48558 800
rect 49054 0 49110 800
rect 49606 0 49662 800
rect 50158 0 50214 800
rect 50710 0 50766 800
rect 51262 0 51318 800
rect 51814 0 51870 800
rect 52366 0 52422 800
rect 52918 0 52974 800
rect 53470 0 53526 800
rect 54022 0 54078 800
rect 54574 0 54630 800
rect 55126 0 55182 800
rect 55678 0 55734 800
rect 56230 0 56286 800
rect 56782 0 56838 800
rect 57334 0 57390 800
rect 57886 0 57942 800
rect 58438 0 58494 800
rect 58990 0 59046 800
rect 59542 0 59598 800
rect 60094 0 60150 800
rect 60646 0 60702 800
rect 61198 0 61254 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62854 0 62910 800
rect 63406 0 63462 800
rect 63958 0 64014 800
rect 64510 0 64566 800
rect 65062 0 65118 800
<< obsm2 >>
rect 938 856 69808 97413
rect 938 734 4838 856
rect 5006 734 5390 856
rect 5558 734 5942 856
rect 6110 734 6494 856
rect 6662 734 7046 856
rect 7214 734 7598 856
rect 7766 734 8150 856
rect 8318 734 8702 856
rect 8870 734 9254 856
rect 9422 734 9806 856
rect 9974 734 10358 856
rect 10526 734 10910 856
rect 11078 734 11462 856
rect 11630 734 12014 856
rect 12182 734 12566 856
rect 12734 734 13118 856
rect 13286 734 13670 856
rect 13838 734 14222 856
rect 14390 734 14774 856
rect 14942 734 15326 856
rect 15494 734 15878 856
rect 16046 734 16430 856
rect 16598 734 16982 856
rect 17150 734 17534 856
rect 17702 734 18086 856
rect 18254 734 18638 856
rect 18806 734 19190 856
rect 19358 734 19742 856
rect 19910 734 20294 856
rect 20462 734 20846 856
rect 21014 734 21398 856
rect 21566 734 21950 856
rect 22118 734 22502 856
rect 22670 734 23054 856
rect 23222 734 23606 856
rect 23774 734 24158 856
rect 24326 734 24710 856
rect 24878 734 25262 856
rect 25430 734 25814 856
rect 25982 734 26366 856
rect 26534 734 26918 856
rect 27086 734 27470 856
rect 27638 734 28022 856
rect 28190 734 28574 856
rect 28742 734 29126 856
rect 29294 734 29678 856
rect 29846 734 30230 856
rect 30398 734 30782 856
rect 30950 734 31334 856
rect 31502 734 31886 856
rect 32054 734 32438 856
rect 32606 734 32990 856
rect 33158 734 33542 856
rect 33710 734 34094 856
rect 34262 734 34646 856
rect 34814 734 35198 856
rect 35366 734 35750 856
rect 35918 734 36302 856
rect 36470 734 36854 856
rect 37022 734 37406 856
rect 37574 734 37958 856
rect 38126 734 38510 856
rect 38678 734 39062 856
rect 39230 734 39614 856
rect 39782 734 40166 856
rect 40334 734 40718 856
rect 40886 734 41270 856
rect 41438 734 41822 856
rect 41990 734 42374 856
rect 42542 734 42926 856
rect 43094 734 43478 856
rect 43646 734 44030 856
rect 44198 734 44582 856
rect 44750 734 45134 856
rect 45302 734 45686 856
rect 45854 734 46238 856
rect 46406 734 46790 856
rect 46958 734 47342 856
rect 47510 734 47894 856
rect 48062 734 48446 856
rect 48614 734 48998 856
rect 49166 734 49550 856
rect 49718 734 50102 856
rect 50270 734 50654 856
rect 50822 734 51206 856
rect 51374 734 51758 856
rect 51926 734 52310 856
rect 52478 734 52862 856
rect 53030 734 53414 856
rect 53582 734 53966 856
rect 54134 734 54518 856
rect 54686 734 55070 856
rect 55238 734 55622 856
rect 55790 734 56174 856
rect 56342 734 56726 856
rect 56894 734 57278 856
rect 57446 734 57830 856
rect 57998 734 58382 856
rect 58550 734 58934 856
rect 59102 734 59486 856
rect 59654 734 60038 856
rect 60206 734 60590 856
rect 60758 734 61142 856
rect 61310 734 61694 856
rect 61862 734 62246 856
rect 62414 734 62798 856
rect 62966 734 63350 856
rect 63518 734 63902 856
rect 64070 734 64454 856
rect 64622 734 65006 856
rect 65174 734 69808 856
<< metal3 >>
rect 0 88272 800 88392
rect 69200 88272 70000 88392
rect 0 87864 800 87984
rect 69200 87864 70000 87984
rect 0 87456 800 87576
rect 69200 87456 70000 87576
rect 0 87048 800 87168
rect 69200 87048 70000 87168
rect 0 86640 800 86760
rect 69200 86640 70000 86760
rect 0 86232 800 86352
rect 69200 86232 70000 86352
rect 0 85824 800 85944
rect 69200 85824 70000 85944
rect 0 85416 800 85536
rect 69200 85416 70000 85536
rect 0 85008 800 85128
rect 69200 85008 70000 85128
rect 0 84600 800 84720
rect 69200 84600 70000 84720
rect 0 84192 800 84312
rect 69200 84192 70000 84312
rect 0 83784 800 83904
rect 69200 83784 70000 83904
rect 0 83376 800 83496
rect 69200 83376 70000 83496
rect 0 82968 800 83088
rect 69200 82968 70000 83088
rect 0 82560 800 82680
rect 69200 82560 70000 82680
rect 0 82152 800 82272
rect 69200 82152 70000 82272
rect 0 81744 800 81864
rect 69200 81744 70000 81864
rect 0 81336 800 81456
rect 69200 81336 70000 81456
rect 0 80928 800 81048
rect 69200 80928 70000 81048
rect 0 80520 800 80640
rect 69200 80520 70000 80640
rect 0 80112 800 80232
rect 69200 80112 70000 80232
rect 0 79704 800 79824
rect 69200 79704 70000 79824
rect 0 79296 800 79416
rect 69200 79296 70000 79416
rect 0 78888 800 79008
rect 69200 78888 70000 79008
rect 0 78480 800 78600
rect 69200 78480 70000 78600
rect 0 78072 800 78192
rect 69200 78072 70000 78192
rect 0 77664 800 77784
rect 69200 77664 70000 77784
rect 0 77256 800 77376
rect 69200 77256 70000 77376
rect 0 76848 800 76968
rect 69200 76848 70000 76968
rect 0 76440 800 76560
rect 69200 76440 70000 76560
rect 0 76032 800 76152
rect 69200 76032 70000 76152
rect 0 75624 800 75744
rect 69200 75624 70000 75744
rect 0 75216 800 75336
rect 69200 75216 70000 75336
rect 0 74808 800 74928
rect 69200 74808 70000 74928
rect 0 74400 800 74520
rect 69200 74400 70000 74520
rect 0 73992 800 74112
rect 69200 73992 70000 74112
rect 0 73584 800 73704
rect 69200 73584 70000 73704
rect 0 73176 800 73296
rect 69200 73176 70000 73296
rect 0 72768 800 72888
rect 69200 72768 70000 72888
rect 0 72360 800 72480
rect 69200 72360 70000 72480
rect 0 71952 800 72072
rect 69200 71952 70000 72072
rect 0 71544 800 71664
rect 69200 71544 70000 71664
rect 0 71136 800 71256
rect 69200 71136 70000 71256
rect 0 70728 800 70848
rect 69200 70728 70000 70848
rect 0 70320 800 70440
rect 69200 70320 70000 70440
rect 0 69912 800 70032
rect 69200 69912 70000 70032
rect 0 69504 800 69624
rect 69200 69504 70000 69624
rect 0 69096 800 69216
rect 69200 69096 70000 69216
rect 0 68688 800 68808
rect 69200 68688 70000 68808
rect 0 68280 800 68400
rect 69200 68280 70000 68400
rect 0 67872 800 67992
rect 69200 67872 70000 67992
rect 0 67464 800 67584
rect 69200 67464 70000 67584
rect 0 67056 800 67176
rect 69200 67056 70000 67176
rect 0 66648 800 66768
rect 69200 66648 70000 66768
rect 0 66240 800 66360
rect 69200 66240 70000 66360
rect 0 65832 800 65952
rect 69200 65832 70000 65952
rect 0 65424 800 65544
rect 69200 65424 70000 65544
rect 0 65016 800 65136
rect 69200 65016 70000 65136
rect 0 64608 800 64728
rect 69200 64608 70000 64728
rect 0 64200 800 64320
rect 69200 64200 70000 64320
rect 0 63792 800 63912
rect 69200 63792 70000 63912
rect 0 63384 800 63504
rect 69200 63384 70000 63504
rect 0 62976 800 63096
rect 69200 62976 70000 63096
rect 0 62568 800 62688
rect 69200 62568 70000 62688
rect 0 62160 800 62280
rect 69200 62160 70000 62280
rect 0 61752 800 61872
rect 69200 61752 70000 61872
rect 0 61344 800 61464
rect 69200 61344 70000 61464
rect 0 60936 800 61056
rect 69200 60936 70000 61056
rect 0 60528 800 60648
rect 69200 60528 70000 60648
rect 0 60120 800 60240
rect 69200 60120 70000 60240
rect 0 59712 800 59832
rect 69200 59712 70000 59832
rect 0 59304 800 59424
rect 69200 59304 70000 59424
rect 0 58896 800 59016
rect 69200 58896 70000 59016
rect 0 58488 800 58608
rect 69200 58488 70000 58608
rect 0 58080 800 58200
rect 69200 58080 70000 58200
rect 0 57672 800 57792
rect 69200 57672 70000 57792
rect 0 57264 800 57384
rect 69200 57264 70000 57384
rect 0 56856 800 56976
rect 69200 56856 70000 56976
rect 0 56448 800 56568
rect 69200 56448 70000 56568
rect 0 56040 800 56160
rect 69200 56040 70000 56160
rect 0 55632 800 55752
rect 69200 55632 70000 55752
rect 0 55224 800 55344
rect 69200 55224 70000 55344
rect 0 54816 800 54936
rect 69200 54816 70000 54936
rect 0 54408 800 54528
rect 69200 54408 70000 54528
rect 0 54000 800 54120
rect 69200 54000 70000 54120
rect 0 53592 800 53712
rect 69200 53592 70000 53712
rect 0 53184 800 53304
rect 69200 53184 70000 53304
rect 0 52776 800 52896
rect 69200 52776 70000 52896
rect 0 52368 800 52488
rect 69200 52368 70000 52488
rect 0 51960 800 52080
rect 69200 51960 70000 52080
rect 0 51552 800 51672
rect 69200 51552 70000 51672
rect 0 51144 800 51264
rect 69200 51144 70000 51264
rect 0 50736 800 50856
rect 69200 50736 70000 50856
rect 0 50328 800 50448
rect 69200 50328 70000 50448
rect 0 49920 800 50040
rect 69200 49920 70000 50040
rect 0 49512 800 49632
rect 69200 49512 70000 49632
rect 0 49104 800 49224
rect 69200 49104 70000 49224
rect 0 48696 800 48816
rect 69200 48696 70000 48816
rect 0 48288 800 48408
rect 69200 48288 70000 48408
rect 0 47880 800 48000
rect 69200 47880 70000 48000
rect 0 47472 800 47592
rect 69200 47472 70000 47592
rect 0 47064 800 47184
rect 69200 47064 70000 47184
rect 0 46656 800 46776
rect 69200 46656 70000 46776
rect 0 46248 800 46368
rect 69200 46248 70000 46368
rect 0 45840 800 45960
rect 69200 45840 70000 45960
rect 0 45432 800 45552
rect 69200 45432 70000 45552
rect 0 45024 800 45144
rect 69200 45024 70000 45144
rect 0 44616 800 44736
rect 69200 44616 70000 44736
rect 0 44208 800 44328
rect 69200 44208 70000 44328
rect 0 43800 800 43920
rect 69200 43800 70000 43920
rect 0 43392 800 43512
rect 69200 43392 70000 43512
rect 0 42984 800 43104
rect 69200 42984 70000 43104
rect 0 42576 800 42696
rect 69200 42576 70000 42696
rect 0 42168 800 42288
rect 69200 42168 70000 42288
rect 0 41760 800 41880
rect 69200 41760 70000 41880
rect 0 41352 800 41472
rect 69200 41352 70000 41472
rect 0 40944 800 41064
rect 69200 40944 70000 41064
rect 0 40536 800 40656
rect 69200 40536 70000 40656
rect 0 40128 800 40248
rect 69200 40128 70000 40248
rect 0 39720 800 39840
rect 69200 39720 70000 39840
rect 0 39312 800 39432
rect 69200 39312 70000 39432
rect 0 38904 800 39024
rect 69200 38904 70000 39024
rect 0 38496 800 38616
rect 69200 38496 70000 38616
rect 0 38088 800 38208
rect 69200 38088 70000 38208
rect 0 37680 800 37800
rect 69200 37680 70000 37800
rect 0 37272 800 37392
rect 69200 37272 70000 37392
rect 0 36864 800 36984
rect 69200 36864 70000 36984
rect 0 36456 800 36576
rect 69200 36456 70000 36576
rect 0 36048 800 36168
rect 69200 36048 70000 36168
rect 0 35640 800 35760
rect 69200 35640 70000 35760
rect 0 35232 800 35352
rect 69200 35232 70000 35352
rect 0 34824 800 34944
rect 69200 34824 70000 34944
rect 0 34416 800 34536
rect 69200 34416 70000 34536
rect 0 34008 800 34128
rect 69200 34008 70000 34128
rect 0 33600 800 33720
rect 69200 33600 70000 33720
rect 0 33192 800 33312
rect 69200 33192 70000 33312
rect 0 32784 800 32904
rect 69200 32784 70000 32904
rect 0 32376 800 32496
rect 69200 32376 70000 32496
rect 0 31968 800 32088
rect 69200 31968 70000 32088
rect 0 31560 800 31680
rect 69200 31560 70000 31680
rect 0 31152 800 31272
rect 69200 31152 70000 31272
rect 0 30744 800 30864
rect 69200 30744 70000 30864
rect 0 30336 800 30456
rect 69200 30336 70000 30456
rect 0 29928 800 30048
rect 69200 29928 70000 30048
rect 0 29520 800 29640
rect 69200 29520 70000 29640
rect 0 29112 800 29232
rect 69200 29112 70000 29232
rect 0 28704 800 28824
rect 69200 28704 70000 28824
rect 0 28296 800 28416
rect 69200 28296 70000 28416
rect 0 27888 800 28008
rect 69200 27888 70000 28008
rect 0 27480 800 27600
rect 69200 27480 70000 27600
rect 0 27072 800 27192
rect 69200 27072 70000 27192
rect 0 26664 800 26784
rect 69200 26664 70000 26784
rect 0 26256 800 26376
rect 69200 26256 70000 26376
rect 0 25848 800 25968
rect 69200 25848 70000 25968
rect 0 25440 800 25560
rect 69200 25440 70000 25560
rect 0 25032 800 25152
rect 69200 25032 70000 25152
rect 0 24624 800 24744
rect 69200 24624 70000 24744
rect 0 24216 800 24336
rect 69200 24216 70000 24336
rect 0 23808 800 23928
rect 69200 23808 70000 23928
rect 0 23400 800 23520
rect 69200 23400 70000 23520
rect 0 22992 800 23112
rect 69200 22992 70000 23112
rect 0 22584 800 22704
rect 69200 22584 70000 22704
rect 0 22176 800 22296
rect 69200 22176 70000 22296
rect 0 21768 800 21888
rect 69200 21768 70000 21888
rect 0 21360 800 21480
rect 69200 21360 70000 21480
rect 0 20952 800 21072
rect 69200 20952 70000 21072
rect 0 20544 800 20664
rect 69200 20544 70000 20664
rect 0 20136 800 20256
rect 69200 20136 70000 20256
rect 0 19728 800 19848
rect 69200 19728 70000 19848
rect 0 19320 800 19440
rect 69200 19320 70000 19440
rect 0 18912 800 19032
rect 69200 18912 70000 19032
rect 0 18504 800 18624
rect 69200 18504 70000 18624
rect 0 18096 800 18216
rect 69200 18096 70000 18216
rect 0 17688 800 17808
rect 69200 17688 70000 17808
rect 0 17280 800 17400
rect 69200 17280 70000 17400
rect 0 16872 800 16992
rect 69200 16872 70000 16992
rect 0 16464 800 16584
rect 69200 16464 70000 16584
rect 0 16056 800 16176
rect 69200 16056 70000 16176
rect 0 15648 800 15768
rect 69200 15648 70000 15768
rect 0 15240 800 15360
rect 69200 15240 70000 15360
rect 0 14832 800 14952
rect 69200 14832 70000 14952
rect 0 14424 800 14544
rect 69200 14424 70000 14544
rect 0 14016 800 14136
rect 69200 14016 70000 14136
rect 0 13608 800 13728
rect 69200 13608 70000 13728
rect 0 13200 800 13320
rect 69200 13200 70000 13320
rect 0 12792 800 12912
rect 69200 12792 70000 12912
rect 0 12384 800 12504
rect 69200 12384 70000 12504
rect 0 11976 800 12096
rect 69200 11976 70000 12096
rect 0 11568 800 11688
rect 69200 11568 70000 11688
<< obsm3 >>
rect 800 88472 69200 97409
rect 880 88192 69120 88472
rect 800 88064 69200 88192
rect 880 87784 69120 88064
rect 800 87656 69200 87784
rect 880 87376 69120 87656
rect 800 87248 69200 87376
rect 880 86968 69120 87248
rect 800 86840 69200 86968
rect 880 86560 69120 86840
rect 800 86432 69200 86560
rect 880 86152 69120 86432
rect 800 86024 69200 86152
rect 880 85744 69120 86024
rect 800 85616 69200 85744
rect 880 85336 69120 85616
rect 800 85208 69200 85336
rect 880 84928 69120 85208
rect 800 84800 69200 84928
rect 880 84520 69120 84800
rect 800 84392 69200 84520
rect 880 84112 69120 84392
rect 800 83984 69200 84112
rect 880 83704 69120 83984
rect 800 83576 69200 83704
rect 880 83296 69120 83576
rect 800 83168 69200 83296
rect 880 82888 69120 83168
rect 800 82760 69200 82888
rect 880 82480 69120 82760
rect 800 82352 69200 82480
rect 880 82072 69120 82352
rect 800 81944 69200 82072
rect 880 81664 69120 81944
rect 800 81536 69200 81664
rect 880 81256 69120 81536
rect 800 81128 69200 81256
rect 880 80848 69120 81128
rect 800 80720 69200 80848
rect 880 80440 69120 80720
rect 800 80312 69200 80440
rect 880 80032 69120 80312
rect 800 79904 69200 80032
rect 880 79624 69120 79904
rect 800 79496 69200 79624
rect 880 79216 69120 79496
rect 800 79088 69200 79216
rect 880 78808 69120 79088
rect 800 78680 69200 78808
rect 880 78400 69120 78680
rect 800 78272 69200 78400
rect 880 77992 69120 78272
rect 800 77864 69200 77992
rect 880 77584 69120 77864
rect 800 77456 69200 77584
rect 880 77176 69120 77456
rect 800 77048 69200 77176
rect 880 76768 69120 77048
rect 800 76640 69200 76768
rect 880 76360 69120 76640
rect 800 76232 69200 76360
rect 880 75952 69120 76232
rect 800 75824 69200 75952
rect 880 75544 69120 75824
rect 800 75416 69200 75544
rect 880 75136 69120 75416
rect 800 75008 69200 75136
rect 880 74728 69120 75008
rect 800 74600 69200 74728
rect 880 74320 69120 74600
rect 800 74192 69200 74320
rect 880 73912 69120 74192
rect 800 73784 69200 73912
rect 880 73504 69120 73784
rect 800 73376 69200 73504
rect 880 73096 69120 73376
rect 800 72968 69200 73096
rect 880 72688 69120 72968
rect 800 72560 69200 72688
rect 880 72280 69120 72560
rect 800 72152 69200 72280
rect 880 71872 69120 72152
rect 800 71744 69200 71872
rect 880 71464 69120 71744
rect 800 71336 69200 71464
rect 880 71056 69120 71336
rect 800 70928 69200 71056
rect 880 70648 69120 70928
rect 800 70520 69200 70648
rect 880 70240 69120 70520
rect 800 70112 69200 70240
rect 880 69832 69120 70112
rect 800 69704 69200 69832
rect 880 69424 69120 69704
rect 800 69296 69200 69424
rect 880 69016 69120 69296
rect 800 68888 69200 69016
rect 880 68608 69120 68888
rect 800 68480 69200 68608
rect 880 68200 69120 68480
rect 800 68072 69200 68200
rect 880 67792 69120 68072
rect 800 67664 69200 67792
rect 880 67384 69120 67664
rect 800 67256 69200 67384
rect 880 66976 69120 67256
rect 800 66848 69200 66976
rect 880 66568 69120 66848
rect 800 66440 69200 66568
rect 880 66160 69120 66440
rect 800 66032 69200 66160
rect 880 65752 69120 66032
rect 800 65624 69200 65752
rect 880 65344 69120 65624
rect 800 65216 69200 65344
rect 880 64936 69120 65216
rect 800 64808 69200 64936
rect 880 64528 69120 64808
rect 800 64400 69200 64528
rect 880 64120 69120 64400
rect 800 63992 69200 64120
rect 880 63712 69120 63992
rect 800 63584 69200 63712
rect 880 63304 69120 63584
rect 800 63176 69200 63304
rect 880 62896 69120 63176
rect 800 62768 69200 62896
rect 880 62488 69120 62768
rect 800 62360 69200 62488
rect 880 62080 69120 62360
rect 800 61952 69200 62080
rect 880 61672 69120 61952
rect 800 61544 69200 61672
rect 880 61264 69120 61544
rect 800 61136 69200 61264
rect 880 60856 69120 61136
rect 800 60728 69200 60856
rect 880 60448 69120 60728
rect 800 60320 69200 60448
rect 880 60040 69120 60320
rect 800 59912 69200 60040
rect 880 59632 69120 59912
rect 800 59504 69200 59632
rect 880 59224 69120 59504
rect 800 59096 69200 59224
rect 880 58816 69120 59096
rect 800 58688 69200 58816
rect 880 58408 69120 58688
rect 800 58280 69200 58408
rect 880 58000 69120 58280
rect 800 57872 69200 58000
rect 880 57592 69120 57872
rect 800 57464 69200 57592
rect 880 57184 69120 57464
rect 800 57056 69200 57184
rect 880 56776 69120 57056
rect 800 56648 69200 56776
rect 880 56368 69120 56648
rect 800 56240 69200 56368
rect 880 55960 69120 56240
rect 800 55832 69200 55960
rect 880 55552 69120 55832
rect 800 55424 69200 55552
rect 880 55144 69120 55424
rect 800 55016 69200 55144
rect 880 54736 69120 55016
rect 800 54608 69200 54736
rect 880 54328 69120 54608
rect 800 54200 69200 54328
rect 880 53920 69120 54200
rect 800 53792 69200 53920
rect 880 53512 69120 53792
rect 800 53384 69200 53512
rect 880 53104 69120 53384
rect 800 52976 69200 53104
rect 880 52696 69120 52976
rect 800 52568 69200 52696
rect 880 52288 69120 52568
rect 800 52160 69200 52288
rect 880 51880 69120 52160
rect 800 51752 69200 51880
rect 880 51472 69120 51752
rect 800 51344 69200 51472
rect 880 51064 69120 51344
rect 800 50936 69200 51064
rect 880 50656 69120 50936
rect 800 50528 69200 50656
rect 880 50248 69120 50528
rect 800 50120 69200 50248
rect 880 49840 69120 50120
rect 800 49712 69200 49840
rect 880 49432 69120 49712
rect 800 49304 69200 49432
rect 880 49024 69120 49304
rect 800 48896 69200 49024
rect 880 48616 69120 48896
rect 800 48488 69200 48616
rect 880 48208 69120 48488
rect 800 48080 69200 48208
rect 880 47800 69120 48080
rect 800 47672 69200 47800
rect 880 47392 69120 47672
rect 800 47264 69200 47392
rect 880 46984 69120 47264
rect 800 46856 69200 46984
rect 880 46576 69120 46856
rect 800 46448 69200 46576
rect 880 46168 69120 46448
rect 800 46040 69200 46168
rect 880 45760 69120 46040
rect 800 45632 69200 45760
rect 880 45352 69120 45632
rect 800 45224 69200 45352
rect 880 44944 69120 45224
rect 800 44816 69200 44944
rect 880 44536 69120 44816
rect 800 44408 69200 44536
rect 880 44128 69120 44408
rect 800 44000 69200 44128
rect 880 43720 69120 44000
rect 800 43592 69200 43720
rect 880 43312 69120 43592
rect 800 43184 69200 43312
rect 880 42904 69120 43184
rect 800 42776 69200 42904
rect 880 42496 69120 42776
rect 800 42368 69200 42496
rect 880 42088 69120 42368
rect 800 41960 69200 42088
rect 880 41680 69120 41960
rect 800 41552 69200 41680
rect 880 41272 69120 41552
rect 800 41144 69200 41272
rect 880 40864 69120 41144
rect 800 40736 69200 40864
rect 880 40456 69120 40736
rect 800 40328 69200 40456
rect 880 40048 69120 40328
rect 800 39920 69200 40048
rect 880 39640 69120 39920
rect 800 39512 69200 39640
rect 880 39232 69120 39512
rect 800 39104 69200 39232
rect 880 38824 69120 39104
rect 800 38696 69200 38824
rect 880 38416 69120 38696
rect 800 38288 69200 38416
rect 880 38008 69120 38288
rect 800 37880 69200 38008
rect 880 37600 69120 37880
rect 800 37472 69200 37600
rect 880 37192 69120 37472
rect 800 37064 69200 37192
rect 880 36784 69120 37064
rect 800 36656 69200 36784
rect 880 36376 69120 36656
rect 800 36248 69200 36376
rect 880 35968 69120 36248
rect 800 35840 69200 35968
rect 880 35560 69120 35840
rect 800 35432 69200 35560
rect 880 35152 69120 35432
rect 800 35024 69200 35152
rect 880 34744 69120 35024
rect 800 34616 69200 34744
rect 880 34336 69120 34616
rect 800 34208 69200 34336
rect 880 33928 69120 34208
rect 800 33800 69200 33928
rect 880 33520 69120 33800
rect 800 33392 69200 33520
rect 880 33112 69120 33392
rect 800 32984 69200 33112
rect 880 32704 69120 32984
rect 800 32576 69200 32704
rect 880 32296 69120 32576
rect 800 32168 69200 32296
rect 880 31888 69120 32168
rect 800 31760 69200 31888
rect 880 31480 69120 31760
rect 800 31352 69200 31480
rect 880 31072 69120 31352
rect 800 30944 69200 31072
rect 880 30664 69120 30944
rect 800 30536 69200 30664
rect 880 30256 69120 30536
rect 800 30128 69200 30256
rect 880 29848 69120 30128
rect 800 29720 69200 29848
rect 880 29440 69120 29720
rect 800 29312 69200 29440
rect 880 29032 69120 29312
rect 800 28904 69200 29032
rect 880 28624 69120 28904
rect 800 28496 69200 28624
rect 880 28216 69120 28496
rect 800 28088 69200 28216
rect 880 27808 69120 28088
rect 800 27680 69200 27808
rect 880 27400 69120 27680
rect 800 27272 69200 27400
rect 880 26992 69120 27272
rect 800 26864 69200 26992
rect 880 26584 69120 26864
rect 800 26456 69200 26584
rect 880 26176 69120 26456
rect 800 26048 69200 26176
rect 880 25768 69120 26048
rect 800 25640 69200 25768
rect 880 25360 69120 25640
rect 800 25232 69200 25360
rect 880 24952 69120 25232
rect 800 24824 69200 24952
rect 880 24544 69120 24824
rect 800 24416 69200 24544
rect 880 24136 69120 24416
rect 800 24008 69200 24136
rect 880 23728 69120 24008
rect 800 23600 69200 23728
rect 880 23320 69120 23600
rect 800 23192 69200 23320
rect 880 22912 69120 23192
rect 800 22784 69200 22912
rect 880 22504 69120 22784
rect 800 22376 69200 22504
rect 880 22096 69120 22376
rect 800 21968 69200 22096
rect 880 21688 69120 21968
rect 800 21560 69200 21688
rect 880 21280 69120 21560
rect 800 21152 69200 21280
rect 880 20872 69120 21152
rect 800 20744 69200 20872
rect 880 20464 69120 20744
rect 800 20336 69200 20464
rect 880 20056 69120 20336
rect 800 19928 69200 20056
rect 880 19648 69120 19928
rect 800 19520 69200 19648
rect 880 19240 69120 19520
rect 800 19112 69200 19240
rect 880 18832 69120 19112
rect 800 18704 69200 18832
rect 880 18424 69120 18704
rect 800 18296 69200 18424
rect 880 18016 69120 18296
rect 800 17888 69200 18016
rect 880 17608 69120 17888
rect 800 17480 69200 17608
rect 880 17200 69120 17480
rect 800 17072 69200 17200
rect 880 16792 69120 17072
rect 800 16664 69200 16792
rect 880 16384 69120 16664
rect 800 16256 69200 16384
rect 880 15976 69120 16256
rect 800 15848 69200 15976
rect 880 15568 69120 15848
rect 800 15440 69200 15568
rect 880 15160 69120 15440
rect 800 15032 69200 15160
rect 880 14752 69120 15032
rect 800 14624 69200 14752
rect 880 14344 69120 14624
rect 800 14216 69200 14344
rect 880 13936 69120 14216
rect 800 13808 69200 13936
rect 880 13528 69120 13808
rect 800 13400 69200 13528
rect 880 13120 69120 13400
rect 800 12992 69200 13120
rect 880 12712 69120 12992
rect 800 12584 69200 12712
rect 880 12304 69120 12584
rect 800 12176 69200 12304
rect 880 11896 69120 12176
rect 800 11768 69200 11896
rect 880 11488 69120 11768
rect 800 2143 69200 11488
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
<< obsm4 >>
rect 7419 2483 19488 75445
rect 19968 2483 34848 75445
rect 35328 2483 50208 75445
rect 50688 2483 65568 75445
rect 66048 2483 66917 75445
<< labels >>
rlabel metal3 s 0 45840 800 45960 6 sram0_addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 sram0_addr0[1]
port 2 nsew signal output
rlabel metal3 s 0 46656 800 46776 6 sram0_addr0[2]
port 3 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 sram0_addr0[3]
port 4 nsew signal output
rlabel metal3 s 0 47472 800 47592 6 sram0_addr0[4]
port 5 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 sram0_addr0[5]
port 6 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 sram0_addr0[6]
port 7 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 sram0_addr0[7]
port 8 nsew signal output
rlabel metal3 s 0 49104 800 49224 6 sram0_addr0[8]
port 9 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 sram0_addr1[0]
port 10 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 sram0_addr1[1]
port 11 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 sram0_addr1[2]
port 12 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 sram0_addr1[3]
port 13 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 sram0_addr1[4]
port 14 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 sram0_addr1[5]
port 15 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 sram0_addr1[6]
port 16 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 sram0_addr1[7]
port 17 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 sram0_addr1[8]
port 18 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 sram0_clk0
port 19 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 sram0_clk1
port 20 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 sram0_csb0[0]
port 21 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 sram0_csb0[1]
port 22 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 sram0_csb1[0]
port 23 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 sram0_csb1[1]
port 24 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 sram0_din0[0]
port 25 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 sram0_din0[10]
port 26 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 sram0_din0[11]
port 27 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 sram0_din0[12]
port 28 nsew signal output
rlabel metal3 s 0 54816 800 54936 6 sram0_din0[13]
port 29 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 sram0_din0[14]
port 30 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 sram0_din0[15]
port 31 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 sram0_din0[16]
port 32 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 sram0_din0[17]
port 33 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 sram0_din0[18]
port 34 nsew signal output
rlabel metal3 s 0 57264 800 57384 6 sram0_din0[19]
port 35 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 sram0_din0[1]
port 36 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 sram0_din0[20]
port 37 nsew signal output
rlabel metal3 s 0 58080 800 58200 6 sram0_din0[21]
port 38 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 sram0_din0[22]
port 39 nsew signal output
rlabel metal3 s 0 58896 800 59016 6 sram0_din0[23]
port 40 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 sram0_din0[24]
port 41 nsew signal output
rlabel metal3 s 0 59712 800 59832 6 sram0_din0[25]
port 42 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 sram0_din0[26]
port 43 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 sram0_din0[27]
port 44 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 sram0_din0[28]
port 45 nsew signal output
rlabel metal3 s 0 61344 800 61464 6 sram0_din0[29]
port 46 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 sram0_din0[2]
port 47 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 sram0_din0[30]
port 48 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 sram0_din0[31]
port 49 nsew signal output
rlabel metal3 s 0 50736 800 50856 6 sram0_din0[3]
port 50 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 sram0_din0[4]
port 51 nsew signal output
rlabel metal3 s 0 51552 800 51672 6 sram0_din0[5]
port 52 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 sram0_din0[6]
port 53 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 sram0_din0[7]
port 54 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 sram0_din0[8]
port 55 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 sram0_din0[9]
port 56 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 sram0_dout0[0]
port 57 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 sram0_dout0[10]
port 58 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 sram0_dout0[11]
port 59 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 sram0_dout0[12]
port 60 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 sram0_dout0[13]
port 61 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 sram0_dout0[14]
port 62 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 sram0_dout0[15]
port 63 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 sram0_dout0[16]
port 64 nsew signal input
rlabel metal3 s 0 69504 800 69624 6 sram0_dout0[17]
port 65 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 sram0_dout0[18]
port 66 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 sram0_dout0[19]
port 67 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 sram0_dout0[1]
port 68 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 sram0_dout0[20]
port 69 nsew signal input
rlabel metal3 s 0 71136 800 71256 6 sram0_dout0[21]
port 70 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 sram0_dout0[22]
port 71 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 sram0_dout0[23]
port 72 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 sram0_dout0[24]
port 73 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 sram0_dout0[25]
port 74 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 sram0_dout0[26]
port 75 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 sram0_dout0[27]
port 76 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 sram0_dout0[28]
port 77 nsew signal input
rlabel metal3 s 0 74400 800 74520 6 sram0_dout0[29]
port 78 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 sram0_dout0[2]
port 79 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 sram0_dout0[30]
port 80 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 sram0_dout0[31]
port 81 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 sram0_dout0[32]
port 82 nsew signal input
rlabel metal3 s 0 76032 800 76152 6 sram0_dout0[33]
port 83 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 sram0_dout0[34]
port 84 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 sram0_dout0[35]
port 85 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 sram0_dout0[36]
port 86 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 sram0_dout0[37]
port 87 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 sram0_dout0[38]
port 88 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 sram0_dout0[39]
port 89 nsew signal input
rlabel metal3 s 0 63792 800 63912 6 sram0_dout0[3]
port 90 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 sram0_dout0[40]
port 91 nsew signal input
rlabel metal3 s 0 79296 800 79416 6 sram0_dout0[41]
port 92 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 sram0_dout0[42]
port 93 nsew signal input
rlabel metal3 s 0 80112 800 80232 6 sram0_dout0[43]
port 94 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 sram0_dout0[44]
port 95 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 sram0_dout0[45]
port 96 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 sram0_dout0[46]
port 97 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 sram0_dout0[47]
port 98 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 sram0_dout0[48]
port 99 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 sram0_dout0[49]
port 100 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 sram0_dout0[4]
port 101 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 sram0_dout0[50]
port 102 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 sram0_dout0[51]
port 103 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 sram0_dout0[52]
port 104 nsew signal input
rlabel metal3 s 0 84192 800 84312 6 sram0_dout0[53]
port 105 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 sram0_dout0[54]
port 106 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 sram0_dout0[55]
port 107 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 sram0_dout0[56]
port 108 nsew signal input
rlabel metal3 s 0 85824 800 85944 6 sram0_dout0[57]
port 109 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 sram0_dout0[58]
port 110 nsew signal input
rlabel metal3 s 0 86640 800 86760 6 sram0_dout0[59]
port 111 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 sram0_dout0[5]
port 112 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 sram0_dout0[60]
port 113 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 sram0_dout0[61]
port 114 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 sram0_dout0[62]
port 115 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 sram0_dout0[63]
port 116 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 sram0_dout0[6]
port 117 nsew signal input
rlabel metal3 s 0 65424 800 65544 6 sram0_dout0[7]
port 118 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 sram0_dout0[8]
port 119 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 sram0_dout0[9]
port 120 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 sram0_dout1[0]
port 121 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 sram0_dout1[10]
port 122 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 sram0_dout1[11]
port 123 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 sram0_dout1[12]
port 124 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 sram0_dout1[13]
port 125 nsew signal input
rlabel metal3 s 0 22176 800 22296 6 sram0_dout1[14]
port 126 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 sram0_dout1[15]
port 127 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 sram0_dout1[16]
port 128 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 sram0_dout1[17]
port 129 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 sram0_dout1[18]
port 130 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 sram0_dout1[19]
port 131 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 sram0_dout1[1]
port 132 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 sram0_dout1[20]
port 133 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 sram0_dout1[21]
port 134 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 sram0_dout1[22]
port 135 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 sram0_dout1[23]
port 136 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 sram0_dout1[24]
port 137 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 sram0_dout1[25]
port 138 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 sram0_dout1[26]
port 139 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 sram0_dout1[27]
port 140 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 sram0_dout1[28]
port 141 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 sram0_dout1[29]
port 142 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 sram0_dout1[2]
port 143 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 sram0_dout1[30]
port 144 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 sram0_dout1[31]
port 145 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 sram0_dout1[32]
port 146 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 sram0_dout1[33]
port 147 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 sram0_dout1[34]
port 148 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 sram0_dout1[35]
port 149 nsew signal input
rlabel metal3 s 0 31152 800 31272 6 sram0_dout1[36]
port 150 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 sram0_dout1[37]
port 151 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 sram0_dout1[38]
port 152 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 sram0_dout1[39]
port 153 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 sram0_dout1[3]
port 154 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 sram0_dout1[40]
port 155 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 sram0_dout1[41]
port 156 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 sram0_dout1[42]
port 157 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 sram0_dout1[43]
port 158 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 sram0_dout1[44]
port 159 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 sram0_dout1[45]
port 160 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 sram0_dout1[46]
port 161 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 sram0_dout1[47]
port 162 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 sram0_dout1[48]
port 163 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 sram0_dout1[49]
port 164 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 sram0_dout1[4]
port 165 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 sram0_dout1[50]
port 166 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 sram0_dout1[51]
port 167 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 sram0_dout1[52]
port 168 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 sram0_dout1[53]
port 169 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 sram0_dout1[54]
port 170 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 sram0_dout1[55]
port 171 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 sram0_dout1[56]
port 172 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 sram0_dout1[57]
port 173 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 sram0_dout1[58]
port 174 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 sram0_dout1[59]
port 175 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 sram0_dout1[5]
port 176 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 sram0_dout1[60]
port 177 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 sram0_dout1[61]
port 178 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 sram0_dout1[62]
port 179 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 sram0_dout1[63]
port 180 nsew signal input
rlabel metal3 s 0 18912 800 19032 6 sram0_dout1[6]
port 181 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 sram0_dout1[7]
port 182 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 sram0_dout1[8]
port 183 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 sram0_dout1[9]
port 184 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 sram0_web0
port 185 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 sram0_wmask0[0]
port 186 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 sram0_wmask0[1]
port 187 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 sram0_wmask0[2]
port 188 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 sram0_wmask0[3]
port 189 nsew signal output
rlabel metal3 s 69200 45840 70000 45960 6 sram1_addr0[0]
port 190 nsew signal output
rlabel metal3 s 69200 46248 70000 46368 6 sram1_addr0[1]
port 191 nsew signal output
rlabel metal3 s 69200 46656 70000 46776 6 sram1_addr0[2]
port 192 nsew signal output
rlabel metal3 s 69200 47064 70000 47184 6 sram1_addr0[3]
port 193 nsew signal output
rlabel metal3 s 69200 47472 70000 47592 6 sram1_addr0[4]
port 194 nsew signal output
rlabel metal3 s 69200 47880 70000 48000 6 sram1_addr0[5]
port 195 nsew signal output
rlabel metal3 s 69200 48288 70000 48408 6 sram1_addr0[6]
port 196 nsew signal output
rlabel metal3 s 69200 48696 70000 48816 6 sram1_addr0[7]
port 197 nsew signal output
rlabel metal3 s 69200 49104 70000 49224 6 sram1_addr0[8]
port 198 nsew signal output
rlabel metal3 s 69200 12792 70000 12912 6 sram1_addr1[0]
port 199 nsew signal output
rlabel metal3 s 69200 13200 70000 13320 6 sram1_addr1[1]
port 200 nsew signal output
rlabel metal3 s 69200 13608 70000 13728 6 sram1_addr1[2]
port 201 nsew signal output
rlabel metal3 s 69200 14016 70000 14136 6 sram1_addr1[3]
port 202 nsew signal output
rlabel metal3 s 69200 14424 70000 14544 6 sram1_addr1[4]
port 203 nsew signal output
rlabel metal3 s 69200 14832 70000 14952 6 sram1_addr1[5]
port 204 nsew signal output
rlabel metal3 s 69200 15240 70000 15360 6 sram1_addr1[6]
port 205 nsew signal output
rlabel metal3 s 69200 15648 70000 15768 6 sram1_addr1[7]
port 206 nsew signal output
rlabel metal3 s 69200 16056 70000 16176 6 sram1_addr1[8]
port 207 nsew signal output
rlabel metal3 s 69200 42576 70000 42696 6 sram1_clk0
port 208 nsew signal output
rlabel metal3 s 69200 11568 70000 11688 6 sram1_clk1
port 209 nsew signal output
rlabel metal3 s 69200 42984 70000 43104 6 sram1_csb0[0]
port 210 nsew signal output
rlabel metal3 s 69200 43392 70000 43512 6 sram1_csb0[1]
port 211 nsew signal output
rlabel metal3 s 69200 11976 70000 12096 6 sram1_csb1[0]
port 212 nsew signal output
rlabel metal3 s 69200 12384 70000 12504 6 sram1_csb1[1]
port 213 nsew signal output
rlabel metal3 s 69200 49512 70000 49632 6 sram1_din0[0]
port 214 nsew signal output
rlabel metal3 s 69200 53592 70000 53712 6 sram1_din0[10]
port 215 nsew signal output
rlabel metal3 s 69200 54000 70000 54120 6 sram1_din0[11]
port 216 nsew signal output
rlabel metal3 s 69200 54408 70000 54528 6 sram1_din0[12]
port 217 nsew signal output
rlabel metal3 s 69200 54816 70000 54936 6 sram1_din0[13]
port 218 nsew signal output
rlabel metal3 s 69200 55224 70000 55344 6 sram1_din0[14]
port 219 nsew signal output
rlabel metal3 s 69200 55632 70000 55752 6 sram1_din0[15]
port 220 nsew signal output
rlabel metal3 s 69200 56040 70000 56160 6 sram1_din0[16]
port 221 nsew signal output
rlabel metal3 s 69200 56448 70000 56568 6 sram1_din0[17]
port 222 nsew signal output
rlabel metal3 s 69200 56856 70000 56976 6 sram1_din0[18]
port 223 nsew signal output
rlabel metal3 s 69200 57264 70000 57384 6 sram1_din0[19]
port 224 nsew signal output
rlabel metal3 s 69200 49920 70000 50040 6 sram1_din0[1]
port 225 nsew signal output
rlabel metal3 s 69200 57672 70000 57792 6 sram1_din0[20]
port 226 nsew signal output
rlabel metal3 s 69200 58080 70000 58200 6 sram1_din0[21]
port 227 nsew signal output
rlabel metal3 s 69200 58488 70000 58608 6 sram1_din0[22]
port 228 nsew signal output
rlabel metal3 s 69200 58896 70000 59016 6 sram1_din0[23]
port 229 nsew signal output
rlabel metal3 s 69200 59304 70000 59424 6 sram1_din0[24]
port 230 nsew signal output
rlabel metal3 s 69200 59712 70000 59832 6 sram1_din0[25]
port 231 nsew signal output
rlabel metal3 s 69200 60120 70000 60240 6 sram1_din0[26]
port 232 nsew signal output
rlabel metal3 s 69200 60528 70000 60648 6 sram1_din0[27]
port 233 nsew signal output
rlabel metal3 s 69200 60936 70000 61056 6 sram1_din0[28]
port 234 nsew signal output
rlabel metal3 s 69200 61344 70000 61464 6 sram1_din0[29]
port 235 nsew signal output
rlabel metal3 s 69200 50328 70000 50448 6 sram1_din0[2]
port 236 nsew signal output
rlabel metal3 s 69200 61752 70000 61872 6 sram1_din0[30]
port 237 nsew signal output
rlabel metal3 s 69200 62160 70000 62280 6 sram1_din0[31]
port 238 nsew signal output
rlabel metal3 s 69200 50736 70000 50856 6 sram1_din0[3]
port 239 nsew signal output
rlabel metal3 s 69200 51144 70000 51264 6 sram1_din0[4]
port 240 nsew signal output
rlabel metal3 s 69200 51552 70000 51672 6 sram1_din0[5]
port 241 nsew signal output
rlabel metal3 s 69200 51960 70000 52080 6 sram1_din0[6]
port 242 nsew signal output
rlabel metal3 s 69200 52368 70000 52488 6 sram1_din0[7]
port 243 nsew signal output
rlabel metal3 s 69200 52776 70000 52896 6 sram1_din0[8]
port 244 nsew signal output
rlabel metal3 s 69200 53184 70000 53304 6 sram1_din0[9]
port 245 nsew signal output
rlabel metal3 s 69200 62568 70000 62688 6 sram1_dout0[0]
port 246 nsew signal input
rlabel metal3 s 69200 66648 70000 66768 6 sram1_dout0[10]
port 247 nsew signal input
rlabel metal3 s 69200 67056 70000 67176 6 sram1_dout0[11]
port 248 nsew signal input
rlabel metal3 s 69200 67464 70000 67584 6 sram1_dout0[12]
port 249 nsew signal input
rlabel metal3 s 69200 67872 70000 67992 6 sram1_dout0[13]
port 250 nsew signal input
rlabel metal3 s 69200 68280 70000 68400 6 sram1_dout0[14]
port 251 nsew signal input
rlabel metal3 s 69200 68688 70000 68808 6 sram1_dout0[15]
port 252 nsew signal input
rlabel metal3 s 69200 69096 70000 69216 6 sram1_dout0[16]
port 253 nsew signal input
rlabel metal3 s 69200 69504 70000 69624 6 sram1_dout0[17]
port 254 nsew signal input
rlabel metal3 s 69200 69912 70000 70032 6 sram1_dout0[18]
port 255 nsew signal input
rlabel metal3 s 69200 70320 70000 70440 6 sram1_dout0[19]
port 256 nsew signal input
rlabel metal3 s 69200 62976 70000 63096 6 sram1_dout0[1]
port 257 nsew signal input
rlabel metal3 s 69200 70728 70000 70848 6 sram1_dout0[20]
port 258 nsew signal input
rlabel metal3 s 69200 71136 70000 71256 6 sram1_dout0[21]
port 259 nsew signal input
rlabel metal3 s 69200 71544 70000 71664 6 sram1_dout0[22]
port 260 nsew signal input
rlabel metal3 s 69200 71952 70000 72072 6 sram1_dout0[23]
port 261 nsew signal input
rlabel metal3 s 69200 72360 70000 72480 6 sram1_dout0[24]
port 262 nsew signal input
rlabel metal3 s 69200 72768 70000 72888 6 sram1_dout0[25]
port 263 nsew signal input
rlabel metal3 s 69200 73176 70000 73296 6 sram1_dout0[26]
port 264 nsew signal input
rlabel metal3 s 69200 73584 70000 73704 6 sram1_dout0[27]
port 265 nsew signal input
rlabel metal3 s 69200 73992 70000 74112 6 sram1_dout0[28]
port 266 nsew signal input
rlabel metal3 s 69200 74400 70000 74520 6 sram1_dout0[29]
port 267 nsew signal input
rlabel metal3 s 69200 63384 70000 63504 6 sram1_dout0[2]
port 268 nsew signal input
rlabel metal3 s 69200 74808 70000 74928 6 sram1_dout0[30]
port 269 nsew signal input
rlabel metal3 s 69200 75216 70000 75336 6 sram1_dout0[31]
port 270 nsew signal input
rlabel metal3 s 69200 75624 70000 75744 6 sram1_dout0[32]
port 271 nsew signal input
rlabel metal3 s 69200 76032 70000 76152 6 sram1_dout0[33]
port 272 nsew signal input
rlabel metal3 s 69200 76440 70000 76560 6 sram1_dout0[34]
port 273 nsew signal input
rlabel metal3 s 69200 76848 70000 76968 6 sram1_dout0[35]
port 274 nsew signal input
rlabel metal3 s 69200 77256 70000 77376 6 sram1_dout0[36]
port 275 nsew signal input
rlabel metal3 s 69200 77664 70000 77784 6 sram1_dout0[37]
port 276 nsew signal input
rlabel metal3 s 69200 78072 70000 78192 6 sram1_dout0[38]
port 277 nsew signal input
rlabel metal3 s 69200 78480 70000 78600 6 sram1_dout0[39]
port 278 nsew signal input
rlabel metal3 s 69200 63792 70000 63912 6 sram1_dout0[3]
port 279 nsew signal input
rlabel metal3 s 69200 78888 70000 79008 6 sram1_dout0[40]
port 280 nsew signal input
rlabel metal3 s 69200 79296 70000 79416 6 sram1_dout0[41]
port 281 nsew signal input
rlabel metal3 s 69200 79704 70000 79824 6 sram1_dout0[42]
port 282 nsew signal input
rlabel metal3 s 69200 80112 70000 80232 6 sram1_dout0[43]
port 283 nsew signal input
rlabel metal3 s 69200 80520 70000 80640 6 sram1_dout0[44]
port 284 nsew signal input
rlabel metal3 s 69200 80928 70000 81048 6 sram1_dout0[45]
port 285 nsew signal input
rlabel metal3 s 69200 81336 70000 81456 6 sram1_dout0[46]
port 286 nsew signal input
rlabel metal3 s 69200 81744 70000 81864 6 sram1_dout0[47]
port 287 nsew signal input
rlabel metal3 s 69200 82152 70000 82272 6 sram1_dout0[48]
port 288 nsew signal input
rlabel metal3 s 69200 82560 70000 82680 6 sram1_dout0[49]
port 289 nsew signal input
rlabel metal3 s 69200 64200 70000 64320 6 sram1_dout0[4]
port 290 nsew signal input
rlabel metal3 s 69200 82968 70000 83088 6 sram1_dout0[50]
port 291 nsew signal input
rlabel metal3 s 69200 83376 70000 83496 6 sram1_dout0[51]
port 292 nsew signal input
rlabel metal3 s 69200 83784 70000 83904 6 sram1_dout0[52]
port 293 nsew signal input
rlabel metal3 s 69200 84192 70000 84312 6 sram1_dout0[53]
port 294 nsew signal input
rlabel metal3 s 69200 84600 70000 84720 6 sram1_dout0[54]
port 295 nsew signal input
rlabel metal3 s 69200 85008 70000 85128 6 sram1_dout0[55]
port 296 nsew signal input
rlabel metal3 s 69200 85416 70000 85536 6 sram1_dout0[56]
port 297 nsew signal input
rlabel metal3 s 69200 85824 70000 85944 6 sram1_dout0[57]
port 298 nsew signal input
rlabel metal3 s 69200 86232 70000 86352 6 sram1_dout0[58]
port 299 nsew signal input
rlabel metal3 s 69200 86640 70000 86760 6 sram1_dout0[59]
port 300 nsew signal input
rlabel metal3 s 69200 64608 70000 64728 6 sram1_dout0[5]
port 301 nsew signal input
rlabel metal3 s 69200 87048 70000 87168 6 sram1_dout0[60]
port 302 nsew signal input
rlabel metal3 s 69200 87456 70000 87576 6 sram1_dout0[61]
port 303 nsew signal input
rlabel metal3 s 69200 87864 70000 87984 6 sram1_dout0[62]
port 304 nsew signal input
rlabel metal3 s 69200 88272 70000 88392 6 sram1_dout0[63]
port 305 nsew signal input
rlabel metal3 s 69200 65016 70000 65136 6 sram1_dout0[6]
port 306 nsew signal input
rlabel metal3 s 69200 65424 70000 65544 6 sram1_dout0[7]
port 307 nsew signal input
rlabel metal3 s 69200 65832 70000 65952 6 sram1_dout0[8]
port 308 nsew signal input
rlabel metal3 s 69200 66240 70000 66360 6 sram1_dout0[9]
port 309 nsew signal input
rlabel metal3 s 69200 16464 70000 16584 6 sram1_dout1[0]
port 310 nsew signal input
rlabel metal3 s 69200 20544 70000 20664 6 sram1_dout1[10]
port 311 nsew signal input
rlabel metal3 s 69200 20952 70000 21072 6 sram1_dout1[11]
port 312 nsew signal input
rlabel metal3 s 69200 21360 70000 21480 6 sram1_dout1[12]
port 313 nsew signal input
rlabel metal3 s 69200 21768 70000 21888 6 sram1_dout1[13]
port 314 nsew signal input
rlabel metal3 s 69200 22176 70000 22296 6 sram1_dout1[14]
port 315 nsew signal input
rlabel metal3 s 69200 22584 70000 22704 6 sram1_dout1[15]
port 316 nsew signal input
rlabel metal3 s 69200 22992 70000 23112 6 sram1_dout1[16]
port 317 nsew signal input
rlabel metal3 s 69200 23400 70000 23520 6 sram1_dout1[17]
port 318 nsew signal input
rlabel metal3 s 69200 23808 70000 23928 6 sram1_dout1[18]
port 319 nsew signal input
rlabel metal3 s 69200 24216 70000 24336 6 sram1_dout1[19]
port 320 nsew signal input
rlabel metal3 s 69200 16872 70000 16992 6 sram1_dout1[1]
port 321 nsew signal input
rlabel metal3 s 69200 24624 70000 24744 6 sram1_dout1[20]
port 322 nsew signal input
rlabel metal3 s 69200 25032 70000 25152 6 sram1_dout1[21]
port 323 nsew signal input
rlabel metal3 s 69200 25440 70000 25560 6 sram1_dout1[22]
port 324 nsew signal input
rlabel metal3 s 69200 25848 70000 25968 6 sram1_dout1[23]
port 325 nsew signal input
rlabel metal3 s 69200 26256 70000 26376 6 sram1_dout1[24]
port 326 nsew signal input
rlabel metal3 s 69200 26664 70000 26784 6 sram1_dout1[25]
port 327 nsew signal input
rlabel metal3 s 69200 27072 70000 27192 6 sram1_dout1[26]
port 328 nsew signal input
rlabel metal3 s 69200 27480 70000 27600 6 sram1_dout1[27]
port 329 nsew signal input
rlabel metal3 s 69200 27888 70000 28008 6 sram1_dout1[28]
port 330 nsew signal input
rlabel metal3 s 69200 28296 70000 28416 6 sram1_dout1[29]
port 331 nsew signal input
rlabel metal3 s 69200 17280 70000 17400 6 sram1_dout1[2]
port 332 nsew signal input
rlabel metal3 s 69200 28704 70000 28824 6 sram1_dout1[30]
port 333 nsew signal input
rlabel metal3 s 69200 29112 70000 29232 6 sram1_dout1[31]
port 334 nsew signal input
rlabel metal3 s 69200 29520 70000 29640 6 sram1_dout1[32]
port 335 nsew signal input
rlabel metal3 s 69200 29928 70000 30048 6 sram1_dout1[33]
port 336 nsew signal input
rlabel metal3 s 69200 30336 70000 30456 6 sram1_dout1[34]
port 337 nsew signal input
rlabel metal3 s 69200 30744 70000 30864 6 sram1_dout1[35]
port 338 nsew signal input
rlabel metal3 s 69200 31152 70000 31272 6 sram1_dout1[36]
port 339 nsew signal input
rlabel metal3 s 69200 31560 70000 31680 6 sram1_dout1[37]
port 340 nsew signal input
rlabel metal3 s 69200 31968 70000 32088 6 sram1_dout1[38]
port 341 nsew signal input
rlabel metal3 s 69200 32376 70000 32496 6 sram1_dout1[39]
port 342 nsew signal input
rlabel metal3 s 69200 17688 70000 17808 6 sram1_dout1[3]
port 343 nsew signal input
rlabel metal3 s 69200 32784 70000 32904 6 sram1_dout1[40]
port 344 nsew signal input
rlabel metal3 s 69200 33192 70000 33312 6 sram1_dout1[41]
port 345 nsew signal input
rlabel metal3 s 69200 33600 70000 33720 6 sram1_dout1[42]
port 346 nsew signal input
rlabel metal3 s 69200 34008 70000 34128 6 sram1_dout1[43]
port 347 nsew signal input
rlabel metal3 s 69200 34416 70000 34536 6 sram1_dout1[44]
port 348 nsew signal input
rlabel metal3 s 69200 34824 70000 34944 6 sram1_dout1[45]
port 349 nsew signal input
rlabel metal3 s 69200 35232 70000 35352 6 sram1_dout1[46]
port 350 nsew signal input
rlabel metal3 s 69200 35640 70000 35760 6 sram1_dout1[47]
port 351 nsew signal input
rlabel metal3 s 69200 36048 70000 36168 6 sram1_dout1[48]
port 352 nsew signal input
rlabel metal3 s 69200 36456 70000 36576 6 sram1_dout1[49]
port 353 nsew signal input
rlabel metal3 s 69200 18096 70000 18216 6 sram1_dout1[4]
port 354 nsew signal input
rlabel metal3 s 69200 36864 70000 36984 6 sram1_dout1[50]
port 355 nsew signal input
rlabel metal3 s 69200 37272 70000 37392 6 sram1_dout1[51]
port 356 nsew signal input
rlabel metal3 s 69200 37680 70000 37800 6 sram1_dout1[52]
port 357 nsew signal input
rlabel metal3 s 69200 38088 70000 38208 6 sram1_dout1[53]
port 358 nsew signal input
rlabel metal3 s 69200 38496 70000 38616 6 sram1_dout1[54]
port 359 nsew signal input
rlabel metal3 s 69200 38904 70000 39024 6 sram1_dout1[55]
port 360 nsew signal input
rlabel metal3 s 69200 39312 70000 39432 6 sram1_dout1[56]
port 361 nsew signal input
rlabel metal3 s 69200 39720 70000 39840 6 sram1_dout1[57]
port 362 nsew signal input
rlabel metal3 s 69200 40128 70000 40248 6 sram1_dout1[58]
port 363 nsew signal input
rlabel metal3 s 69200 40536 70000 40656 6 sram1_dout1[59]
port 364 nsew signal input
rlabel metal3 s 69200 18504 70000 18624 6 sram1_dout1[5]
port 365 nsew signal input
rlabel metal3 s 69200 40944 70000 41064 6 sram1_dout1[60]
port 366 nsew signal input
rlabel metal3 s 69200 41352 70000 41472 6 sram1_dout1[61]
port 367 nsew signal input
rlabel metal3 s 69200 41760 70000 41880 6 sram1_dout1[62]
port 368 nsew signal input
rlabel metal3 s 69200 42168 70000 42288 6 sram1_dout1[63]
port 369 nsew signal input
rlabel metal3 s 69200 18912 70000 19032 6 sram1_dout1[6]
port 370 nsew signal input
rlabel metal3 s 69200 19320 70000 19440 6 sram1_dout1[7]
port 371 nsew signal input
rlabel metal3 s 69200 19728 70000 19848 6 sram1_dout1[8]
port 372 nsew signal input
rlabel metal3 s 69200 20136 70000 20256 6 sram1_dout1[9]
port 373 nsew signal input
rlabel metal3 s 69200 43800 70000 43920 6 sram1_web0
port 374 nsew signal output
rlabel metal3 s 69200 44208 70000 44328 6 sram1_wmask0[0]
port 375 nsew signal output
rlabel metal3 s 69200 44616 70000 44736 6 sram1_wmask0[1]
port 376 nsew signal output
rlabel metal3 s 69200 45024 70000 45144 6 sram1_wmask0[2]
port 377 nsew signal output
rlabel metal3 s 69200 45432 70000 45552 6 sram1_wmask0[3]
port 378 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 379 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 379 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 379 nsew power bidirectional
rlabel metal2 s 62302 0 62358 800 6 vga_b[0]
port 380 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 vga_b[1]
port 381 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 vga_g[0]
port 382 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 vga_g[1]
port 383 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 vga_hsync
port 384 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 vga_r[0]
port 385 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 vga_r[1]
port 386 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 vga_vsync
port 387 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 video_irq[0]
port 388 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 video_irq[1]
port 389 nsew signal output
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 390 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 390 nsew ground bidirectional
rlabel metal2 s 5998 0 6054 800 6 wb_ack_o
port 391 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wb_adr_i[0]
port 392 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wb_adr_i[10]
port 393 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wb_adr_i[11]
port 394 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wb_adr_i[12]
port 395 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wb_adr_i[13]
port 396 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wb_adr_i[14]
port 397 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wb_adr_i[15]
port 398 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wb_adr_i[16]
port 399 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wb_adr_i[17]
port 400 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wb_adr_i[18]
port 401 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wb_adr_i[19]
port 402 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wb_adr_i[1]
port 403 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wb_adr_i[20]
port 404 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wb_adr_i[21]
port 405 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 wb_adr_i[22]
port 406 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wb_adr_i[23]
port 407 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wb_adr_i[2]
port 408 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wb_adr_i[3]
port 409 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wb_adr_i[4]
port 410 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wb_adr_i[5]
port 411 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wb_adr_i[6]
port 412 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wb_adr_i[7]
port 413 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wb_adr_i[8]
port 414 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wb_adr_i[9]
port 415 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wb_clk_i
port 416 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wb_cyc_i
port 417 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wb_data_i[0]
port 418 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wb_data_i[10]
port 419 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wb_data_i[11]
port 420 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wb_data_i[12]
port 421 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wb_data_i[13]
port 422 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wb_data_i[14]
port 423 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wb_data_i[15]
port 424 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wb_data_i[16]
port 425 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wb_data_i[17]
port 426 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wb_data_i[18]
port 427 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wb_data_i[19]
port 428 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wb_data_i[1]
port 429 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 wb_data_i[20]
port 430 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 wb_data_i[21]
port 431 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wb_data_i[22]
port 432 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 wb_data_i[23]
port 433 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 wb_data_i[24]
port 434 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wb_data_i[25]
port 435 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 wb_data_i[26]
port 436 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wb_data_i[27]
port 437 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 wb_data_i[28]
port 438 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 wb_data_i[29]
port 439 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wb_data_i[2]
port 440 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wb_data_i[30]
port 441 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wb_data_i[31]
port 442 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wb_data_i[3]
port 443 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wb_data_i[4]
port 444 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wb_data_i[5]
port 445 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wb_data_i[6]
port 446 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wb_data_i[7]
port 447 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wb_data_i[8]
port 448 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wb_data_i[9]
port 449 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wb_data_o[0]
port 450 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wb_data_o[10]
port 451 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wb_data_o[11]
port 452 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wb_data_o[12]
port 453 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wb_data_o[13]
port 454 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wb_data_o[14]
port 455 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wb_data_o[15]
port 456 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 wb_data_o[16]
port 457 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 wb_data_o[17]
port 458 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 wb_data_o[18]
port 459 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 wb_data_o[19]
port 460 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wb_data_o[1]
port 461 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 wb_data_o[20]
port 462 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 wb_data_o[21]
port 463 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 wb_data_o[22]
port 464 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 wb_data_o[23]
port 465 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 wb_data_o[24]
port 466 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 wb_data_o[25]
port 467 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 wb_data_o[26]
port 468 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 wb_data_o[27]
port 469 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 wb_data_o[28]
port 470 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wb_data_o[29]
port 471 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wb_data_o[2]
port 472 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 wb_data_o[30]
port 473 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 wb_data_o[31]
port 474 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 wb_data_o[3]
port 475 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wb_data_o[4]
port 476 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wb_data_o[5]
port 477 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wb_data_o[6]
port 478 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 wb_data_o[7]
port 479 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wb_data_o[8]
port 480 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wb_data_o[9]
port 481 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wb_error_o
port 482 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 wb_rst_i
port 483 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wb_sel_i[0]
port 484 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wb_sel_i[1]
port 485 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wb_sel_i[2]
port 486 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wb_sel_i[3]
port 487 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wb_stall_o
port 488 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 wb_stb_i
port 489 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wb_we_i
port 490 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8284318
string GDS_FILE /mnt/f/WSL/ASIC/ExperiarSoC/openlane/Video/runs/23_05_11_00_24/results/signoff/Video.magic.gds
string GDS_START 1006448
<< end >>

