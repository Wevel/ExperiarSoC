magic
tech sky130A
magscale 1 2
timestamp 1651272818
<< viali >>
rect 38025 37417 38059 37451
rect 30021 37213 30055 37247
rect 37841 37213 37875 37247
rect 30205 37077 30239 37111
rect 29929 36873 29963 36907
rect 4077 36737 4111 36771
rect 12357 36737 12391 36771
rect 17509 36669 17543 36703
rect 17693 36669 17727 36703
rect 18061 36669 18095 36703
rect 24593 36669 24627 36703
rect 24777 36669 24811 36703
rect 25053 36669 25087 36703
rect 3157 36533 3191 36567
rect 3893 36533 3927 36567
rect 4721 36533 4755 36567
rect 8677 36533 8711 36567
rect 9137 36533 9171 36567
rect 12541 36533 12575 36567
rect 20545 36533 20579 36567
rect 26985 36533 27019 36567
rect 12541 36329 12575 36363
rect 17509 36329 17543 36363
rect 17969 36329 18003 36363
rect 25329 36329 25363 36363
rect 5273 36193 5307 36227
rect 8953 36193 8987 36227
rect 9781 36193 9815 36227
rect 11989 36193 12023 36227
rect 12633 36193 12667 36227
rect 19441 36193 19475 36227
rect 20913 36193 20947 36227
rect 22201 36193 22235 36227
rect 26617 36193 26651 36227
rect 27629 36193 27663 36227
rect 3249 36125 3283 36159
rect 3801 36125 3835 36159
rect 7665 36125 7699 36159
rect 12725 36125 12759 36159
rect 13369 36125 13403 36159
rect 14105 36125 14139 36159
rect 16037 36125 16071 36159
rect 18153 36125 18187 36159
rect 21741 36125 21775 36159
rect 24409 36125 24443 36159
rect 26157 36125 26191 36159
rect 3985 36057 4019 36091
rect 9137 36057 9171 36091
rect 12449 36057 12483 36091
rect 19625 36057 19659 36091
rect 21925 36057 21959 36091
rect 26801 36057 26835 36091
rect 12909 35989 12943 36023
rect 13553 35989 13587 36023
rect 19717 35785 19751 35819
rect 20821 35785 20855 35819
rect 5273 35717 5307 35751
rect 11989 35717 12023 35751
rect 12633 35717 12667 35751
rect 7573 35649 7607 35683
rect 10241 35649 10275 35683
rect 11713 35649 11747 35683
rect 12449 35649 12483 35683
rect 15945 35649 15979 35683
rect 16681 35649 16715 35683
rect 19533 35649 19567 35683
rect 20637 35649 20671 35683
rect 21833 35649 21867 35683
rect 30021 35649 30055 35683
rect 30288 35649 30322 35683
rect 32393 35649 32427 35683
rect 2973 35581 3007 35615
rect 3433 35581 3467 35615
rect 3617 35581 3651 35615
rect 7757 35581 7791 35615
rect 9413 35581 9447 35615
rect 11897 35581 11931 35615
rect 14197 35581 14231 35615
rect 16865 35581 16899 35615
rect 18245 35581 18279 35615
rect 23121 35581 23155 35615
rect 23305 35581 23339 35615
rect 23765 35581 23799 35615
rect 26433 35581 26467 35615
rect 26985 35581 27019 35615
rect 27169 35581 27203 35615
rect 28365 35581 28399 35615
rect 32137 35581 32171 35615
rect 16129 35513 16163 35547
rect 10057 35445 10091 35479
rect 11529 35445 11563 35479
rect 11989 35445 12023 35479
rect 22477 35445 22511 35479
rect 31401 35445 31435 35479
rect 33517 35445 33551 35479
rect 3249 35241 3283 35275
rect 3801 35241 3835 35275
rect 8033 35241 8067 35275
rect 12725 35241 12759 35275
rect 12909 35241 12943 35275
rect 16405 35241 16439 35275
rect 16865 35241 16899 35275
rect 17785 35241 17819 35275
rect 18245 35241 18279 35275
rect 26065 35241 26099 35275
rect 32137 35241 32171 35275
rect 6101 35105 6135 35139
rect 7021 35105 7055 35139
rect 9137 35105 9171 35139
rect 9321 35105 9355 35139
rect 10517 35105 10551 35139
rect 11989 35105 12023 35139
rect 13093 35105 13127 35139
rect 14105 35105 14139 35139
rect 15209 35105 15243 35139
rect 17969 35105 18003 35139
rect 21925 35105 21959 35139
rect 23765 35105 23799 35139
rect 24685 35105 24719 35139
rect 26709 35105 26743 35139
rect 28365 35105 28399 35139
rect 29561 35105 29595 35139
rect 3065 35037 3099 35071
rect 3985 35037 4019 35071
rect 6285 35037 6319 35071
rect 6745 35037 6779 35071
rect 8217 35037 8251 35071
rect 12265 35037 12299 35071
rect 12909 35037 12943 35071
rect 16589 35037 16623 35071
rect 16681 35037 16715 35071
rect 16865 35037 16899 35071
rect 18061 35037 18095 35071
rect 24409 35037 24443 35071
rect 25881 35037 25915 35071
rect 31953 35037 31987 35071
rect 4445 34969 4479 35003
rect 13185 34969 13219 35003
rect 14289 34969 14323 35003
rect 17785 34969 17819 35003
rect 22109 34969 22143 35003
rect 26893 34969 26927 35003
rect 29828 34969 29862 35003
rect 30941 34901 30975 34935
rect 6745 34697 6779 34731
rect 8125 34697 8159 34731
rect 11529 34697 11563 34731
rect 12449 34697 12483 34731
rect 13369 34697 13403 34731
rect 16681 34697 16715 34731
rect 18061 34697 18095 34731
rect 18981 34697 19015 34731
rect 21189 34697 21223 34731
rect 29837 34697 29871 34731
rect 30297 34697 30331 34731
rect 3341 34629 3375 34663
rect 7205 34629 7239 34663
rect 7665 34629 7699 34663
rect 3157 34561 3191 34595
rect 6929 34561 6963 34595
rect 7941 34561 7975 34595
rect 11713 34561 11747 34595
rect 11805 34561 11839 34595
rect 11989 34561 12023 34595
rect 12633 34561 12667 34595
rect 12909 34561 12943 34595
rect 13553 34561 13587 34595
rect 15945 34561 15979 34595
rect 16865 34561 16899 34595
rect 17141 34561 17175 34595
rect 17601 34561 17635 34595
rect 17893 34561 17927 34595
rect 18521 34561 18555 34595
rect 18797 34561 18831 34595
rect 21005 34561 21039 34595
rect 24317 34561 24351 34595
rect 29653 34561 29687 34595
rect 30481 34561 30515 34595
rect 32965 34561 32999 34595
rect 33232 34561 33266 34595
rect 4353 34493 4387 34527
rect 7113 34493 7147 34527
rect 7849 34493 7883 34527
rect 12725 34493 12759 34527
rect 16957 34493 16991 34527
rect 17693 34493 17727 34527
rect 18613 34493 18647 34527
rect 21833 34493 21867 34527
rect 22017 34493 22051 34527
rect 22293 34493 22327 34527
rect 24501 34493 24535 34527
rect 24777 34493 24811 34527
rect 2697 34357 2731 34391
rect 5641 34357 5675 34391
rect 7205 34357 7239 34391
rect 7665 34357 7699 34391
rect 11989 34357 12023 34391
rect 12633 34357 12667 34391
rect 16129 34357 16163 34391
rect 17141 34357 17175 34391
rect 17877 34357 17911 34391
rect 18521 34357 18555 34391
rect 19441 34357 19475 34391
rect 34345 34357 34379 34391
rect 7297 34153 7331 34187
rect 7757 34153 7791 34187
rect 13093 34153 13127 34187
rect 15669 34153 15703 34187
rect 17325 34153 17359 34187
rect 18245 34153 18279 34187
rect 19257 34153 19291 34187
rect 21833 34153 21867 34187
rect 23213 34153 23247 34187
rect 29745 34153 29779 34187
rect 30573 34153 30607 34187
rect 31861 34153 31895 34187
rect 32873 34153 32907 34187
rect 16313 34085 16347 34119
rect 18705 34085 18739 34119
rect 20913 34085 20947 34119
rect 4629 34017 4663 34051
rect 6285 34017 6319 34051
rect 7665 34017 7699 34051
rect 17417 34017 17451 34051
rect 18337 34017 18371 34051
rect 19349 34017 19383 34051
rect 24869 34017 24903 34051
rect 27629 34017 27663 34051
rect 30113 34017 30147 34051
rect 30941 34017 30975 34051
rect 31493 34017 31527 34051
rect 1409 33949 1443 33983
rect 2053 33949 2087 33983
rect 7481 33949 7515 33983
rect 11345 33949 11379 33983
rect 12357 33949 12391 33983
rect 12633 33949 12667 33983
rect 13277 33949 13311 33983
rect 15485 33949 15519 33983
rect 16129 33949 16163 33983
rect 17601 33949 17635 33983
rect 18521 33949 18555 33983
rect 19533 33949 19567 33983
rect 20729 33949 20763 33983
rect 24593 33949 24627 33983
rect 26065 33949 26099 33983
rect 26341 33949 26375 33983
rect 27353 33949 27387 33983
rect 29929 33949 29963 33983
rect 30757 33949 30791 33983
rect 31677 33949 31711 33983
rect 32689 33949 32723 33983
rect 37473 33949 37507 33983
rect 38117 33949 38151 33983
rect 6101 33881 6135 33915
rect 7757 33881 7791 33915
rect 17325 33881 17359 33915
rect 18245 33881 18279 33915
rect 19257 33881 19291 33915
rect 1593 33813 1627 33847
rect 11161 33813 11195 33847
rect 16773 33813 16807 33847
rect 17785 33813 17819 33847
rect 19717 33813 19751 33847
rect 37933 33813 37967 33847
rect 10425 33609 10459 33643
rect 16129 33609 16163 33643
rect 19809 33609 19843 33643
rect 32505 33609 32539 33643
rect 4629 33541 4663 33575
rect 8033 33541 8067 33575
rect 7757 33473 7791 33507
rect 10241 33473 10275 33507
rect 12449 33473 12483 33507
rect 16681 33473 16715 33507
rect 18613 33473 18647 33507
rect 18705 33473 18739 33507
rect 18889 33473 18923 33507
rect 19349 33473 19383 33507
rect 19625 33473 19659 33507
rect 32321 33473 32355 33507
rect 2789 33405 2823 33439
rect 2973 33405 3007 33439
rect 7941 33405 7975 33439
rect 12173 33405 12207 33439
rect 16957 33405 16991 33439
rect 19441 33405 19475 33439
rect 24501 33405 24535 33439
rect 24685 33405 24719 33439
rect 25605 33405 25639 33439
rect 32137 33405 32171 33439
rect 7113 33269 7147 33303
rect 7573 33269 7607 33303
rect 8033 33269 8067 33303
rect 10885 33269 10919 33303
rect 11621 33269 11655 33303
rect 18429 33269 18463 33303
rect 18613 33269 18647 33303
rect 19349 33269 19383 33303
rect 20269 33269 20303 33303
rect 27169 33269 27203 33303
rect 11897 33065 11931 33099
rect 17233 33065 17267 33099
rect 18337 33065 18371 33099
rect 24593 33065 24627 33099
rect 4077 32929 4111 32963
rect 11805 32929 11839 32963
rect 14933 32929 14967 32963
rect 15393 32929 15427 32963
rect 22845 32929 22879 32963
rect 25605 32929 25639 32963
rect 27445 32929 27479 32963
rect 3801 32861 3835 32895
rect 7757 32861 7791 32895
rect 11621 32861 11655 32895
rect 12449 32861 12483 32895
rect 14657 32861 14691 32895
rect 17049 32861 17083 32895
rect 18153 32861 18187 32895
rect 19257 32861 19291 32895
rect 22569 32861 22603 32895
rect 11897 32793 11931 32827
rect 27261 32793 27295 32827
rect 7573 32725 7607 32759
rect 11437 32725 11471 32759
rect 19901 32725 19935 32759
rect 25605 32521 25639 32555
rect 4721 32453 4755 32487
rect 7389 32453 7423 32487
rect 12633 32453 12667 32487
rect 1409 32385 1443 32419
rect 2053 32385 2087 32419
rect 7205 32385 7239 32419
rect 14289 32385 14323 32419
rect 17969 32385 18003 32419
rect 18705 32385 18739 32419
rect 23673 32385 23707 32419
rect 25421 32385 25455 32419
rect 2881 32317 2915 32351
rect 3065 32317 3099 32351
rect 9045 32317 9079 32351
rect 12449 32317 12483 32351
rect 18245 32317 18279 32351
rect 19349 32317 19383 32351
rect 23397 32317 23431 32351
rect 1593 32181 1627 32215
rect 5365 32181 5399 32215
rect 18889 32181 18923 32215
rect 2881 31977 2915 32011
rect 18521 31977 18555 32011
rect 24409 31977 24443 32011
rect 24593 31977 24627 32011
rect 37657 31909 37691 31943
rect 5273 31841 5307 31875
rect 5825 31841 5859 31875
rect 6929 31841 6963 31875
rect 11529 31841 11563 31875
rect 16589 31841 16623 31875
rect 30205 31841 30239 31875
rect 32413 31841 32447 31875
rect 33609 31841 33643 31875
rect 7205 31773 7239 31807
rect 11805 31773 11839 31807
rect 12817 31773 12851 31807
rect 14105 31773 14139 31807
rect 15669 31773 15703 31807
rect 16129 31773 16163 31807
rect 18613 31773 18647 31807
rect 19441 31773 19475 31807
rect 24593 31773 24627 31807
rect 24685 31773 24719 31807
rect 36277 31773 36311 31807
rect 5641 31705 5675 31739
rect 16313 31705 16347 31739
rect 24869 31705 24903 31739
rect 29929 31705 29963 31739
rect 32137 31705 32171 31739
rect 33333 31705 33367 31739
rect 36522 31705 36556 31739
rect 13001 31637 13035 31671
rect 23765 31637 23799 31671
rect 25421 31637 25455 31671
rect 29561 31637 29595 31671
rect 30021 31637 30055 31671
rect 30849 31637 30883 31671
rect 31769 31637 31803 31671
rect 32229 31637 32263 31671
rect 32965 31637 32999 31671
rect 33425 31637 33459 31671
rect 3709 31433 3743 31467
rect 22293 31433 22327 31467
rect 26065 31433 26099 31467
rect 31585 31433 31619 31467
rect 32505 31433 32539 31467
rect 32873 31433 32907 31467
rect 34529 31433 34563 31467
rect 2513 31365 2547 31399
rect 9137 31365 9171 31399
rect 10977 31365 11011 31399
rect 11897 31365 11931 31399
rect 13001 31365 13035 31399
rect 14657 31365 14691 31399
rect 17049 31365 17083 31399
rect 18061 31365 18095 31399
rect 19717 31365 19751 31399
rect 30573 31365 30607 31399
rect 31217 31365 31251 31399
rect 35510 31365 35544 31399
rect 1409 31297 1443 31331
rect 3893 31297 3927 31331
rect 4537 31297 4571 31331
rect 5549 31297 5583 31331
rect 12173 31297 12207 31331
rect 17233 31297 17267 31331
rect 19901 31297 19935 31331
rect 21833 31297 21867 31331
rect 22109 31297 22143 31331
rect 25605 31297 25639 31331
rect 25881 31297 25915 31331
rect 29561 31297 29595 31331
rect 31033 31297 31067 31331
rect 31309 31297 31343 31331
rect 31401 31297 31435 31331
rect 34345 31297 34379 31331
rect 2881 31229 2915 31263
rect 5825 31229 5859 31263
rect 6837 31229 6871 31263
rect 7297 31229 7331 31263
rect 7481 31229 7515 31263
rect 12081 31229 12115 31263
rect 12817 31229 12851 31263
rect 21925 31229 21959 31263
rect 23305 31229 23339 31263
rect 23489 31229 23523 31263
rect 23765 31229 23799 31263
rect 25697 31229 25731 31263
rect 29653 31229 29687 31263
rect 29837 31229 29871 31263
rect 32965 31229 32999 31263
rect 33149 31229 33183 31263
rect 35265 31229 35299 31263
rect 1593 31161 1627 31195
rect 2678 31093 2712 31127
rect 2789 31093 2823 31127
rect 3157 31093 3191 31127
rect 4353 31093 4387 31127
rect 11989 31093 12023 31127
rect 12357 31093 12391 31127
rect 21833 31093 21867 31127
rect 25605 31093 25639 31127
rect 29193 31093 29227 31127
rect 36645 31093 36679 31127
rect 7481 30889 7515 30923
rect 8401 30889 8435 30923
rect 9413 30889 9447 30923
rect 9873 30889 9907 30923
rect 10333 30889 10367 30923
rect 15209 30889 15243 30923
rect 19441 30889 19475 30923
rect 20913 30889 20947 30923
rect 21649 30889 21683 30923
rect 22017 30889 22051 30923
rect 22937 30889 22971 30923
rect 23397 30889 23431 30923
rect 24409 30889 24443 30923
rect 24869 30889 24903 30923
rect 29009 30889 29043 30923
rect 29561 30889 29595 30923
rect 30757 30889 30791 30923
rect 31953 30889 31987 30923
rect 33057 30889 33091 30923
rect 35633 30889 35667 30923
rect 1409 30821 1443 30855
rect 7941 30821 7975 30855
rect 8953 30821 8987 30855
rect 19257 30821 19291 30855
rect 21097 30821 21131 30855
rect 3985 30753 4019 30787
rect 4261 30753 4295 30787
rect 10241 30753 10275 30787
rect 11345 30753 11379 30787
rect 14749 30753 14783 30787
rect 17693 30753 17727 30787
rect 17969 30753 18003 30787
rect 18705 30753 18739 30787
rect 20729 30753 20763 30787
rect 21649 30753 21683 30787
rect 24501 30753 24535 30787
rect 30205 30753 30239 30787
rect 31309 30753 31343 30787
rect 33701 30753 33735 30787
rect 3249 30685 3283 30719
rect 3801 30685 3835 30719
rect 7297 30685 7331 30719
rect 8125 30685 8159 30719
rect 8217 30685 8251 30719
rect 9137 30685 9171 30719
rect 9229 30685 9263 30719
rect 10064 30685 10098 30719
rect 11161 30685 11195 30719
rect 15393 30685 15427 30719
rect 19441 30685 19475 30719
rect 19533 30685 19567 30719
rect 20913 30685 20947 30719
rect 21833 30685 21867 30719
rect 22753 30685 22787 30719
rect 24685 30685 24719 30719
rect 28457 30685 28491 30719
rect 28641 30685 28675 30719
rect 28825 30685 28859 30719
rect 29929 30685 29963 30719
rect 31217 30685 31251 30719
rect 32137 30685 32171 30719
rect 32321 30685 32355 30719
rect 32505 30685 32539 30719
rect 33517 30685 33551 30719
rect 35449 30685 35483 30719
rect 8401 30617 8435 30651
rect 9413 30617 9447 30651
rect 10333 30617 10367 30651
rect 13001 30617 13035 30651
rect 14565 30617 14599 30651
rect 18521 30617 18555 30651
rect 19717 30617 19751 30651
rect 20637 30617 20671 30651
rect 21557 30617 21591 30651
rect 24409 30617 24443 30651
rect 25329 30617 25363 30651
rect 28733 30617 28767 30651
rect 32229 30617 32263 30651
rect 16681 30549 16715 30583
rect 27997 30549 28031 30583
rect 30021 30549 30055 30583
rect 31125 30549 31159 30583
rect 33425 30549 33459 30583
rect 3893 30345 3927 30379
rect 4813 30345 4847 30379
rect 4353 30277 4387 30311
rect 5273 30277 5307 30311
rect 11989 30277 12023 30311
rect 13921 30277 13955 30311
rect 19257 30277 19291 30311
rect 29285 30277 29319 30311
rect 32505 30277 32539 30311
rect 4077 30209 4111 30243
rect 4997 30209 5031 30243
rect 10977 30209 11011 30243
rect 12265 30209 12299 30243
rect 13369 30209 13403 30243
rect 14105 30209 14139 30243
rect 18061 30209 18095 30243
rect 18981 30209 19015 30243
rect 20453 30209 20487 30243
rect 22017 30209 22051 30243
rect 29101 30209 29135 30243
rect 29377 30209 29411 30243
rect 29469 30209 29503 30243
rect 32321 30209 32355 30243
rect 35521 30209 35555 30243
rect 4169 30141 4203 30175
rect 5089 30141 5123 30175
rect 8217 30141 8251 30175
rect 9137 30141 9171 30175
rect 9321 30141 9355 30175
rect 12173 30141 12207 30175
rect 18337 30141 18371 30175
rect 19165 30141 19199 30175
rect 22661 30141 22695 30175
rect 22845 30141 22879 30175
rect 23673 30141 23707 30175
rect 30757 30141 30791 30175
rect 31033 30141 31067 30175
rect 32137 30141 32171 30175
rect 35265 30141 35299 30175
rect 12449 30073 12483 30107
rect 18797 30073 18831 30107
rect 20637 30073 20671 30107
rect 22201 30073 22235 30107
rect 31493 30073 31527 30107
rect 4353 30005 4387 30039
rect 5273 30005 5307 30039
rect 11989 30005 12023 30039
rect 13277 30005 13311 30039
rect 14841 30005 14875 30039
rect 18981 30005 19015 30039
rect 19809 30005 19843 30039
rect 28641 30005 28675 30039
rect 29653 30005 29687 30039
rect 36645 30005 36679 30039
rect 38117 30005 38151 30039
rect 1593 29801 1627 29835
rect 3893 29801 3927 29835
rect 4353 29801 4387 29835
rect 7665 29801 7699 29835
rect 9505 29801 9539 29835
rect 11805 29801 11839 29835
rect 21649 29801 21683 29835
rect 21833 29801 21867 29835
rect 22293 29801 22327 29835
rect 22753 29801 22787 29835
rect 30665 29801 30699 29835
rect 35081 29801 35115 29835
rect 23213 29733 23247 29767
rect 32321 29733 32355 29767
rect 4261 29665 4295 29699
rect 12541 29665 12575 29699
rect 15669 29665 15703 29699
rect 17785 29665 17819 29699
rect 21557 29665 21591 29699
rect 22385 29665 22419 29699
rect 28549 29665 28583 29699
rect 29009 29665 29043 29699
rect 31861 29665 31895 29699
rect 36737 29665 36771 29699
rect 37841 29665 37875 29699
rect 37933 29665 37967 29699
rect 1409 29597 1443 29631
rect 2053 29597 2087 29631
rect 4077 29597 4111 29631
rect 4353 29597 4387 29631
rect 12265 29597 12299 29631
rect 15945 29597 15979 29631
rect 18061 29597 18095 29631
rect 20545 29597 20579 29631
rect 21649 29597 21683 29631
rect 22569 29597 22603 29631
rect 34897 29597 34931 29631
rect 36553 29597 36587 29631
rect 36645 29597 36679 29631
rect 37749 29597 37783 29631
rect 9413 29529 9447 29563
rect 21373 29529 21407 29563
rect 22293 29529 22327 29563
rect 28825 29529 28859 29563
rect 30757 29529 30791 29563
rect 14105 29461 14139 29495
rect 15209 29461 15243 29495
rect 20729 29461 20763 29495
rect 29745 29461 29779 29495
rect 36185 29461 36219 29495
rect 37381 29461 37415 29495
rect 17141 29257 17175 29291
rect 18153 29257 18187 29291
rect 20269 29257 20303 29291
rect 30481 29257 30515 29291
rect 30205 29189 30239 29223
rect 31309 29189 31343 29223
rect 15025 29121 15059 29155
rect 15117 29121 15151 29155
rect 15301 29121 15335 29155
rect 15761 29121 15795 29155
rect 17233 29121 17267 29155
rect 18245 29121 18279 29155
rect 19073 29121 19107 29155
rect 20085 29121 20119 29155
rect 23489 29121 23523 29155
rect 24133 29121 24167 29155
rect 29929 29121 29963 29155
rect 30113 29121 30147 29155
rect 30297 29121 30331 29155
rect 3065 29053 3099 29087
rect 3525 29053 3559 29087
rect 3709 29053 3743 29087
rect 4169 29053 4203 29087
rect 13001 29053 13035 29087
rect 13829 29053 13863 29087
rect 14013 29053 14047 29087
rect 18797 29053 18831 29087
rect 28825 29053 28859 29087
rect 29101 29053 29135 29087
rect 29285 29053 29319 29087
rect 11713 28985 11747 29019
rect 15945 28985 15979 29019
rect 23029 28985 23063 29019
rect 24317 28985 24351 29019
rect 31493 28985 31527 29019
rect 8677 28917 8711 28951
rect 9229 28917 9263 28951
rect 14841 28917 14875 28951
rect 15301 28917 15335 28951
rect 20729 28917 20763 28951
rect 23673 28917 23707 28951
rect 3249 28713 3283 28747
rect 4445 28713 4479 28747
rect 15853 28713 15887 28747
rect 24409 28713 24443 28747
rect 30297 28713 30331 28747
rect 31125 28713 31159 28747
rect 33609 28713 33643 28747
rect 3985 28645 4019 28679
rect 4353 28577 4387 28611
rect 8953 28577 8987 28611
rect 9781 28577 9815 28611
rect 13001 28577 13035 28611
rect 14657 28577 14691 28611
rect 14933 28577 14967 28611
rect 15669 28577 15703 28611
rect 23305 28577 23339 28611
rect 24501 28577 24535 28611
rect 29745 28577 29779 28611
rect 1409 28509 1443 28543
rect 2605 28509 2639 28543
rect 3065 28509 3099 28543
rect 4169 28509 4203 28543
rect 4445 28509 4479 28543
rect 5733 28509 5767 28543
rect 13277 28509 13311 28543
rect 15853 28509 15887 28543
rect 23029 28509 23063 28543
rect 24685 28509 24719 28543
rect 25513 28509 25547 28543
rect 29929 28509 29963 28543
rect 5549 28441 5583 28475
rect 9137 28441 9171 28475
rect 15577 28441 15611 28475
rect 24409 28441 24443 28475
rect 33701 28441 33735 28475
rect 1593 28373 1627 28407
rect 4997 28373 5031 28407
rect 16037 28373 16071 28407
rect 22569 28373 22603 28407
rect 24869 28373 24903 28407
rect 29837 28373 29871 28407
rect 5089 28169 5123 28203
rect 29653 28169 29687 28203
rect 30021 28169 30055 28203
rect 34161 28169 34195 28203
rect 1409 28101 1443 28135
rect 15853 28101 15887 28135
rect 23673 28101 23707 28135
rect 32505 28101 32539 28135
rect 2789 28033 2823 28067
rect 5273 28033 5307 28067
rect 9137 28033 9171 28067
rect 14933 28033 14967 28067
rect 15577 28033 15611 28067
rect 16865 28033 16899 28067
rect 25513 28033 25547 28067
rect 27261 28033 27295 28067
rect 32689 28033 32723 28067
rect 33977 28033 34011 28067
rect 2973 27965 3007 27999
rect 3249 27965 3283 27999
rect 9321 27965 9355 27999
rect 9689 27965 9723 27999
rect 15669 27965 15703 27999
rect 19441 27965 19475 27999
rect 19717 27965 19751 27999
rect 25329 27965 25363 27999
rect 26985 27965 27019 27999
rect 30113 27965 30147 27999
rect 30297 27965 30331 27999
rect 33793 27965 33827 27999
rect 13369 27829 13403 27863
rect 14289 27829 14323 27863
rect 14749 27829 14783 27863
rect 15393 27829 15427 27863
rect 15577 27829 15611 27863
rect 16681 27829 16715 27863
rect 20729 27829 20763 27863
rect 26157 27829 26191 27863
rect 3065 27625 3099 27659
rect 4261 27625 4295 27659
rect 16865 27625 16899 27659
rect 3801 27557 3835 27591
rect 10333 27557 10367 27591
rect 23857 27557 23891 27591
rect 33885 27557 33919 27591
rect 4169 27489 4203 27523
rect 14565 27489 14599 27523
rect 14749 27489 14783 27523
rect 15761 27489 15795 27523
rect 17049 27489 17083 27523
rect 19993 27489 20027 27523
rect 26065 27489 26099 27523
rect 26249 27489 26283 27523
rect 26985 27489 27019 27523
rect 33517 27489 33551 27523
rect 35817 27489 35851 27523
rect 37013 27489 37047 27523
rect 3249 27421 3283 27455
rect 3985 27421 4019 27455
rect 4261 27421 4295 27455
rect 9045 27421 9079 27455
rect 9321 27421 9355 27455
rect 10517 27421 10551 27455
rect 11161 27421 11195 27455
rect 17141 27421 17175 27455
rect 17877 27421 17911 27455
rect 18521 27421 18555 27455
rect 20453 27421 20487 27455
rect 20729 27421 20763 27455
rect 23673 27421 23707 27455
rect 26709 27421 26743 27455
rect 33701 27421 33735 27455
rect 35541 27421 35575 27455
rect 35633 27421 35667 27455
rect 36737 27421 36771 27455
rect 16865 27353 16899 27387
rect 19809 27353 19843 27387
rect 24409 27353 24443 27387
rect 17325 27285 17359 27319
rect 18061 27285 18095 27319
rect 32045 27285 32079 27319
rect 35173 27285 35207 27319
rect 36369 27285 36403 27319
rect 36829 27285 36863 27319
rect 9781 27081 9815 27115
rect 24409 27081 24443 27115
rect 31493 27081 31527 27115
rect 32781 27081 32815 27115
rect 34069 27081 34103 27115
rect 36737 27081 36771 27115
rect 9321 27013 9355 27047
rect 14473 27013 14507 27047
rect 18705 27013 18739 27047
rect 23949 27013 23983 27047
rect 32505 27013 32539 27047
rect 37657 27013 37691 27047
rect 1409 26945 1443 26979
rect 2053 26945 2087 26979
rect 9597 26945 9631 26979
rect 10425 26945 10459 26979
rect 17233 26945 17267 26979
rect 18521 26945 18555 26979
rect 24225 26945 24259 26979
rect 29837 26945 29871 26979
rect 32229 26945 32263 26979
rect 32413 26945 32447 26979
rect 32597 26945 32631 26979
rect 33977 26945 34011 26979
rect 34805 26945 34839 26979
rect 36369 26945 36403 26979
rect 37841 26945 37875 26979
rect 9413 26877 9447 26911
rect 14289 26877 14323 26911
rect 14749 26877 14783 26911
rect 17509 26877 17543 26911
rect 19441 26877 19475 26911
rect 24041 26877 24075 26911
rect 27997 26877 28031 26911
rect 29653 26877 29687 26911
rect 34253 26877 34287 26911
rect 36093 26877 36127 26911
rect 36277 26877 36311 26911
rect 1593 26741 1627 26775
rect 4721 26741 4755 26775
rect 5181 26741 5215 26775
rect 9413 26741 9447 26775
rect 10609 26741 10643 26775
rect 24225 26741 24259 26775
rect 33609 26741 33643 26775
rect 4537 26537 4571 26571
rect 14381 26537 14415 26571
rect 16129 26537 16163 26571
rect 16497 26537 16531 26571
rect 18061 26537 18095 26571
rect 33057 26537 33091 26571
rect 36461 26537 36495 26571
rect 32597 26469 32631 26503
rect 35265 26469 35299 26503
rect 38025 26469 38059 26503
rect 5181 26401 5215 26435
rect 6837 26401 6871 26435
rect 11437 26401 11471 26435
rect 11621 26401 11655 26435
rect 11897 26401 11931 26435
rect 14841 26401 14875 26435
rect 19717 26401 19751 26435
rect 27997 26401 28031 26435
rect 31401 26401 31435 26435
rect 33517 26401 33551 26435
rect 33701 26401 33735 26435
rect 35909 26401 35943 26435
rect 37105 26401 37139 26435
rect 4721 26333 4755 26367
rect 8401 26333 8435 26367
rect 9137 26333 9171 26367
rect 15117 26333 15151 26367
rect 16273 26333 16307 26367
rect 16405 26333 16439 26367
rect 16589 26333 16623 26367
rect 17049 26333 17083 26367
rect 18705 26333 18739 26367
rect 19257 26333 19291 26367
rect 27721 26333 27755 26367
rect 29561 26333 29595 26367
rect 32045 26333 32079 26367
rect 32321 26333 32355 26367
rect 32413 26333 32447 26367
rect 35725 26333 35759 26367
rect 37841 26333 37875 26367
rect 5365 26265 5399 26299
rect 9321 26265 9355 26299
rect 10977 26265 11011 26299
rect 19441 26265 19475 26299
rect 25973 26265 26007 26299
rect 26709 26265 26743 26299
rect 31217 26265 31251 26299
rect 32229 26265 32263 26299
rect 33425 26265 33459 26299
rect 36921 26265 36955 26299
rect 35633 26197 35667 26231
rect 36829 26197 36863 26231
rect 2881 25993 2915 26027
rect 4721 25993 4755 26027
rect 5365 25993 5399 26027
rect 8953 25993 8987 26027
rect 10333 25993 10367 26027
rect 36001 25993 36035 26027
rect 36369 25993 36403 26027
rect 4261 25925 4295 25959
rect 14105 25925 14139 25959
rect 30941 25925 30975 25959
rect 32597 25925 32631 25959
rect 36461 25925 36495 25959
rect 1409 25857 1443 25891
rect 2421 25857 2455 25891
rect 2697 25857 2731 25891
rect 3065 25857 3099 25891
rect 4537 25857 4571 25891
rect 5181 25857 5215 25891
rect 6561 25857 6595 25891
rect 9137 25857 9171 25891
rect 9413 25857 9447 25891
rect 9873 25857 9907 25891
rect 10149 25857 10183 25891
rect 10977 25857 11011 25891
rect 11713 25857 11747 25891
rect 12357 25857 12391 25891
rect 22293 25857 22327 25891
rect 27261 25857 27295 25891
rect 32413 25857 32447 25891
rect 32689 25857 32723 25891
rect 32781 25857 32815 25891
rect 4445 25789 4479 25823
rect 9229 25789 9263 25823
rect 10057 25789 10091 25823
rect 13461 25789 13495 25823
rect 13921 25789 13955 25823
rect 15301 25789 15335 25823
rect 26985 25789 27019 25823
rect 29285 25789 29319 25823
rect 31125 25789 31159 25823
rect 36645 25789 36679 25823
rect 1593 25721 1627 25755
rect 10793 25721 10827 25755
rect 22477 25721 22511 25755
rect 33517 25721 33551 25755
rect 2605 25653 2639 25687
rect 4537 25653 4571 25687
rect 6377 25653 6411 25687
rect 9413 25653 9447 25687
rect 10149 25653 10183 25687
rect 11529 25653 11563 25687
rect 12173 25653 12207 25687
rect 23121 25653 23155 25687
rect 25329 25653 25363 25687
rect 25789 25653 25823 25687
rect 26341 25653 26375 25687
rect 32965 25653 32999 25687
rect 35541 25653 35575 25687
rect 37657 25653 37691 25687
rect 4169 25449 4203 25483
rect 4353 25449 4387 25483
rect 11253 25449 11287 25483
rect 11713 25449 11747 25483
rect 19441 25449 19475 25483
rect 21833 25449 21867 25483
rect 25697 25449 25731 25483
rect 25881 25449 25915 25483
rect 26341 25449 26375 25483
rect 26801 25449 26835 25483
rect 32413 25449 32447 25483
rect 1409 25381 1443 25415
rect 4077 25313 4111 25347
rect 4813 25313 4847 25347
rect 4997 25313 5031 25347
rect 5549 25313 5583 25347
rect 9781 25313 9815 25347
rect 11529 25313 11563 25347
rect 21649 25313 21683 25347
rect 25513 25313 25547 25347
rect 26433 25313 26467 25347
rect 27997 25313 28031 25347
rect 31769 25313 31803 25347
rect 2605 25245 2639 25279
rect 3249 25245 3283 25279
rect 4169 25245 4203 25279
rect 8401 25245 8435 25279
rect 8953 25245 8987 25279
rect 11437 25245 11471 25279
rect 19257 25245 19291 25279
rect 21557 25245 21591 25279
rect 21833 25245 21867 25279
rect 25697 25245 25731 25279
rect 26617 25245 26651 25279
rect 27721 25245 27755 25279
rect 30389 25245 30423 25279
rect 30665 25245 30699 25279
rect 32045 25245 32079 25279
rect 32873 25245 32907 25279
rect 33057 25245 33091 25279
rect 33241 25245 33275 25279
rect 3893 25177 3927 25211
rect 9137 25177 9171 25211
rect 11713 25177 11747 25211
rect 22569 25177 22603 25211
rect 22753 25177 22787 25211
rect 25421 25177 25455 25211
rect 26341 25177 26375 25211
rect 33149 25177 33183 25211
rect 33885 25177 33919 25211
rect 3065 25109 3099 25143
rect 22017 25109 22051 25143
rect 24961 25109 24995 25143
rect 29837 25109 29871 25143
rect 31953 25109 31987 25143
rect 33425 25109 33459 25143
rect 36185 25109 36219 25143
rect 9229 24905 9263 24939
rect 26341 24905 26375 24939
rect 2789 24837 2823 24871
rect 21833 24837 21867 24871
rect 25421 24837 25455 24871
rect 2605 24769 2639 24803
rect 5549 24769 5583 24803
rect 9413 24769 9447 24803
rect 10057 24769 10091 24803
rect 10333 24769 10367 24803
rect 17233 24769 17267 24803
rect 17785 24769 17819 24803
rect 18337 24769 18371 24803
rect 20637 24769 20671 24803
rect 22109 24769 22143 24803
rect 23029 24769 23063 24803
rect 25697 24769 25731 24803
rect 26985 24769 27019 24803
rect 27261 24769 27295 24803
rect 30113 24769 30147 24803
rect 30665 24769 30699 24803
rect 3065 24701 3099 24735
rect 5825 24701 5859 24735
rect 10241 24701 10275 24735
rect 15117 24701 15151 24735
rect 15669 24701 15703 24735
rect 15853 24701 15887 24735
rect 20361 24701 20395 24735
rect 21925 24701 21959 24735
rect 23213 24701 23247 24735
rect 23489 24701 23523 24735
rect 25513 24701 25547 24735
rect 27077 24701 27111 24735
rect 29653 24701 29687 24735
rect 29929 24701 29963 24735
rect 9873 24633 9907 24667
rect 22293 24633 22327 24667
rect 27445 24633 27479 24667
rect 33149 24633 33183 24667
rect 6377 24565 6411 24599
rect 10333 24565 10367 24599
rect 21833 24565 21867 24599
rect 25421 24565 25455 24599
rect 25881 24565 25915 24599
rect 26985 24565 27019 24599
rect 30757 24565 30791 24599
rect 31309 24565 31343 24599
rect 32505 24565 32539 24599
rect 1593 24361 1627 24395
rect 3893 24361 3927 24395
rect 4353 24361 4387 24395
rect 14289 24361 14323 24395
rect 17141 24361 17175 24395
rect 18153 24361 18187 24395
rect 18337 24361 18371 24395
rect 22937 24361 22971 24395
rect 23857 24361 23891 24395
rect 25605 24361 25639 24395
rect 26065 24361 26099 24395
rect 16681 24293 16715 24327
rect 24593 24293 24627 24327
rect 4261 24225 4295 24259
rect 15945 24225 15979 24259
rect 16221 24225 16255 24259
rect 16957 24225 16991 24259
rect 17969 24225 18003 24259
rect 21741 24225 21775 24259
rect 27537 24225 27571 24259
rect 32321 24225 32355 24259
rect 33333 24225 33367 24259
rect 1409 24157 1443 24191
rect 2053 24157 2087 24191
rect 4077 24157 4111 24191
rect 4997 24157 5031 24191
rect 5641 24157 5675 24191
rect 6101 24157 6135 24191
rect 16865 24157 16899 24191
rect 18153 24157 18187 24191
rect 19441 24157 19475 24191
rect 20177 24157 20211 24191
rect 20453 24157 20487 24191
rect 21465 24157 21499 24191
rect 22753 24157 22787 24191
rect 23673 24157 23707 24191
rect 24409 24157 24443 24191
rect 25053 24157 25087 24191
rect 25789 24157 25823 24191
rect 25881 24157 25915 24191
rect 26617 24157 26651 24191
rect 27261 24157 27295 24191
rect 32597 24157 32631 24191
rect 33517 24157 33551 24191
rect 4353 24089 4387 24123
rect 17141 24089 17175 24123
rect 17877 24089 17911 24123
rect 25605 24089 25639 24123
rect 4813 24021 4847 24055
rect 5457 24021 5491 24055
rect 19257 24021 19291 24055
rect 26801 24021 26835 24055
rect 33701 24021 33735 24055
rect 17601 23817 17635 23851
rect 24041 23817 24075 23851
rect 27629 23817 27663 23851
rect 18061 23749 18095 23783
rect 29837 23749 29871 23783
rect 4813 23681 4847 23715
rect 7205 23681 7239 23715
rect 16872 23681 16906 23715
rect 17141 23681 17175 23715
rect 17785 23681 17819 23715
rect 19081 23681 19115 23715
rect 20361 23681 20395 23715
rect 22109 23681 22143 23715
rect 23121 23681 23155 23715
rect 23397 23681 23431 23715
rect 25881 23681 25915 23715
rect 30021 23681 30055 23715
rect 34345 23681 34379 23715
rect 16957 23613 16991 23647
rect 17877 23613 17911 23647
rect 20085 23613 20119 23647
rect 21833 23613 21867 23647
rect 23213 23613 23247 23647
rect 24593 23613 24627 23647
rect 24869 23613 24903 23647
rect 28181 23613 28215 23647
rect 7389 23545 7423 23579
rect 18889 23545 18923 23579
rect 23581 23545 23615 23579
rect 4629 23477 4663 23511
rect 12357 23477 12391 23511
rect 15301 23477 15335 23511
rect 16681 23477 16715 23511
rect 17141 23477 17175 23511
rect 18061 23477 18095 23511
rect 23121 23477 23155 23511
rect 27077 23477 27111 23511
rect 30481 23477 30515 23511
rect 32689 23477 32723 23511
rect 34529 23477 34563 23511
rect 34989 23477 35023 23511
rect 4445 23273 4479 23307
rect 6653 23273 6687 23307
rect 12541 23273 12575 23307
rect 13277 23273 13311 23307
rect 17785 23273 17819 23307
rect 18521 23273 18555 23307
rect 20361 23273 20395 23307
rect 36185 23273 36219 23307
rect 3985 23205 4019 23239
rect 4353 23137 4387 23171
rect 10609 23137 10643 23171
rect 16865 23137 16899 23171
rect 17693 23137 17727 23171
rect 18337 23137 18371 23171
rect 20269 23137 20303 23171
rect 27445 23137 27479 23171
rect 27629 23137 27663 23171
rect 30665 23137 30699 23171
rect 1409 23069 1443 23103
rect 2605 23069 2639 23103
rect 3249 23069 3283 23103
rect 4169 23069 4203 23103
rect 7665 23069 7699 23103
rect 10885 23069 10919 23103
rect 11345 23069 11379 23103
rect 12725 23069 12759 23103
rect 13461 23069 13495 23103
rect 17509 23069 17543 23103
rect 17785 23069 17819 23103
rect 18245 23069 18279 23103
rect 18521 23069 18555 23103
rect 20361 23069 20395 23103
rect 29929 23069 29963 23103
rect 30849 23069 30883 23103
rect 31033 23069 31067 23103
rect 31677 23069 31711 23103
rect 33977 23069 34011 23103
rect 34805 23069 34839 23103
rect 4445 23001 4479 23035
rect 7849 23001 7883 23035
rect 15025 23001 15059 23035
rect 16681 23001 16715 23035
rect 20085 23001 20119 23035
rect 25789 23001 25823 23035
rect 35050 23001 35084 23035
rect 1593 22933 1627 22967
rect 3065 22933 3099 22967
rect 17325 22933 17359 22967
rect 18705 22933 18739 22967
rect 20545 22933 20579 22967
rect 22937 22933 22971 22967
rect 25237 22933 25271 22967
rect 30113 22933 30147 22967
rect 31493 22933 31527 22967
rect 34161 22933 34195 22967
rect 6377 22729 6411 22763
rect 29929 22729 29963 22763
rect 30665 22729 30699 22763
rect 31125 22729 31159 22763
rect 33885 22729 33919 22763
rect 1409 22661 1443 22695
rect 2973 22661 3007 22695
rect 7665 22661 7699 22695
rect 18153 22661 18187 22695
rect 19073 22661 19107 22695
rect 35142 22661 35176 22695
rect 2789 22593 2823 22627
rect 5273 22593 5307 22627
rect 6561 22593 6595 22627
rect 10149 22593 10183 22627
rect 11529 22593 11563 22627
rect 16037 22593 16071 22627
rect 16865 22593 16899 22627
rect 17877 22593 17911 22627
rect 18797 22593 18831 22627
rect 19533 22593 19567 22627
rect 20821 22593 20855 22627
rect 22845 22593 22879 22627
rect 23121 22593 23155 22627
rect 24777 22593 24811 22627
rect 27445 22593 27479 22627
rect 29561 22593 29595 22627
rect 29745 22593 29779 22627
rect 30757 22593 30791 22627
rect 33701 22593 33735 22627
rect 3249 22525 3283 22559
rect 9873 22525 9907 22559
rect 18061 22525 18095 22559
rect 18981 22525 19015 22559
rect 23029 22525 23063 22559
rect 30481 22525 30515 22559
rect 33057 22525 33091 22559
rect 33517 22525 33551 22559
rect 34897 22525 34931 22559
rect 12173 22457 12207 22491
rect 16681 22457 16715 22491
rect 22385 22457 22419 22491
rect 23305 22457 23339 22491
rect 27629 22457 27663 22491
rect 5089 22389 5123 22423
rect 5825 22389 5859 22423
rect 7113 22389 7147 22423
rect 11713 22389 11747 22423
rect 13093 22389 13127 22423
rect 15025 22389 15059 22423
rect 15853 22389 15887 22423
rect 17693 22389 17727 22423
rect 18153 22389 18187 22423
rect 18613 22389 18647 22423
rect 18797 22389 18831 22423
rect 19717 22389 19751 22423
rect 20637 22389 20671 22423
rect 23121 22389 23155 22423
rect 24961 22389 24995 22423
rect 29009 22389 29043 22423
rect 34437 22389 34471 22423
rect 36277 22389 36311 22423
rect 4261 22185 4295 22219
rect 4445 22185 4479 22219
rect 10149 22185 10183 22219
rect 29561 22185 29595 22219
rect 4169 22049 4203 22083
rect 5917 22049 5951 22083
rect 9045 22049 9079 22083
rect 10333 22049 10367 22083
rect 11161 22049 11195 22083
rect 12633 22049 12667 22083
rect 14933 22049 14967 22083
rect 15117 22049 15151 22083
rect 15393 22049 15427 22083
rect 20361 22049 20395 22083
rect 20729 22049 20763 22083
rect 27629 22049 27663 22083
rect 30205 22049 30239 22083
rect 33057 22049 33091 22083
rect 2697 21981 2731 22015
rect 4261 21981 4295 22015
rect 4997 21981 5031 22015
rect 5641 21981 5675 22015
rect 6929 21981 6963 22015
rect 7665 21981 7699 22015
rect 9505 21981 9539 22015
rect 10425 21981 10459 22015
rect 19717 21981 19751 22015
rect 20177 21981 20211 22015
rect 23581 21981 23615 22015
rect 27813 21981 27847 22015
rect 31125 21981 31159 22015
rect 33793 21981 33827 22015
rect 34161 21981 34195 22015
rect 35265 21981 35299 22015
rect 36093 21981 36127 22015
rect 3985 21913 4019 21947
rect 10149 21913 10183 21947
rect 11345 21913 11379 21947
rect 17601 21913 17635 21947
rect 18153 21913 18187 21947
rect 25973 21913 26007 21947
rect 31392 21913 31426 21947
rect 33977 21913 34011 21947
rect 36338 21913 36372 21947
rect 5181 21845 5215 21879
rect 7113 21845 7147 21879
rect 7849 21845 7883 21879
rect 9689 21845 9723 21879
rect 10609 21845 10643 21879
rect 13553 21845 13587 21879
rect 18245 21845 18279 21879
rect 22477 21845 22511 21879
rect 29009 21845 29043 21879
rect 29929 21845 29963 21879
rect 30021 21845 30055 21879
rect 32505 21845 32539 21879
rect 35449 21845 35483 21879
rect 37473 21845 37507 21879
rect 6837 21641 6871 21675
rect 10701 21641 10735 21675
rect 32137 21641 32171 21675
rect 35909 21641 35943 21675
rect 38025 21641 38059 21675
rect 2881 21573 2915 21607
rect 11713 21573 11747 21607
rect 19625 21573 19659 21607
rect 30012 21573 30046 21607
rect 1409 21505 1443 21539
rect 2053 21505 2087 21539
rect 2697 21505 2731 21539
rect 4537 21505 4571 21539
rect 5457 21505 5491 21539
rect 6377 21505 6411 21539
rect 6561 21505 6595 21539
rect 6653 21505 6687 21539
rect 7297 21505 7331 21539
rect 9689 21505 9723 21539
rect 10885 21505 10919 21539
rect 11529 21505 11563 21539
rect 13829 21505 13863 21539
rect 14565 21505 14599 21539
rect 17141 21505 17175 21539
rect 25237 21505 25271 21539
rect 25973 21505 26007 21539
rect 37841 21505 37875 21539
rect 8953 21437 8987 21471
rect 9413 21437 9447 21471
rect 12541 21437 12575 21471
rect 17417 21437 17451 21471
rect 19441 21437 19475 21471
rect 19901 21437 19935 21471
rect 23673 21437 23707 21471
rect 25053 21437 25087 21471
rect 29745 21437 29779 21471
rect 1593 21301 1627 21335
rect 5273 21301 5307 21335
rect 6377 21301 6411 21335
rect 7481 21301 7515 21335
rect 7941 21301 7975 21335
rect 14013 21301 14047 21335
rect 26249 21301 26283 21335
rect 31125 21301 31159 21335
rect 4629 21097 4663 21131
rect 8309 21097 8343 21131
rect 11253 21097 11287 21131
rect 11897 21097 11931 21131
rect 12357 21097 12391 21131
rect 19717 21097 19751 21131
rect 24409 21097 24443 21131
rect 25329 21097 25363 21131
rect 29929 21097 29963 21131
rect 30481 21097 30515 21131
rect 4537 20961 4571 20995
rect 5273 20961 5307 20995
rect 5549 20961 5583 20995
rect 9321 20961 9355 20995
rect 9597 20961 9631 20995
rect 11069 20961 11103 20995
rect 11989 20961 12023 20995
rect 18153 20961 18187 20995
rect 24501 20961 24535 20995
rect 28457 20961 28491 20995
rect 31033 20961 31067 20995
rect 4353 20893 4387 20927
rect 4629 20893 4663 20927
rect 5089 20893 5123 20927
rect 11253 20893 11287 20927
rect 12173 20893 12207 20927
rect 12909 20893 12943 20927
rect 16313 20893 16347 20927
rect 17877 20893 17911 20927
rect 22661 20893 22695 20927
rect 22937 20893 22971 20927
rect 24409 20893 24443 20927
rect 24685 20893 24719 20927
rect 25513 20893 25547 20927
rect 28917 20893 28951 20927
rect 10977 20825 11011 20859
rect 11897 20825 11931 20859
rect 28733 20825 28767 20859
rect 30941 20825 30975 20859
rect 4169 20757 4203 20791
rect 11437 20757 11471 20791
rect 13093 20757 13127 20791
rect 24869 20757 24903 20791
rect 25973 20757 26007 20791
rect 30849 20757 30883 20791
rect 5457 20553 5491 20587
rect 11621 20553 11655 20587
rect 12725 20553 12759 20587
rect 14013 20553 14047 20587
rect 24685 20553 24719 20587
rect 26065 20553 26099 20587
rect 7665 20485 7699 20519
rect 16865 20485 16899 20519
rect 24225 20485 24259 20519
rect 1409 20417 1443 20451
rect 2053 20417 2087 20451
rect 3341 20417 3375 20451
rect 4997 20417 5031 20451
rect 5181 20417 5215 20451
rect 5273 20417 5307 20451
rect 11805 20417 11839 20451
rect 12909 20417 12943 20451
rect 16681 20417 16715 20451
rect 24501 20417 24535 20451
rect 25881 20417 25915 20451
rect 7481 20349 7515 20383
rect 8033 20349 8067 20383
rect 17141 20349 17175 20383
rect 24317 20349 24351 20383
rect 20085 20281 20119 20315
rect 1593 20213 1627 20247
rect 3157 20213 3191 20247
rect 5273 20213 5307 20247
rect 13369 20213 13403 20247
rect 19533 20213 19567 20247
rect 23673 20213 23707 20247
rect 24409 20213 24443 20247
rect 5181 20009 5215 20043
rect 8033 20009 8067 20043
rect 22937 20009 22971 20043
rect 24409 20009 24443 20043
rect 36001 20009 36035 20043
rect 37105 20009 37139 20043
rect 12081 19941 12115 19975
rect 7573 19873 7607 19907
rect 12541 19873 12575 19907
rect 14933 19873 14967 19907
rect 16957 19873 16991 19907
rect 17969 19873 18003 19907
rect 24501 19873 24535 19907
rect 25329 19873 25363 19907
rect 36461 19873 36495 19907
rect 37565 19873 37599 19907
rect 37657 19873 37691 19907
rect 2421 19805 2455 19839
rect 7297 19805 7331 19839
rect 12817 19805 12851 19839
rect 14473 19805 14507 19839
rect 16773 19805 16807 19839
rect 19625 19805 19659 19839
rect 22293 19805 22327 19839
rect 22753 19805 22787 19839
rect 23397 19805 23431 19839
rect 24409 19805 24443 19839
rect 24685 19805 24719 19839
rect 26065 19805 26099 19839
rect 26341 19805 26375 19839
rect 14657 19737 14691 19771
rect 36553 19737 36587 19771
rect 20913 19669 20947 19703
rect 23581 19669 23615 19703
rect 24869 19669 24903 19703
rect 36461 19669 36495 19703
rect 37473 19669 37507 19703
rect 5365 19465 5399 19499
rect 8401 19465 8435 19499
rect 19809 19465 19843 19499
rect 22017 19465 22051 19499
rect 24593 19465 24627 19499
rect 2605 19397 2639 19431
rect 18797 19397 18831 19431
rect 20729 19397 20763 19431
rect 23305 19397 23339 19431
rect 27261 19397 27295 19431
rect 28917 19397 28951 19431
rect 2421 19329 2455 19363
rect 5549 19329 5583 19363
rect 6837 19329 6871 19363
rect 8217 19329 8251 19363
rect 12173 19329 12207 19363
rect 12817 19329 12851 19363
rect 14473 19329 14507 19363
rect 16865 19329 16899 19363
rect 19901 19329 19935 19363
rect 21833 19329 21867 19363
rect 22477 19329 22511 19363
rect 24133 19329 24167 19363
rect 24317 19329 24351 19363
rect 24409 19329 24443 19363
rect 32321 19329 32355 19363
rect 32505 19329 32539 19363
rect 35613 19329 35647 19363
rect 2881 19261 2915 19295
rect 7481 19261 7515 19295
rect 29101 19261 29135 19295
rect 33057 19261 33091 19295
rect 34805 19261 34839 19295
rect 35357 19261 35391 19295
rect 18981 19193 19015 19227
rect 7021 19125 7055 19159
rect 12357 19125 12391 19159
rect 13001 19125 13035 19159
rect 13461 19125 13495 19159
rect 18153 19125 18187 19159
rect 20821 19125 20855 19159
rect 22661 19125 22695 19159
rect 24409 19125 24443 19159
rect 32413 19125 32447 19159
rect 36737 19125 36771 19159
rect 6009 18921 6043 18955
rect 7665 18921 7699 18955
rect 12633 18921 12667 18955
rect 14289 18921 14323 18955
rect 18521 18921 18555 18955
rect 23581 18921 23615 18955
rect 24409 18921 24443 18955
rect 29653 18921 29687 18955
rect 34989 18921 35023 18955
rect 36829 18921 36863 18955
rect 8125 18853 8159 18887
rect 33977 18853 34011 18887
rect 5825 18785 5859 18819
rect 6653 18785 6687 18819
rect 7205 18785 7239 18819
rect 7757 18785 7791 18819
rect 23121 18785 23155 18819
rect 24501 18785 24535 18819
rect 28549 18785 28583 18819
rect 35449 18785 35483 18819
rect 37841 18785 37875 18819
rect 1409 18717 1443 18751
rect 2053 18717 2087 18751
rect 5089 18717 5123 18751
rect 5733 18717 5767 18751
rect 7941 18717 7975 18751
rect 9597 18717 9631 18751
rect 11989 18717 12023 18751
rect 12817 18717 12851 18751
rect 12909 18717 12943 18751
rect 14105 18717 14139 18751
rect 17601 18717 17635 18751
rect 18337 18717 18371 18751
rect 19349 18717 19383 18751
rect 19717 18717 19751 18751
rect 19993 18717 20027 18751
rect 20729 18717 20763 18751
rect 21649 18717 21683 18751
rect 22845 18717 22879 18751
rect 24409 18717 24443 18751
rect 24685 18717 24719 18751
rect 25789 18717 25823 18751
rect 26433 18717 26467 18751
rect 29009 18717 29043 18751
rect 30757 18717 30791 18751
rect 32597 18717 32631 18751
rect 32689 18717 32723 18751
rect 32873 18717 32907 18751
rect 32965 18717 32999 18751
rect 33793 18717 33827 18751
rect 34805 18717 34839 18751
rect 34989 18717 35023 18751
rect 37414 18717 37448 18751
rect 37933 18717 37967 18751
rect 6009 18649 6043 18683
rect 7665 18649 7699 18683
rect 8953 18649 8987 18683
rect 12633 18649 12667 18683
rect 28825 18649 28859 18683
rect 31002 18649 31036 18683
rect 35694 18649 35728 18683
rect 1593 18581 1627 18615
rect 5549 18581 5583 18615
rect 12173 18581 12207 18615
rect 13093 18581 13127 18615
rect 20637 18581 20671 18615
rect 21833 18581 21867 18615
rect 24869 18581 24903 18615
rect 25973 18581 26007 18615
rect 26617 18581 26651 18615
rect 32137 18581 32171 18615
rect 33149 18581 33183 18615
rect 37289 18581 37323 18615
rect 37473 18581 37507 18615
rect 25421 18377 25455 18411
rect 29837 18377 29871 18411
rect 29929 18377 29963 18411
rect 30297 18377 30331 18411
rect 32781 18377 32815 18411
rect 35357 18377 35391 18411
rect 35909 18377 35943 18411
rect 36093 18377 36127 18411
rect 37473 18377 37507 18411
rect 13185 18309 13219 18343
rect 17785 18309 17819 18343
rect 24685 18309 24719 18343
rect 27169 18309 27203 18343
rect 28825 18309 28859 18343
rect 30757 18309 30791 18343
rect 32413 18309 32447 18343
rect 32597 18309 32631 18343
rect 3157 18241 3191 18275
rect 4169 18241 4203 18275
rect 4721 18241 4755 18275
rect 5549 18241 5583 18275
rect 5825 18241 5859 18275
rect 6377 18241 6411 18275
rect 6653 18241 6687 18275
rect 7297 18241 7331 18275
rect 7573 18241 7607 18275
rect 9137 18241 9171 18275
rect 12081 18241 12115 18275
rect 12357 18241 12391 18275
rect 17601 18241 17635 18275
rect 21281 18241 21315 18275
rect 22385 18241 22419 18275
rect 24869 18241 24903 18275
rect 30941 18241 30975 18275
rect 35265 18241 35299 18275
rect 35449 18241 35483 18275
rect 36034 18241 36068 18275
rect 36461 18241 36495 18275
rect 36553 18241 36587 18275
rect 37473 18241 37507 18275
rect 5641 18173 5675 18207
rect 6561 18173 6595 18207
rect 7389 18173 7423 18207
rect 8217 18173 8251 18207
rect 9321 18173 9355 18207
rect 9689 18173 9723 18207
rect 12265 18173 12299 18207
rect 13001 18173 13035 18207
rect 14841 18173 14875 18207
rect 18245 18173 18279 18207
rect 24409 18173 24443 18207
rect 26985 18173 27019 18207
rect 29745 18173 29779 18207
rect 4905 18105 4939 18139
rect 3249 18037 3283 18071
rect 5365 18037 5399 18071
rect 5825 18037 5859 18071
rect 6469 18037 6503 18071
rect 6837 18037 6871 18071
rect 7297 18037 7331 18071
rect 7757 18037 7791 18071
rect 12357 18037 12391 18071
rect 12541 18037 12575 18071
rect 20085 18037 20119 18071
rect 22293 18037 22327 18071
rect 31125 18037 31159 18071
rect 2513 17833 2547 17867
rect 3939 17833 3973 17867
rect 7757 17833 7791 17867
rect 8401 17833 8435 17867
rect 9413 17833 9447 17867
rect 10241 17833 10275 17867
rect 12357 17833 12391 17867
rect 16129 17833 16163 17867
rect 18245 17833 18279 17867
rect 29653 17833 29687 17867
rect 30757 17833 30791 17867
rect 32597 17833 32631 17867
rect 38025 17833 38059 17867
rect 4077 17765 4111 17799
rect 9781 17765 9815 17799
rect 2605 17697 2639 17731
rect 4169 17697 4203 17731
rect 5089 17697 5123 17731
rect 5549 17697 5583 17731
rect 9413 17697 9447 17731
rect 12449 17697 12483 17731
rect 20085 17697 20119 17731
rect 21925 17697 21959 17731
rect 1409 17629 1443 17663
rect 2513 17629 2547 17663
rect 9597 17629 9631 17663
rect 10425 17629 10459 17663
rect 12265 17629 12299 17663
rect 12541 17629 12575 17663
rect 13185 17629 13219 17663
rect 14105 17629 14139 17663
rect 16313 17629 16347 17663
rect 30573 17629 30607 17663
rect 31217 17629 31251 17663
rect 33149 17629 33183 17663
rect 35265 17629 35299 17663
rect 37381 17629 37415 17663
rect 37841 17629 37875 17663
rect 3801 17561 3835 17595
rect 5273 17561 5307 17595
rect 9321 17561 9355 17595
rect 18153 17561 18187 17595
rect 19257 17561 19291 17595
rect 20269 17561 20303 17595
rect 31484 17561 31518 17595
rect 1593 17493 1627 17527
rect 2881 17493 2915 17527
rect 4445 17493 4479 17527
rect 12725 17493 12759 17527
rect 13369 17493 13403 17527
rect 17601 17493 17635 17527
rect 3433 17289 3467 17323
rect 5457 17289 5491 17323
rect 18797 17289 18831 17323
rect 20821 17289 20855 17323
rect 29561 17289 29595 17323
rect 30389 17289 30423 17323
rect 31401 17289 31435 17323
rect 35633 17289 35667 17323
rect 1409 17221 1443 17255
rect 2973 17221 3007 17255
rect 3985 17221 4019 17255
rect 13553 17221 13587 17255
rect 18153 17221 18187 17255
rect 22477 17221 22511 17255
rect 23397 17221 23431 17255
rect 30481 17221 30515 17255
rect 2145 17153 2179 17187
rect 3249 17153 3283 17187
rect 4261 17153 4295 17187
rect 5641 17153 5675 17187
rect 12449 17153 12483 17187
rect 12725 17153 12759 17187
rect 13369 17153 13403 17187
rect 22753 17153 22787 17187
rect 23673 17153 23707 17187
rect 27261 17153 27295 17187
rect 31217 17153 31251 17187
rect 2237 17085 2271 17119
rect 3065 17085 3099 17119
rect 4077 17085 4111 17119
rect 12633 17085 12667 17119
rect 15117 17085 15151 17119
rect 18521 17085 18555 17119
rect 22661 17085 22695 17119
rect 23489 17085 23523 17119
rect 30573 17085 30607 17119
rect 2145 16949 2179 16983
rect 2513 16949 2547 16983
rect 3249 16949 3283 16983
rect 4077 16949 4111 16983
rect 4445 16949 4479 16983
rect 9137 16949 9171 16983
rect 12725 16949 12759 16983
rect 12909 16949 12943 16983
rect 18318 16949 18352 16983
rect 18429 16949 18463 16983
rect 22477 16949 22511 16983
rect 22937 16949 22971 16983
rect 23397 16949 23431 16983
rect 23857 16949 23891 16983
rect 27077 16949 27111 16983
rect 30021 16949 30055 16983
rect 2973 16745 3007 16779
rect 3966 16745 4000 16779
rect 4077 16745 4111 16779
rect 12725 16745 12759 16779
rect 18337 16745 18371 16779
rect 23397 16745 23431 16779
rect 28549 16745 28583 16779
rect 35265 16745 35299 16779
rect 17233 16677 17267 16711
rect 30481 16677 30515 16711
rect 4169 16609 4203 16643
rect 9137 16609 9171 16643
rect 9689 16609 9723 16643
rect 12725 16609 12759 16643
rect 18337 16609 18371 16643
rect 19901 16609 19935 16643
rect 20177 16609 20211 16643
rect 23305 16609 23339 16643
rect 26617 16609 26651 16643
rect 35817 16609 35851 16643
rect 2605 16541 2639 16575
rect 3801 16541 3835 16575
rect 7757 16541 7791 16575
rect 12909 16541 12943 16575
rect 18153 16541 18187 16575
rect 18429 16541 18463 16575
rect 23121 16541 23155 16575
rect 23397 16541 23431 16575
rect 26884 16541 26918 16575
rect 30113 16541 30147 16575
rect 30297 16541 30331 16575
rect 2789 16473 2823 16507
rect 4537 16473 4571 16507
rect 9321 16473 9355 16507
rect 12633 16473 12667 16507
rect 17049 16473 17083 16507
rect 36084 16473 36118 16507
rect 7573 16405 7607 16439
rect 13093 16405 13127 16439
rect 16405 16405 16439 16439
rect 18613 16405 18647 16439
rect 23581 16405 23615 16439
rect 27997 16405 28031 16439
rect 29561 16405 29595 16439
rect 37197 16405 37231 16439
rect 9413 16201 9447 16235
rect 27169 16201 27203 16235
rect 28457 16201 28491 16235
rect 36277 16201 36311 16235
rect 28365 16133 28399 16167
rect 35173 16133 35207 16167
rect 1409 16065 1443 16099
rect 2053 16065 2087 16099
rect 3157 16065 3191 16099
rect 6561 16065 6595 16099
rect 9597 16065 9631 16099
rect 12909 16065 12943 16099
rect 16681 16065 16715 16099
rect 16957 16065 16991 16099
rect 17785 16065 17819 16099
rect 24869 16065 24903 16099
rect 27353 16065 27387 16099
rect 34897 16065 34931 16099
rect 35633 16065 35667 16099
rect 35817 16065 35851 16099
rect 35909 16065 35943 16099
rect 36001 16065 36035 16099
rect 16865 15997 16899 16031
rect 22569 15997 22603 16031
rect 22753 15997 22787 16031
rect 23489 15997 23523 16031
rect 27537 15997 27571 16031
rect 28641 15997 28675 16031
rect 35173 15997 35207 16031
rect 3249 15929 3283 15963
rect 17969 15929 18003 15963
rect 27997 15929 28031 15963
rect 1593 15861 1627 15895
rect 6377 15861 6411 15895
rect 12725 15861 12759 15895
rect 13369 15861 13403 15895
rect 16865 15861 16899 15895
rect 17141 15861 17175 15895
rect 20821 15861 20855 15895
rect 25053 15861 25087 15895
rect 34989 15861 35023 15895
rect 17325 15657 17359 15691
rect 23213 15657 23247 15691
rect 32689 15657 32723 15691
rect 35817 15657 35851 15691
rect 36093 15657 36127 15691
rect 16221 15589 16255 15623
rect 5733 15521 5767 15555
rect 16313 15521 16347 15555
rect 18705 15521 18739 15555
rect 19257 15521 19291 15555
rect 20821 15521 20855 15555
rect 22201 15521 22235 15555
rect 25145 15521 25179 15555
rect 35817 15521 35851 15555
rect 5457 15453 5491 15487
rect 6193 15453 6227 15487
rect 7481 15453 7515 15487
rect 8953 15453 8987 15487
rect 12633 15453 12667 15487
rect 13277 15453 13311 15487
rect 13461 15453 13495 15487
rect 15945 15453 15979 15487
rect 16092 15453 16126 15487
rect 17141 15453 17175 15487
rect 19533 15453 19567 15487
rect 23397 15453 23431 15487
rect 25421 15453 25455 15487
rect 30021 15453 30055 15487
rect 32505 15453 32539 15487
rect 35725 15453 35759 15487
rect 16681 15385 16715 15419
rect 21005 15385 21039 15419
rect 30205 15385 30239 15419
rect 12173 15317 12207 15351
rect 13461 15317 13495 15351
rect 15393 15317 15427 15351
rect 17877 15317 17911 15351
rect 27813 15317 27847 15351
rect 28457 15317 28491 15351
rect 9689 15113 9723 15147
rect 19717 15113 19751 15147
rect 20545 15113 20579 15147
rect 29745 15113 29779 15147
rect 4169 15045 4203 15079
rect 7573 15045 7607 15079
rect 10149 15045 10183 15079
rect 12725 15045 12759 15079
rect 18613 15045 18647 15079
rect 24409 15045 24443 15079
rect 26065 15045 26099 15079
rect 27169 15045 27203 15079
rect 28825 15045 28859 15079
rect 35449 15045 35483 15079
rect 1409 14977 1443 15011
rect 2053 14977 2087 15011
rect 7389 14977 7423 15011
rect 9873 14977 9907 15011
rect 12541 14977 12575 15011
rect 19257 14977 19291 15011
rect 19533 14977 19567 15011
rect 20361 14977 20395 15011
rect 22661 14977 22695 15011
rect 35265 14977 35299 15011
rect 35541 14977 35575 15011
rect 3985 14909 4019 14943
rect 4445 14909 4479 14943
rect 7849 14909 7883 14943
rect 10057 14909 10091 14943
rect 13001 14909 13035 14943
rect 16129 14909 16163 14943
rect 16773 14909 16807 14943
rect 16957 14909 16991 14943
rect 19441 14909 19475 14943
rect 26249 14909 26283 14943
rect 26985 14909 27019 14943
rect 35265 14841 35299 14875
rect 1593 14773 1627 14807
rect 9873 14773 9907 14807
rect 19349 14773 19383 14807
rect 3249 14569 3283 14603
rect 9413 14569 9447 14603
rect 10333 14569 10367 14603
rect 19349 14569 19383 14603
rect 19809 14569 19843 14603
rect 33977 14569 34011 14603
rect 34897 14569 34931 14603
rect 5365 14433 5399 14467
rect 6009 14433 6043 14467
rect 6469 14433 6503 14467
rect 9597 14433 9631 14467
rect 10517 14433 10551 14467
rect 19441 14433 19475 14467
rect 22109 14433 22143 14467
rect 27169 14433 27203 14467
rect 30297 14433 30331 14467
rect 34713 14433 34747 14467
rect 3985 14365 4019 14399
rect 5089 14365 5123 14399
rect 9413 14365 9447 14399
rect 10333 14365 10367 14399
rect 15761 14365 15795 14399
rect 16221 14365 16255 14399
rect 18061 14365 18095 14399
rect 19625 14365 19659 14399
rect 21189 14365 21223 14399
rect 21649 14365 21683 14399
rect 26985 14365 27019 14399
rect 30113 14365 30147 14399
rect 33149 14365 33183 14399
rect 33333 14365 33367 14399
rect 33793 14365 33827 14399
rect 33977 14365 34011 14399
rect 34989 14365 35023 14399
rect 6193 14297 6227 14331
rect 9689 14297 9723 14331
rect 10609 14297 10643 14331
rect 16405 14297 16439 14331
rect 18705 14297 18739 14331
rect 19349 14297 19383 14331
rect 21833 14297 21867 14331
rect 29009 14297 29043 14331
rect 30205 14297 30239 14331
rect 37381 14297 37415 14331
rect 38025 14297 38059 14331
rect 9229 14229 9263 14263
rect 10149 14229 10183 14263
rect 26157 14229 26191 14263
rect 26617 14229 26651 14263
rect 27077 14229 27111 14263
rect 29745 14229 29779 14263
rect 33149 14229 33183 14263
rect 34161 14229 34195 14263
rect 34713 14229 34747 14263
rect 37933 14229 37967 14263
rect 15761 14025 15795 14059
rect 16865 14025 16899 14059
rect 17325 14025 17359 14059
rect 19257 14025 19291 14059
rect 21189 14025 21223 14059
rect 26341 14025 26375 14059
rect 30205 14025 30239 14059
rect 32229 14025 32263 14059
rect 35357 14025 35391 14059
rect 37381 14025 37415 14059
rect 5181 13957 5215 13991
rect 13001 13957 13035 13991
rect 28549 13957 28583 13991
rect 34161 13957 34195 13991
rect 36277 13957 36311 13991
rect 5365 13889 5399 13923
rect 7297 13889 7331 13923
rect 8677 13889 8711 13923
rect 12081 13889 12115 13923
rect 16681 13889 16715 13923
rect 17509 13889 17543 13923
rect 21005 13889 21039 13923
rect 29009 13889 29043 13923
rect 29193 13889 29227 13923
rect 30297 13889 30331 13923
rect 31033 13889 31067 13923
rect 33342 13889 33376 13923
rect 34345 13889 34379 13923
rect 34437 13889 34471 13923
rect 34989 13889 35023 13923
rect 35449 13889 35483 13923
rect 36461 13889 36495 13923
rect 37289 13889 37323 13923
rect 3985 13821 4019 13855
rect 7021 13821 7055 13855
rect 8861 13821 8895 13855
rect 9137 13821 9171 13855
rect 12357 13821 12391 13855
rect 14657 13821 14691 13855
rect 14841 13821 14875 13855
rect 29837 13821 29871 13855
rect 30021 13821 30055 13855
rect 30757 13821 30791 13855
rect 30849 13821 30883 13855
rect 33609 13821 33643 13855
rect 35081 13821 35115 13855
rect 35173 13753 35207 13787
rect 29377 13685 29411 13719
rect 31217 13685 31251 13719
rect 9045 13481 9079 13515
rect 10057 13481 10091 13515
rect 11621 13481 11655 13515
rect 13277 13481 13311 13515
rect 16129 13481 16163 13515
rect 16773 13481 16807 13515
rect 17233 13481 17267 13515
rect 19717 13481 19751 13515
rect 20177 13481 20211 13515
rect 28365 13481 28399 13515
rect 30941 13481 30975 13515
rect 33425 13481 33459 13515
rect 36461 13481 36495 13515
rect 10885 13413 10919 13447
rect 15301 13413 15335 13447
rect 16313 13413 16347 13447
rect 27905 13413 27939 13447
rect 5181 13345 5215 13379
rect 6837 13345 6871 13379
rect 16037 13345 16071 13379
rect 16865 13345 16899 13379
rect 17693 13345 17727 13379
rect 19901 13345 19935 13379
rect 26525 13345 26559 13379
rect 32137 13345 32171 13379
rect 1409 13277 1443 13311
rect 2053 13277 2087 13311
rect 7021 13277 7055 13311
rect 8401 13277 8435 13311
rect 9229 13277 9263 13311
rect 10241 13277 10275 13311
rect 11437 13277 11471 13311
rect 12541 13277 12575 13311
rect 15117 13277 15151 13311
rect 16129 13277 16163 13311
rect 17049 13277 17083 13311
rect 19993 13277 20027 13311
rect 22385 13277 22419 13311
rect 26065 13277 26099 13311
rect 29561 13277 29595 13311
rect 33149 13277 33183 13311
rect 35081 13277 35115 13311
rect 15853 13209 15887 13243
rect 16773 13209 16807 13243
rect 19717 13209 19751 13243
rect 25881 13209 25915 13243
rect 26792 13209 26826 13243
rect 29828 13209 29862 13243
rect 33425 13209 33459 13243
rect 35326 13209 35360 13243
rect 1593 13141 1627 13175
rect 25697 13141 25731 13175
rect 29009 13141 29043 13175
rect 33241 13141 33275 13175
rect 10701 12937 10735 12971
rect 12081 12937 12115 12971
rect 15485 12937 15519 12971
rect 17049 12937 17083 12971
rect 20085 12937 20119 12971
rect 26985 12937 27019 12971
rect 29837 12937 29871 12971
rect 34529 12937 34563 12971
rect 2513 12869 2547 12903
rect 2789 12801 2823 12835
rect 5457 12801 5491 12835
rect 8401 12801 8435 12835
rect 12633 12801 12667 12835
rect 12909 12801 12943 12835
rect 14657 12801 14691 12835
rect 17141 12801 17175 12835
rect 18245 12801 18279 12835
rect 19349 12801 19383 12835
rect 22293 12801 22327 12835
rect 27169 12801 27203 12835
rect 30021 12801 30055 12835
rect 34437 12801 34471 12835
rect 34713 12801 34747 12835
rect 2605 12733 2639 12767
rect 8585 12733 8619 12767
rect 9781 12733 9815 12767
rect 14933 12733 14967 12767
rect 18521 12733 18555 12767
rect 22477 12733 22511 12767
rect 23489 12733 23523 12767
rect 19533 12665 19567 12699
rect 34713 12665 34747 12699
rect 2513 12597 2547 12631
rect 2973 12597 3007 12631
rect 4813 12597 4847 12631
rect 35265 12597 35299 12631
rect 2605 12393 2639 12427
rect 10701 12393 10735 12427
rect 14197 12393 14231 12427
rect 20177 12393 20211 12427
rect 22845 12393 22879 12427
rect 35449 12393 35483 12427
rect 37381 12393 37415 12427
rect 10517 12325 10551 12359
rect 2605 12257 2639 12291
rect 5273 12257 5307 12291
rect 5733 12257 5767 12291
rect 9781 12257 9815 12291
rect 10057 12257 10091 12291
rect 10793 12257 10827 12291
rect 18245 12257 18279 12291
rect 26525 12257 26559 12291
rect 36001 12257 36035 12291
rect 1409 12189 1443 12223
rect 2513 12189 2547 12223
rect 10701 12189 10735 12223
rect 11437 12189 11471 12223
rect 12357 12189 12391 12223
rect 18521 12189 18555 12223
rect 19441 12189 19475 12223
rect 22293 12189 22327 12223
rect 23029 12189 23063 12223
rect 36257 12189 36291 12223
rect 5457 12121 5491 12155
rect 10977 12121 11011 12155
rect 22109 12121 22143 12155
rect 25697 12121 25731 12155
rect 25881 12121 25915 12155
rect 1593 12053 1627 12087
rect 2881 12053 2915 12087
rect 11621 12053 11655 12087
rect 12541 12053 12575 12087
rect 13369 12053 13403 12087
rect 19625 12053 19659 12087
rect 26065 12053 26099 12087
rect 6377 11849 6411 11883
rect 11713 11849 11747 11883
rect 19901 11849 19935 11883
rect 22293 11849 22327 11883
rect 25513 11849 25547 11883
rect 29837 11849 29871 11883
rect 30573 11849 30607 11883
rect 1409 11781 1443 11815
rect 20361 11781 20395 11815
rect 21833 11781 21867 11815
rect 6561 11713 6595 11747
rect 10517 11713 10551 11747
rect 10793 11713 10827 11747
rect 13093 11713 13127 11747
rect 13645 11713 13679 11747
rect 16957 11713 16991 11747
rect 18613 11713 18647 11747
rect 19257 11713 19291 11747
rect 20085 11713 20119 11747
rect 22017 11713 22051 11747
rect 22109 11713 22143 11747
rect 25881 11713 25915 11747
rect 26985 11713 27019 11747
rect 30021 11713 30055 11747
rect 10609 11645 10643 11679
rect 12817 11645 12851 11679
rect 13829 11645 13863 11679
rect 17233 11645 17267 11679
rect 20177 11645 20211 11679
rect 25973 11645 26007 11679
rect 26065 11645 26099 11679
rect 18797 11577 18831 11611
rect 10609 11509 10643 11543
rect 10977 11509 11011 11543
rect 15945 11509 15979 11543
rect 19441 11509 19475 11543
rect 20085 11509 20119 11543
rect 21833 11509 21867 11543
rect 27169 11509 27203 11543
rect 2513 11305 2547 11339
rect 10977 11305 11011 11339
rect 11897 11305 11931 11339
rect 15393 11305 15427 11339
rect 15577 11305 15611 11339
rect 16865 11305 16899 11339
rect 17325 11305 17359 11339
rect 18613 11305 18647 11339
rect 20361 11305 20395 11339
rect 21281 11305 21315 11339
rect 22201 11305 22235 11339
rect 28641 11305 28675 11339
rect 32873 11305 32907 11339
rect 10793 11237 10827 11271
rect 21741 11237 21775 11271
rect 30757 11237 30791 11271
rect 2605 11169 2639 11203
rect 11161 11169 11195 11203
rect 11989 11169 12023 11203
rect 13185 11169 13219 11203
rect 15761 11169 15795 11203
rect 21373 11169 21407 11203
rect 22293 11169 22327 11203
rect 24961 11169 24995 11203
rect 25421 11169 25455 11203
rect 2789 11101 2823 11135
rect 10977 11101 11011 11135
rect 11897 11101 11931 11135
rect 13001 11101 13035 11135
rect 14197 11101 14231 11135
rect 15577 11101 15611 11135
rect 15853 11101 15887 11135
rect 19257 11101 19291 11135
rect 20545 11101 20579 11135
rect 20637 11101 20671 11135
rect 21557 11101 21591 11135
rect 22477 11101 22511 11135
rect 23581 11101 23615 11135
rect 27261 11101 27295 11135
rect 32689 11101 32723 11135
rect 2513 11033 2547 11067
rect 11253 11033 11287 11067
rect 12173 11033 12207 11067
rect 20361 11033 20395 11067
rect 21281 11033 21315 11067
rect 22201 11033 22235 11067
rect 25145 11033 25179 11067
rect 27506 11033 27540 11067
rect 2973 10965 3007 10999
rect 11713 10965 11747 10999
rect 14381 10965 14415 10999
rect 19441 10965 19475 10999
rect 20821 10965 20855 10999
rect 22661 10965 22695 10999
rect 23765 10965 23799 10999
rect 29653 10965 29687 10999
rect 4537 10761 4571 10795
rect 15945 10761 15979 10795
rect 22109 10761 22143 10795
rect 30389 10761 30423 10795
rect 31125 10761 31159 10795
rect 10793 10693 10827 10727
rect 12541 10693 12575 10727
rect 13461 10693 13495 10727
rect 14933 10693 14967 10727
rect 29745 10693 29779 10727
rect 30297 10693 30331 10727
rect 1409 10625 1443 10659
rect 2053 10625 2087 10659
rect 2881 10625 2915 10659
rect 3111 10625 3145 10659
rect 4077 10625 4111 10659
rect 4353 10625 4387 10659
rect 10517 10625 10551 10659
rect 12265 10625 12299 10659
rect 13185 10625 13219 10659
rect 14013 10625 14047 10659
rect 15117 10625 15151 10659
rect 15209 10625 15243 10659
rect 17417 10625 17451 10659
rect 17601 10625 17635 10659
rect 17877 10625 17911 10659
rect 18429 10625 18463 10659
rect 19533 10625 19567 10659
rect 20177 10625 20211 10659
rect 23029 10625 23063 10659
rect 30941 10625 30975 10659
rect 34713 10625 34747 10659
rect 34897 10625 34931 10659
rect 3249 10557 3283 10591
rect 4169 10557 4203 10591
rect 9321 10557 9355 10591
rect 9597 10557 9631 10591
rect 10701 10557 10735 10591
rect 12449 10557 12483 10591
rect 13277 10557 13311 10591
rect 1593 10489 1627 10523
rect 3525 10489 3559 10523
rect 10333 10489 10367 10523
rect 17233 10489 17267 10523
rect 34713 10489 34747 10523
rect 3046 10421 3080 10455
rect 4077 10421 4111 10455
rect 10609 10421 10643 10455
rect 12081 10421 12115 10455
rect 12541 10421 12575 10455
rect 13001 10421 13035 10455
rect 13461 10421 13495 10455
rect 14197 10421 14231 10455
rect 15117 10421 15151 10455
rect 15393 10421 15427 10455
rect 19717 10421 19751 10455
rect 20361 10421 20395 10455
rect 23213 10421 23247 10455
rect 1961 10217 1995 10251
rect 2513 10217 2547 10251
rect 2973 10217 3007 10251
rect 12449 10217 12483 10251
rect 15117 10217 15151 10251
rect 16037 10217 16071 10251
rect 19717 10217 19751 10251
rect 20637 10217 20671 10251
rect 21281 10217 21315 10251
rect 2605 10081 2639 10115
rect 11069 10081 11103 10115
rect 15209 10081 15243 10115
rect 19533 10081 19567 10115
rect 20453 10081 20487 10115
rect 21373 10081 21407 10115
rect 24409 10081 24443 10115
rect 26065 10081 26099 10115
rect 30481 10081 30515 10115
rect 1869 10013 1903 10047
rect 2513 10013 2547 10047
rect 2789 10013 2823 10047
rect 5273 10013 5307 10047
rect 7113 10013 7147 10047
rect 10149 10013 10183 10047
rect 12633 10013 12667 10047
rect 15025 10013 15059 10047
rect 15301 10013 15335 10047
rect 19717 10013 19751 10047
rect 20637 10013 20671 10047
rect 21557 10013 21591 10047
rect 26249 10013 26283 10047
rect 30849 10013 30883 10047
rect 30941 10013 30975 10047
rect 31493 10013 31527 10047
rect 31677 10013 31711 10047
rect 34989 10013 35023 10047
rect 38117 10013 38151 10047
rect 5540 9945 5574 9979
rect 10333 9945 10367 9979
rect 16957 9945 16991 9979
rect 19441 9945 19475 9979
rect 20361 9945 20395 9979
rect 21281 9945 21315 9979
rect 31401 9945 31435 9979
rect 35234 9945 35268 9979
rect 6653 9877 6687 9911
rect 13093 9877 13127 9911
rect 15485 9877 15519 9911
rect 18613 9877 18647 9911
rect 19901 9877 19935 9911
rect 20821 9877 20855 9911
rect 21741 9877 21775 9911
rect 29929 9877 29963 9911
rect 30757 9877 30791 9911
rect 34161 9877 34195 9911
rect 36369 9877 36403 9911
rect 2973 9673 3007 9707
rect 10701 9673 10735 9707
rect 31401 9673 31435 9707
rect 3617 9605 3651 9639
rect 3801 9605 3835 9639
rect 7849 9605 7883 9639
rect 20545 9605 20579 9639
rect 29377 9605 29411 9639
rect 33609 9605 33643 9639
rect 34529 9605 34563 9639
rect 35256 9605 35290 9639
rect 1409 9537 1443 9571
rect 2513 9537 2547 9571
rect 2789 9537 2823 9571
rect 3433 9537 3467 9571
rect 5641 9537 5675 9571
rect 10885 9537 10919 9571
rect 11529 9537 11563 9571
rect 15485 9537 15519 9571
rect 16129 9537 16163 9571
rect 20729 9537 20763 9571
rect 20821 9537 20855 9571
rect 23949 9537 23983 9571
rect 28641 9537 28675 9571
rect 30277 9537 30311 9571
rect 33333 9537 33367 9571
rect 34069 9537 34103 9571
rect 34253 9537 34287 9571
rect 34437 9537 34471 9571
rect 2697 9469 2731 9503
rect 7665 9469 7699 9503
rect 9505 9469 9539 9503
rect 11805 9469 11839 9503
rect 24225 9469 24259 9503
rect 26985 9469 27019 9503
rect 27261 9469 27295 9503
rect 29561 9469 29595 9503
rect 30021 9469 30055 9503
rect 34345 9469 34379 9503
rect 34989 9469 35023 9503
rect 1593 9401 1627 9435
rect 5457 9401 5491 9435
rect 21005 9401 21039 9435
rect 28825 9401 28859 9435
rect 33425 9401 33459 9435
rect 2789 9333 2823 9367
rect 6377 9333 6411 9367
rect 15301 9333 15335 9367
rect 15945 9333 15979 9367
rect 20545 9333 20579 9367
rect 32781 9333 32815 9367
rect 33517 9333 33551 9367
rect 36369 9333 36403 9367
rect 2973 9129 3007 9163
rect 5549 9129 5583 9163
rect 20637 9129 20671 9163
rect 29009 9129 29043 9163
rect 34069 9129 34103 9163
rect 1409 9061 1443 9095
rect 31309 9061 31343 9095
rect 36001 9061 36035 9095
rect 6561 8993 6595 9027
rect 12725 8993 12759 9027
rect 15577 8993 15611 9027
rect 16589 8993 16623 9027
rect 20729 8993 20763 9027
rect 27077 8993 27111 9027
rect 29745 8993 29779 9027
rect 35449 8993 35483 9027
rect 5181 8925 5215 8959
rect 5365 8925 5399 8959
rect 10977 8925 11011 8959
rect 11897 8925 11931 8959
rect 13001 8925 13035 8959
rect 15393 8925 15427 8959
rect 19901 8925 19935 8959
rect 20913 8925 20947 8959
rect 25237 8925 25271 8959
rect 29929 8925 29963 8959
rect 31217 8925 31251 8959
rect 31493 8925 31527 8959
rect 35173 8925 35207 8959
rect 35357 8925 35391 8959
rect 36093 8925 36127 8959
rect 2605 8857 2639 8891
rect 2789 8857 2823 8891
rect 6377 8857 6411 8891
rect 20637 8857 20671 8891
rect 25421 8857 25455 8891
rect 30021 8857 30055 8891
rect 6009 8789 6043 8823
rect 6469 8789 6503 8823
rect 11161 8789 11195 8823
rect 12081 8789 12115 8823
rect 19717 8789 19751 8823
rect 21097 8789 21131 8823
rect 30389 8789 30423 8823
rect 31677 8789 31711 8823
rect 34989 8789 35023 8823
rect 5273 8585 5307 8619
rect 6377 8585 6411 8619
rect 6929 8585 6963 8619
rect 7297 8585 7331 8619
rect 28365 8585 28399 8619
rect 29837 8585 29871 8619
rect 34989 8585 35023 8619
rect 5641 8517 5675 8551
rect 9321 8517 9355 8551
rect 12173 8517 12207 8551
rect 13829 8517 13863 8551
rect 16865 8517 16899 8551
rect 35541 8517 35575 8551
rect 35725 8517 35759 8551
rect 5457 8449 5491 8483
rect 5549 8449 5583 8483
rect 5825 8449 5859 8483
rect 23765 8449 23799 8483
rect 24041 8449 24075 8483
rect 25145 8449 25179 8483
rect 25881 8449 25915 8483
rect 26065 8449 26099 8483
rect 26985 8449 27019 8483
rect 27252 8449 27286 8483
rect 30021 8449 30055 8483
rect 30849 8449 30883 8483
rect 31309 8449 31343 8483
rect 34529 8449 34563 8483
rect 34805 8449 34839 8483
rect 35449 8449 35483 8483
rect 7389 8381 7423 8415
rect 7573 8381 7607 8415
rect 9137 8381 9171 8415
rect 10977 8381 11011 8415
rect 11989 8381 12023 8415
rect 30205 8381 30239 8415
rect 34621 8381 34655 8415
rect 16681 8313 16715 8347
rect 25329 8313 25363 8347
rect 28825 8313 28859 8347
rect 34069 8313 34103 8347
rect 35725 8313 35759 8347
rect 26249 8245 26283 8279
rect 30757 8245 30791 8279
rect 1593 8041 1627 8075
rect 30389 8041 30423 8075
rect 35357 8041 35391 8075
rect 6653 7905 6687 7939
rect 6837 7905 6871 7939
rect 11161 7905 11195 7939
rect 11437 7905 11471 7939
rect 15301 7905 15335 7939
rect 15761 7905 15795 7939
rect 19349 7905 19383 7939
rect 19533 7905 19567 7939
rect 19809 7905 19843 7939
rect 22661 7905 22695 7939
rect 25329 7905 25363 7939
rect 26985 7905 27019 7939
rect 1409 7837 1443 7871
rect 2053 7837 2087 7871
rect 6561 7837 6595 7871
rect 10977 7837 11011 7871
rect 15117 7837 15151 7871
rect 17693 7837 17727 7871
rect 22937 7837 22971 7871
rect 27169 7837 27203 7871
rect 35173 7837 35207 7871
rect 35357 7837 35391 7871
rect 21833 7769 21867 7803
rect 22017 7769 22051 7803
rect 6193 7701 6227 7735
rect 17877 7701 17911 7735
rect 18521 7701 18555 7735
rect 22201 7701 22235 7735
rect 35541 7701 35575 7735
rect 5457 7497 5491 7531
rect 10057 7497 10091 7531
rect 10149 7497 10183 7531
rect 19993 7497 20027 7531
rect 20913 7497 20947 7531
rect 21281 7497 21315 7531
rect 23949 7497 23983 7531
rect 25605 7497 25639 7531
rect 26065 7497 26099 7531
rect 27169 7497 27203 7531
rect 30665 7497 30699 7531
rect 12633 7429 12667 7463
rect 14289 7429 14323 7463
rect 25973 7429 26007 7463
rect 27997 7429 28031 7463
rect 29653 7429 29687 7463
rect 33609 7429 33643 7463
rect 5365 7361 5399 7395
rect 15301 7361 15335 7395
rect 15393 7361 15427 7395
rect 17233 7361 17267 7395
rect 20821 7361 20855 7395
rect 21833 7361 21867 7395
rect 23121 7361 23155 7395
rect 26985 7361 27019 7395
rect 30113 7361 30147 7395
rect 30205 7361 30239 7395
rect 30389 7361 30423 7395
rect 30481 7361 30515 7395
rect 32137 7361 32171 7395
rect 5641 7293 5675 7327
rect 10333 7293 10367 7327
rect 12449 7293 12483 7327
rect 15485 7293 15519 7327
rect 20729 7293 20763 7327
rect 22109 7293 22143 7327
rect 26157 7293 26191 7327
rect 27813 7293 27847 7327
rect 17049 7225 17083 7259
rect 32321 7225 32355 7259
rect 4997 7157 5031 7191
rect 9689 7157 9723 7191
rect 14933 7157 14967 7191
rect 23305 7157 23339 7191
rect 36185 7157 36219 7191
rect 28917 6953 28951 6987
rect 30573 6953 30607 6987
rect 5181 6817 5215 6851
rect 9597 6817 9631 6851
rect 15577 6817 15611 6851
rect 16773 6817 16807 6851
rect 26617 6817 26651 6851
rect 29929 6817 29963 6851
rect 34161 6817 34195 6851
rect 35725 6817 35759 6851
rect 35909 6817 35943 6851
rect 1409 6749 1443 6783
rect 2053 6749 2087 6783
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 7941 6749 7975 6783
rect 8033 6749 8067 6783
rect 8309 6749 8343 6783
rect 9413 6749 9447 6783
rect 15853 6749 15887 6783
rect 17049 6749 17083 6783
rect 18061 6749 18095 6783
rect 18153 6749 18187 6783
rect 18429 6749 18463 6783
rect 19349 6749 19383 6783
rect 22201 6749 22235 6783
rect 26157 6749 26191 6783
rect 28825 6749 28859 6783
rect 29009 6749 29043 6783
rect 29745 6749 29779 6783
rect 30389 6749 30423 6783
rect 31401 6749 31435 6783
rect 33241 6749 33275 6783
rect 33885 6749 33919 6783
rect 34069 6749 34103 6783
rect 35633 6749 35667 6783
rect 36369 6749 36403 6783
rect 8125 6681 8159 6715
rect 18245 6681 18279 6715
rect 20177 6681 20211 6715
rect 21934 6681 21968 6715
rect 29561 6681 29595 6715
rect 32996 6681 33030 6715
rect 36614 6681 36648 6715
rect 1593 6613 1627 6647
rect 3801 6613 3835 6647
rect 4721 6613 4755 6647
rect 5733 6613 5767 6647
rect 7757 6613 7791 6647
rect 8953 6613 8987 6647
rect 9321 6613 9355 6647
rect 15761 6613 15795 6647
rect 16221 6613 16255 6647
rect 16957 6613 16991 6647
rect 17417 6613 17451 6647
rect 17877 6613 17911 6647
rect 20085 6613 20119 6647
rect 20821 6613 20855 6647
rect 25973 6613 26007 6647
rect 31861 6613 31895 6647
rect 33701 6613 33735 6647
rect 35909 6613 35943 6647
rect 37749 6613 37783 6647
rect 3617 6409 3651 6443
rect 8401 6409 8435 6443
rect 14565 6409 14599 6443
rect 14657 6409 14691 6443
rect 15761 6409 15795 6443
rect 21833 6409 21867 6443
rect 33425 6409 33459 6443
rect 36461 6409 36495 6443
rect 4813 6341 4847 6375
rect 25605 6341 25639 6375
rect 33977 6341 34011 6375
rect 2237 6273 2271 6307
rect 2504 6273 2538 6307
rect 4629 6273 4663 6307
rect 4721 6273 4755 6307
rect 4997 6273 5031 6307
rect 17233 6273 17267 6307
rect 22017 6273 22051 6307
rect 23949 6273 23983 6307
rect 32229 6273 32263 6307
rect 33333 6273 33367 6307
rect 33517 6273 33551 6307
rect 35817 6273 35851 6307
rect 36001 6273 36035 6307
rect 36093 6273 36127 6307
rect 36185 6273 36219 6307
rect 37841 6273 37875 6307
rect 14841 6205 14875 6239
rect 25789 6205 25823 6239
rect 35265 6205 35299 6239
rect 5549 6137 5583 6171
rect 17049 6137 17083 6171
rect 4445 6069 4479 6103
rect 14197 6069 14231 6103
rect 20453 6069 20487 6103
rect 20913 6069 20947 6103
rect 32229 6069 32263 6103
rect 38025 6069 38059 6103
rect 2697 5865 2731 5899
rect 4353 5865 4387 5899
rect 9045 5797 9079 5831
rect 6009 5729 6043 5763
rect 8125 5729 8159 5763
rect 16313 5729 16347 5763
rect 19809 5729 19843 5763
rect 22477 5729 22511 5763
rect 26709 5729 26743 5763
rect 30113 5729 30147 5763
rect 30297 5729 30331 5763
rect 31585 5729 31619 5763
rect 2881 5661 2915 5695
rect 4537 5661 4571 5695
rect 4905 5661 4939 5695
rect 5733 5661 5767 5695
rect 7941 5661 7975 5695
rect 10241 5661 10275 5695
rect 14289 5661 14323 5695
rect 14381 5661 14415 5695
rect 14657 5661 14691 5695
rect 19717 5661 19751 5695
rect 20453 5661 20487 5695
rect 22017 5661 22051 5695
rect 26985 5661 27019 5695
rect 31401 5661 31435 5695
rect 4629 5593 4663 5627
rect 4721 5593 4755 5627
rect 14473 5593 14507 5627
rect 22201 5593 22235 5627
rect 3893 5525 3927 5559
rect 5365 5525 5399 5559
rect 5825 5525 5859 5559
rect 6653 5525 6687 5559
rect 7757 5525 7791 5559
rect 10333 5525 10367 5559
rect 14105 5525 14139 5559
rect 15209 5525 15243 5559
rect 19257 5525 19291 5559
rect 19625 5525 19659 5559
rect 20637 5525 20671 5559
rect 30389 5525 30423 5559
rect 30757 5525 30791 5559
rect 31217 5525 31251 5559
rect 1593 5321 1627 5355
rect 4537 5321 4571 5355
rect 6469 5321 6503 5355
rect 6929 5321 6963 5355
rect 8401 5321 8435 5355
rect 8769 5321 8803 5355
rect 10517 5321 10551 5355
rect 11897 5321 11931 5355
rect 12357 5321 12391 5355
rect 15485 5321 15519 5355
rect 20729 5321 20763 5355
rect 26341 5321 26375 5355
rect 27629 5321 27663 5355
rect 28457 5321 28491 5355
rect 29837 5321 29871 5355
rect 31033 5321 31067 5355
rect 5365 5253 5399 5287
rect 18429 5253 18463 5287
rect 20085 5253 20119 5287
rect 1409 5185 1443 5219
rect 2053 5185 2087 5219
rect 3801 5185 3835 5219
rect 5181 5185 5215 5219
rect 5273 5185 5307 5219
rect 5549 5185 5583 5219
rect 6837 5185 6871 5219
rect 10609 5185 10643 5219
rect 12265 5185 12299 5219
rect 15577 5185 15611 5219
rect 18245 5185 18279 5219
rect 18521 5185 18555 5219
rect 18613 5185 18647 5219
rect 3985 5117 4019 5151
rect 7021 5117 7055 5151
rect 8861 5117 8895 5151
rect 9045 5117 9079 5151
rect 10333 5117 10367 5151
rect 12449 5117 12483 5151
rect 15301 5117 15335 5151
rect 27721 5117 27755 5151
rect 27905 5117 27939 5151
rect 3617 4981 3651 5015
rect 4997 4981 5031 5015
rect 10977 4981 11011 5015
rect 15945 4981 15979 5015
rect 18797 4981 18831 5015
rect 27261 4981 27295 5015
rect 34713 4981 34747 5015
rect 4905 4777 4939 4811
rect 6837 4777 6871 4811
rect 15853 4777 15887 4811
rect 19717 4777 19751 4811
rect 23765 4777 23799 4811
rect 35265 4777 35299 4811
rect 36369 4777 36403 4811
rect 11069 4709 11103 4743
rect 12449 4709 12483 4743
rect 4077 4641 4111 4675
rect 6285 4641 6319 4675
rect 7481 4641 7515 4675
rect 14473 4641 14507 4675
rect 15209 4641 15243 4675
rect 20177 4641 20211 4675
rect 20361 4641 20395 4675
rect 25053 4641 25087 4675
rect 26801 4641 26835 4675
rect 28089 4641 28123 4675
rect 28273 4641 28307 4675
rect 35357 4641 35391 4675
rect 3249 4573 3283 4607
rect 4261 4573 4295 4607
rect 5733 4573 5767 4607
rect 7297 4573 7331 4607
rect 10517 4573 10551 4607
rect 10701 4573 10735 4607
rect 10885 4573 10919 4607
rect 11713 4573 11747 4607
rect 11897 4573 11931 4607
rect 14289 4573 14323 4607
rect 15485 4573 15519 4607
rect 18061 4573 18095 4607
rect 18245 4573 18279 4607
rect 20085 4573 20119 4607
rect 21005 4573 21039 4607
rect 26985 4573 27019 4607
rect 27169 4573 27203 4607
rect 28825 4573 28859 4607
rect 31033 4573 31067 4607
rect 34838 4573 34872 4607
rect 35942 4573 35976 4607
rect 36461 4573 36495 4607
rect 36921 4573 36955 4607
rect 37013 4573 37047 4607
rect 10793 4505 10827 4539
rect 15393 4505 15427 4539
rect 24869 4505 24903 4539
rect 27997 4505 28031 4539
rect 3065 4437 3099 4471
rect 4445 4437 4479 4471
rect 7205 4437 7239 4471
rect 11529 4437 11563 4471
rect 14105 4437 14139 4471
rect 17877 4437 17911 4471
rect 24409 4437 24443 4471
rect 24777 4437 24811 4471
rect 27629 4437 27663 4471
rect 29009 4437 29043 4471
rect 31217 4437 31251 4471
rect 34713 4437 34747 4471
rect 34897 4437 34931 4471
rect 35817 4437 35851 4471
rect 36001 4437 36035 4471
rect 4261 4233 4295 4267
rect 11529 4233 11563 4267
rect 12081 4233 12115 4267
rect 14657 4233 14691 4267
rect 15853 4233 15887 4267
rect 27997 4233 28031 4267
rect 1409 4097 1443 4131
rect 2053 4097 2087 4131
rect 3148 4097 3182 4131
rect 4905 4097 4939 4131
rect 7941 4097 7975 4131
rect 10517 4097 10551 4131
rect 13829 4097 13863 4131
rect 15393 4097 15427 4131
rect 15485 4097 15519 4131
rect 17325 4097 17359 4131
rect 19165 4097 19199 4131
rect 19349 4097 19383 4131
rect 19809 4097 19843 4131
rect 23489 4097 23523 4131
rect 23673 4097 23707 4131
rect 24685 4097 24719 4131
rect 27169 4097 27203 4131
rect 27353 4097 27387 4131
rect 29110 4097 29144 4131
rect 29377 4097 29411 4131
rect 29837 4097 29871 4131
rect 33885 4097 33919 4131
rect 34069 4097 34103 4131
rect 35164 4097 35198 4131
rect 2881 4029 2915 4063
rect 15209 4029 15243 4063
rect 18981 4029 19015 4063
rect 23029 4029 23063 4063
rect 23765 4029 23799 4063
rect 24869 4029 24903 4063
rect 34897 4029 34931 4063
rect 1593 3961 1627 3995
rect 4721 3893 4755 3927
rect 5457 3893 5491 3927
rect 7757 3893 7791 3927
rect 10701 3893 10735 3927
rect 13645 3893 13679 3927
rect 17509 3893 17543 3927
rect 19993 3893 20027 3927
rect 24501 3893 24535 3927
rect 27537 3893 27571 3927
rect 34069 3893 34103 3927
rect 36277 3893 36311 3927
rect 2789 3689 2823 3723
rect 16405 3689 16439 3723
rect 21005 3689 21039 3723
rect 22937 3689 22971 3723
rect 29653 3689 29687 3723
rect 30573 3689 30607 3723
rect 32505 3689 32539 3723
rect 35173 3689 35207 3723
rect 5181 3621 5215 3655
rect 9781 3621 9815 3655
rect 29009 3621 29043 3655
rect 2053 3553 2087 3587
rect 23397 3553 23431 3587
rect 23489 3553 23523 3587
rect 27629 3553 27663 3587
rect 31125 3553 31159 3587
rect 1409 3485 1443 3519
rect 2697 3485 2731 3519
rect 3801 3485 3835 3519
rect 10894 3485 10928 3519
rect 11161 3485 11195 3519
rect 17518 3485 17552 3519
rect 17785 3485 17819 3519
rect 18245 3485 18279 3519
rect 19625 3485 19659 3519
rect 19892 3485 19926 3519
rect 24593 3485 24627 3519
rect 34989 3485 35023 3519
rect 35173 3485 35207 3519
rect 4068 3417 4102 3451
rect 23305 3417 23339 3451
rect 27896 3417 27930 3451
rect 31370 3417 31404 3451
rect 1593 3349 1627 3383
rect 5733 3349 5767 3383
rect 11713 3349 11747 3383
rect 24409 3349 24443 3383
rect 8861 3145 8895 3179
rect 14565 3145 14599 3179
rect 22845 3145 22879 3179
rect 24777 3145 24811 3179
rect 27813 3145 27847 3179
rect 32781 3145 32815 3179
rect 34713 3145 34747 3179
rect 9505 3077 9539 3111
rect 15025 3077 15059 3111
rect 19441 3077 19475 3111
rect 23664 3077 23698 3111
rect 33600 3077 33634 3111
rect 1685 3009 1719 3043
rect 7481 3009 7515 3043
rect 7748 3009 7782 3043
rect 13185 3009 13219 3043
rect 13452 3009 13486 3043
rect 23397 3009 23431 3043
rect 27629 3009 27663 3043
rect 33333 3009 33367 3043
rect 1501 2873 1535 2907
rect 2605 2805 2639 2839
rect 3065 2805 3099 2839
rect 3709 2805 3743 2839
rect 2881 2601 2915 2635
rect 2697 2397 2731 2431
rect 37841 2397 37875 2431
rect 1869 2329 1903 2363
rect 2237 2329 2271 2363
rect 38025 2261 38059 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 38010 37448 38016 37460
rect 37971 37420 38016 37448
rect 38010 37408 38016 37420
rect 38068 37408 38074 37460
rect 29914 37204 29920 37256
rect 29972 37244 29978 37256
rect 30009 37247 30067 37253
rect 30009 37244 30021 37247
rect 29972 37216 30021 37244
rect 29972 37204 29978 37216
rect 30009 37213 30021 37216
rect 30055 37213 30067 37247
rect 37826 37244 37832 37256
rect 37787 37216 37832 37244
rect 30009 37207 30067 37213
rect 37826 37204 37832 37216
rect 37884 37204 37890 37256
rect 30190 37108 30196 37120
rect 30151 37080 30196 37108
rect 30190 37068 30196 37080
rect 30248 37068 30254 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 29914 36904 29920 36916
rect 29875 36876 29920 36904
rect 29914 36864 29920 36876
rect 29972 36864 29978 36916
rect 3970 36796 3976 36848
rect 4028 36836 4034 36848
rect 4028 36808 22094 36836
rect 4028 36796 4034 36808
rect 4065 36771 4123 36777
rect 4065 36737 4077 36771
rect 4111 36737 4123 36771
rect 12342 36768 12348 36780
rect 12303 36740 12348 36768
rect 4065 36731 4123 36737
rect 4080 36700 4108 36731
rect 12342 36728 12348 36740
rect 12400 36728 12406 36780
rect 16390 36700 16396 36712
rect 4080 36672 16396 36700
rect 16390 36660 16396 36672
rect 16448 36660 16454 36712
rect 17494 36700 17500 36712
rect 17455 36672 17500 36700
rect 17494 36660 17500 36672
rect 17552 36660 17558 36712
rect 17681 36703 17739 36709
rect 17681 36669 17693 36703
rect 17727 36700 17739 36703
rect 17954 36700 17960 36712
rect 17727 36672 17960 36700
rect 17727 36669 17739 36672
rect 17681 36663 17739 36669
rect 17954 36660 17960 36672
rect 18012 36660 18018 36712
rect 18046 36660 18052 36712
rect 18104 36700 18110 36712
rect 18104 36672 18149 36700
rect 18104 36660 18110 36672
rect 4062 36592 4068 36644
rect 4120 36632 4126 36644
rect 15194 36632 15200 36644
rect 4120 36604 15200 36632
rect 4120 36592 4126 36604
rect 15194 36592 15200 36604
rect 15252 36592 15258 36644
rect 22066 36632 22094 36808
rect 24578 36700 24584 36712
rect 24539 36672 24584 36700
rect 24578 36660 24584 36672
rect 24636 36660 24642 36712
rect 24762 36700 24768 36712
rect 24723 36672 24768 36700
rect 24762 36660 24768 36672
rect 24820 36660 24826 36712
rect 25041 36703 25099 36709
rect 25041 36669 25053 36703
rect 25087 36669 25099 36703
rect 25041 36663 25099 36669
rect 25056 36632 25084 36663
rect 27614 36632 27620 36644
rect 22066 36604 27620 36632
rect 27614 36592 27620 36604
rect 27672 36592 27678 36644
rect 3142 36564 3148 36576
rect 3103 36536 3148 36564
rect 3142 36524 3148 36536
rect 3200 36524 3206 36576
rect 3878 36564 3884 36576
rect 3839 36536 3884 36564
rect 3878 36524 3884 36536
rect 3936 36524 3942 36576
rect 4706 36564 4712 36576
rect 4667 36536 4712 36564
rect 4706 36524 4712 36536
rect 4764 36524 4770 36576
rect 8665 36567 8723 36573
rect 8665 36533 8677 36567
rect 8711 36564 8723 36567
rect 8938 36564 8944 36576
rect 8711 36536 8944 36564
rect 8711 36533 8723 36536
rect 8665 36527 8723 36533
rect 8938 36524 8944 36536
rect 8996 36524 9002 36576
rect 9122 36564 9128 36576
rect 9083 36536 9128 36564
rect 9122 36524 9128 36536
rect 9180 36524 9186 36576
rect 12529 36567 12587 36573
rect 12529 36533 12541 36567
rect 12575 36564 12587 36567
rect 12618 36564 12624 36576
rect 12575 36536 12624 36564
rect 12575 36533 12587 36536
rect 12529 36527 12587 36533
rect 12618 36524 12624 36536
rect 12676 36524 12682 36576
rect 19426 36524 19432 36576
rect 19484 36564 19490 36576
rect 20533 36567 20591 36573
rect 20533 36564 20545 36567
rect 19484 36536 20545 36564
rect 19484 36524 19490 36536
rect 20533 36533 20545 36536
rect 20579 36533 20591 36567
rect 20533 36527 20591 36533
rect 26602 36524 26608 36576
rect 26660 36564 26666 36576
rect 26973 36567 27031 36573
rect 26973 36564 26985 36567
rect 26660 36536 26985 36564
rect 26660 36524 26666 36536
rect 26973 36533 26985 36536
rect 27019 36533 27031 36567
rect 26973 36527 27031 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 12526 36360 12532 36372
rect 12487 36332 12532 36360
rect 12526 36320 12532 36332
rect 12584 36320 12590 36372
rect 17494 36360 17500 36372
rect 17455 36332 17500 36360
rect 17494 36320 17500 36332
rect 17552 36320 17558 36372
rect 17954 36360 17960 36372
rect 17915 36332 17960 36360
rect 17954 36320 17960 36332
rect 18012 36320 18018 36372
rect 24578 36320 24584 36372
rect 24636 36360 24642 36372
rect 25317 36363 25375 36369
rect 25317 36360 25329 36363
rect 24636 36332 25329 36360
rect 24636 36320 24642 36332
rect 25317 36329 25329 36332
rect 25363 36329 25375 36363
rect 25317 36323 25375 36329
rect 3786 36252 3792 36304
rect 3844 36292 3850 36304
rect 3844 36264 22232 36292
rect 3844 36252 3850 36264
rect 5258 36224 5264 36236
rect 5219 36196 5264 36224
rect 5258 36184 5264 36196
rect 5316 36184 5322 36236
rect 8938 36224 8944 36236
rect 8899 36196 8944 36224
rect 8938 36184 8944 36196
rect 8996 36184 9002 36236
rect 9766 36224 9772 36236
rect 9727 36196 9772 36224
rect 9766 36184 9772 36196
rect 9824 36184 9830 36236
rect 11977 36227 12035 36233
rect 11977 36193 11989 36227
rect 12023 36224 12035 36227
rect 12434 36224 12440 36236
rect 12023 36196 12440 36224
rect 12023 36193 12035 36196
rect 11977 36187 12035 36193
rect 12434 36184 12440 36196
rect 12492 36184 12498 36236
rect 12621 36227 12679 36233
rect 12621 36193 12633 36227
rect 12667 36224 12679 36227
rect 13814 36224 13820 36236
rect 12667 36196 13820 36224
rect 12667 36193 12679 36196
rect 12621 36187 12679 36193
rect 13814 36184 13820 36196
rect 13872 36184 13878 36236
rect 19426 36224 19432 36236
rect 19387 36196 19432 36224
rect 19426 36184 19432 36196
rect 19484 36184 19490 36236
rect 20898 36224 20904 36236
rect 20859 36196 20904 36224
rect 20898 36184 20904 36196
rect 20956 36184 20962 36236
rect 22204 36233 22232 36264
rect 22189 36227 22247 36233
rect 22189 36193 22201 36227
rect 22235 36224 22247 36227
rect 23566 36224 23572 36236
rect 22235 36196 23572 36224
rect 22235 36193 22247 36196
rect 22189 36187 22247 36193
rect 23566 36184 23572 36196
rect 23624 36184 23630 36236
rect 26602 36224 26608 36236
rect 26563 36196 26608 36224
rect 26602 36184 26608 36196
rect 26660 36184 26666 36236
rect 27614 36224 27620 36236
rect 27575 36196 27620 36224
rect 27614 36184 27620 36196
rect 27672 36184 27678 36236
rect 3237 36159 3295 36165
rect 3237 36125 3249 36159
rect 3283 36156 3295 36159
rect 3789 36159 3847 36165
rect 3789 36156 3801 36159
rect 3283 36128 3801 36156
rect 3283 36125 3295 36128
rect 3237 36119 3295 36125
rect 3789 36125 3801 36128
rect 3835 36125 3847 36159
rect 3789 36119 3847 36125
rect 7558 36116 7564 36168
rect 7616 36156 7622 36168
rect 7653 36159 7711 36165
rect 7653 36156 7665 36159
rect 7616 36128 7665 36156
rect 7616 36116 7622 36128
rect 7653 36125 7665 36128
rect 7699 36125 7711 36159
rect 7653 36119 7711 36125
rect 12713 36159 12771 36165
rect 12713 36125 12725 36159
rect 12759 36156 12771 36159
rect 12802 36156 12808 36168
rect 12759 36128 12808 36156
rect 12759 36125 12771 36128
rect 12713 36119 12771 36125
rect 12802 36116 12808 36128
rect 12860 36116 12866 36168
rect 13357 36159 13415 36165
rect 13357 36156 13369 36159
rect 12912 36128 13369 36156
rect 3326 36048 3332 36100
rect 3384 36088 3390 36100
rect 3973 36091 4031 36097
rect 3973 36088 3985 36091
rect 3384 36060 3985 36088
rect 3384 36048 3390 36060
rect 3973 36057 3985 36060
rect 4019 36057 4031 36091
rect 3973 36051 4031 36057
rect 9125 36091 9183 36097
rect 9125 36057 9137 36091
rect 9171 36088 9183 36091
rect 11974 36088 11980 36100
rect 9171 36060 11980 36088
rect 9171 36057 9183 36060
rect 9125 36051 9183 36057
rect 11974 36048 11980 36060
rect 12032 36048 12038 36100
rect 12437 36091 12495 36097
rect 12437 36057 12449 36091
rect 12483 36057 12495 36091
rect 12437 36051 12495 36057
rect 12452 36020 12480 36051
rect 12710 36020 12716 36032
rect 12452 35992 12716 36020
rect 12710 35980 12716 35992
rect 12768 35980 12774 36032
rect 12912 36029 12940 36128
rect 13357 36125 13369 36128
rect 13403 36125 13415 36159
rect 14090 36156 14096 36168
rect 14051 36128 14096 36156
rect 13357 36119 13415 36125
rect 14090 36116 14096 36128
rect 14148 36116 14154 36168
rect 16022 36156 16028 36168
rect 15983 36128 16028 36156
rect 16022 36116 16028 36128
rect 16080 36116 16086 36168
rect 18138 36156 18144 36168
rect 18099 36128 18144 36156
rect 18138 36116 18144 36128
rect 18196 36116 18202 36168
rect 21726 36156 21732 36168
rect 21687 36128 21732 36156
rect 21726 36116 21732 36128
rect 21784 36116 21790 36168
rect 24302 36116 24308 36168
rect 24360 36156 24366 36168
rect 24397 36159 24455 36165
rect 24397 36156 24409 36159
rect 24360 36128 24409 36156
rect 24360 36116 24366 36128
rect 24397 36125 24409 36128
rect 24443 36125 24455 36159
rect 26142 36156 26148 36168
rect 26103 36128 26148 36156
rect 24397 36119 24455 36125
rect 26142 36116 26148 36128
rect 26200 36116 26206 36168
rect 19613 36091 19671 36097
rect 19613 36057 19625 36091
rect 19659 36057 19671 36091
rect 21910 36088 21916 36100
rect 21871 36060 21916 36088
rect 19613 36051 19671 36057
rect 12897 36023 12955 36029
rect 12897 35989 12909 36023
rect 12943 35989 12955 36023
rect 13538 36020 13544 36032
rect 13499 35992 13544 36020
rect 12897 35983 12955 35989
rect 13538 35980 13544 35992
rect 13596 35980 13602 36032
rect 19426 35980 19432 36032
rect 19484 36020 19490 36032
rect 19628 36020 19656 36051
rect 21910 36048 21916 36060
rect 21968 36048 21974 36100
rect 26786 36088 26792 36100
rect 26747 36060 26792 36088
rect 26786 36048 26792 36060
rect 26844 36048 26850 36100
rect 19484 35992 19656 36020
rect 19484 35980 19490 35992
rect 20898 35980 20904 36032
rect 20956 36020 20962 36032
rect 25590 36020 25596 36032
rect 20956 35992 25596 36020
rect 20956 35980 20962 35992
rect 25590 35980 25596 35992
rect 25648 35980 25654 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 16850 35816 16856 35828
rect 11992 35788 16856 35816
rect 5258 35748 5264 35760
rect 5219 35720 5264 35748
rect 5258 35708 5264 35720
rect 5316 35708 5322 35760
rect 11992 35757 12020 35788
rect 16850 35776 16856 35788
rect 16908 35776 16914 35828
rect 19426 35776 19432 35828
rect 19484 35816 19490 35828
rect 19705 35819 19763 35825
rect 19705 35816 19717 35819
rect 19484 35788 19717 35816
rect 19484 35776 19490 35788
rect 19705 35785 19717 35788
rect 19751 35785 19763 35819
rect 19705 35779 19763 35785
rect 20809 35819 20867 35825
rect 20809 35785 20821 35819
rect 20855 35816 20867 35819
rect 21910 35816 21916 35828
rect 20855 35788 21916 35816
rect 20855 35785 20867 35788
rect 20809 35779 20867 35785
rect 21910 35776 21916 35788
rect 21968 35776 21974 35828
rect 11977 35751 12035 35757
rect 11977 35717 11989 35751
rect 12023 35717 12035 35751
rect 12618 35748 12624 35760
rect 12579 35720 12624 35748
rect 11977 35711 12035 35717
rect 12618 35708 12624 35720
rect 12676 35708 12682 35760
rect 15194 35708 15200 35760
rect 15252 35748 15258 35760
rect 20898 35748 20904 35760
rect 15252 35720 20904 35748
rect 15252 35708 15258 35720
rect 20898 35708 20904 35720
rect 20956 35708 20962 35760
rect 30024 35720 32168 35748
rect 7558 35680 7564 35692
rect 7519 35652 7564 35680
rect 7558 35640 7564 35652
rect 7616 35640 7622 35692
rect 10229 35683 10287 35689
rect 10229 35649 10241 35683
rect 10275 35680 10287 35683
rect 11514 35680 11520 35692
rect 10275 35652 11520 35680
rect 10275 35649 10287 35652
rect 10229 35643 10287 35649
rect 11514 35640 11520 35652
rect 11572 35640 11578 35692
rect 11701 35683 11759 35689
rect 11701 35649 11713 35683
rect 11747 35680 11759 35683
rect 12434 35680 12440 35692
rect 11747 35652 12112 35680
rect 12395 35652 12440 35680
rect 11747 35649 11759 35652
rect 11701 35643 11759 35649
rect 2961 35615 3019 35621
rect 2961 35581 2973 35615
rect 3007 35612 3019 35615
rect 3421 35615 3479 35621
rect 3421 35612 3433 35615
rect 3007 35584 3433 35612
rect 3007 35581 3019 35584
rect 2961 35575 3019 35581
rect 3421 35581 3433 35584
rect 3467 35581 3479 35615
rect 3421 35575 3479 35581
rect 3605 35615 3663 35621
rect 3605 35581 3617 35615
rect 3651 35612 3663 35615
rect 3786 35612 3792 35624
rect 3651 35584 3792 35612
rect 3651 35581 3663 35584
rect 3605 35575 3663 35581
rect 3786 35572 3792 35584
rect 3844 35572 3850 35624
rect 7745 35615 7803 35621
rect 7745 35581 7757 35615
rect 7791 35612 7803 35615
rect 8018 35612 8024 35624
rect 7791 35584 8024 35612
rect 7791 35581 7803 35584
rect 7745 35575 7803 35581
rect 8018 35572 8024 35584
rect 8076 35572 8082 35624
rect 9401 35615 9459 35621
rect 9401 35581 9413 35615
rect 9447 35612 9459 35615
rect 9766 35612 9772 35624
rect 9447 35584 9772 35612
rect 9447 35581 9459 35584
rect 9401 35575 9459 35581
rect 9766 35572 9772 35584
rect 9824 35572 9830 35624
rect 11882 35612 11888 35624
rect 11843 35584 11888 35612
rect 11882 35572 11888 35584
rect 11940 35572 11946 35624
rect 12084 35612 12112 35652
rect 12434 35640 12440 35652
rect 12492 35640 12498 35692
rect 15930 35680 15936 35692
rect 15891 35652 15936 35680
rect 15930 35640 15936 35652
rect 15988 35640 15994 35692
rect 16022 35640 16028 35692
rect 16080 35680 16086 35692
rect 16669 35683 16727 35689
rect 16669 35680 16681 35683
rect 16080 35652 16681 35680
rect 16080 35640 16086 35652
rect 16669 35649 16681 35652
rect 16715 35649 16727 35683
rect 16669 35643 16727 35649
rect 18966 35640 18972 35692
rect 19024 35680 19030 35692
rect 19521 35683 19579 35689
rect 19521 35680 19533 35683
rect 19024 35652 19533 35680
rect 19024 35640 19030 35652
rect 19521 35649 19533 35652
rect 19567 35649 19579 35683
rect 20622 35680 20628 35692
rect 20583 35652 20628 35680
rect 19521 35643 19579 35649
rect 20622 35640 20628 35652
rect 20680 35640 20686 35692
rect 21726 35640 21732 35692
rect 21784 35680 21790 35692
rect 21821 35683 21879 35689
rect 21821 35680 21833 35683
rect 21784 35652 21833 35680
rect 21784 35640 21790 35652
rect 21821 35649 21833 35652
rect 21867 35649 21879 35683
rect 21821 35643 21879 35649
rect 29546 35640 29552 35692
rect 29604 35680 29610 35692
rect 30024 35689 30052 35720
rect 30282 35689 30288 35692
rect 30009 35683 30067 35689
rect 30009 35680 30021 35683
rect 29604 35652 30021 35680
rect 29604 35640 29610 35652
rect 30009 35649 30021 35652
rect 30055 35649 30067 35683
rect 30009 35643 30067 35649
rect 30276 35643 30288 35689
rect 30340 35680 30346 35692
rect 30340 35652 30376 35680
rect 30282 35640 30288 35643
rect 30340 35640 30346 35652
rect 32140 35624 32168 35720
rect 32214 35640 32220 35692
rect 32272 35680 32278 35692
rect 32381 35683 32439 35689
rect 32381 35680 32393 35683
rect 32272 35652 32393 35680
rect 32272 35640 32278 35652
rect 32381 35649 32393 35652
rect 32427 35649 32439 35683
rect 32381 35643 32439 35649
rect 12802 35612 12808 35624
rect 12084 35584 12808 35612
rect 12802 35572 12808 35584
rect 12860 35572 12866 35624
rect 14185 35615 14243 35621
rect 14185 35581 14197 35615
rect 14231 35581 14243 35615
rect 14185 35575 14243 35581
rect 16853 35615 16911 35621
rect 16853 35581 16865 35615
rect 16899 35581 16911 35615
rect 18230 35612 18236 35624
rect 18191 35584 18236 35612
rect 16853 35575 16911 35581
rect 4062 35504 4068 35556
rect 4120 35544 4126 35556
rect 14200 35544 14228 35575
rect 4120 35516 14228 35544
rect 4120 35504 4126 35516
rect 9306 35436 9312 35488
rect 9364 35476 9370 35488
rect 10045 35479 10103 35485
rect 10045 35476 10057 35479
rect 9364 35448 10057 35476
rect 9364 35436 9370 35448
rect 10045 35445 10057 35448
rect 10091 35445 10103 35479
rect 10045 35439 10103 35445
rect 10134 35436 10140 35488
rect 10192 35476 10198 35488
rect 11517 35479 11575 35485
rect 11517 35476 11529 35479
rect 10192 35448 11529 35476
rect 10192 35436 10198 35448
rect 11517 35445 11529 35448
rect 11563 35445 11575 35479
rect 11517 35439 11575 35445
rect 11977 35479 12035 35485
rect 11977 35445 11989 35479
rect 12023 35476 12035 35479
rect 12526 35476 12532 35488
rect 12023 35448 12532 35476
rect 12023 35445 12035 35448
rect 11977 35439 12035 35445
rect 12526 35436 12532 35448
rect 12584 35436 12590 35488
rect 14200 35476 14228 35516
rect 16117 35547 16175 35553
rect 16117 35513 16129 35547
rect 16163 35544 16175 35547
rect 16868 35544 16896 35575
rect 18230 35572 18236 35584
rect 18288 35572 18294 35624
rect 23106 35612 23112 35624
rect 23067 35584 23112 35612
rect 23106 35572 23112 35584
rect 23164 35572 23170 35624
rect 23290 35612 23296 35624
rect 23251 35584 23296 35612
rect 23290 35572 23296 35584
rect 23348 35572 23354 35624
rect 23750 35612 23756 35624
rect 23711 35584 23756 35612
rect 23750 35572 23756 35584
rect 23808 35572 23814 35624
rect 26421 35615 26479 35621
rect 26421 35581 26433 35615
rect 26467 35612 26479 35615
rect 26973 35615 27031 35621
rect 26973 35612 26985 35615
rect 26467 35584 26985 35612
rect 26467 35581 26479 35584
rect 26421 35575 26479 35581
rect 26973 35581 26985 35584
rect 27019 35581 27031 35615
rect 27154 35612 27160 35624
rect 27115 35584 27160 35612
rect 26973 35575 27031 35581
rect 27154 35572 27160 35584
rect 27212 35572 27218 35624
rect 27614 35572 27620 35624
rect 27672 35612 27678 35624
rect 28350 35612 28356 35624
rect 27672 35584 28356 35612
rect 27672 35572 27678 35584
rect 28350 35572 28356 35584
rect 28408 35572 28414 35624
rect 32122 35612 32128 35624
rect 32083 35584 32128 35612
rect 32122 35572 32128 35584
rect 32180 35572 32186 35624
rect 16163 35516 16896 35544
rect 16163 35513 16175 35516
rect 16117 35507 16175 35513
rect 14274 35476 14280 35488
rect 14187 35448 14280 35476
rect 14274 35436 14280 35448
rect 14332 35476 14338 35488
rect 18046 35476 18052 35488
rect 14332 35448 18052 35476
rect 14332 35436 14338 35448
rect 18046 35436 18052 35448
rect 18104 35476 18110 35488
rect 18322 35476 18328 35488
rect 18104 35448 18328 35476
rect 18104 35436 18110 35448
rect 18322 35436 18328 35448
rect 18380 35436 18386 35488
rect 21910 35436 21916 35488
rect 21968 35476 21974 35488
rect 22465 35479 22523 35485
rect 22465 35476 22477 35479
rect 21968 35448 22477 35476
rect 21968 35436 21974 35448
rect 22465 35445 22477 35448
rect 22511 35445 22523 35479
rect 22465 35439 22523 35445
rect 29914 35436 29920 35488
rect 29972 35476 29978 35488
rect 31389 35479 31447 35485
rect 31389 35476 31401 35479
rect 29972 35448 31401 35476
rect 29972 35436 29978 35448
rect 31389 35445 31401 35448
rect 31435 35445 31447 35479
rect 33502 35476 33508 35488
rect 33463 35448 33508 35476
rect 31389 35439 31447 35445
rect 33502 35436 33508 35448
rect 33560 35436 33566 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 3237 35275 3295 35281
rect 3237 35241 3249 35275
rect 3283 35272 3295 35275
rect 3326 35272 3332 35284
rect 3283 35244 3332 35272
rect 3283 35241 3295 35244
rect 3237 35235 3295 35241
rect 3326 35232 3332 35244
rect 3384 35232 3390 35284
rect 3786 35272 3792 35284
rect 3747 35244 3792 35272
rect 3786 35232 3792 35244
rect 3844 35232 3850 35284
rect 8018 35272 8024 35284
rect 7979 35244 8024 35272
rect 8018 35232 8024 35244
rect 8076 35232 8082 35284
rect 12342 35232 12348 35284
rect 12400 35272 12406 35284
rect 12713 35275 12771 35281
rect 12713 35272 12725 35275
rect 12400 35244 12725 35272
rect 12400 35232 12406 35244
rect 12713 35241 12725 35244
rect 12759 35241 12771 35275
rect 12713 35235 12771 35241
rect 12897 35275 12955 35281
rect 12897 35241 12909 35275
rect 12943 35241 12955 35275
rect 16390 35272 16396 35284
rect 16351 35244 16396 35272
rect 12897 35235 12955 35241
rect 10134 35204 10140 35216
rect 3068 35176 10140 35204
rect 3068 35077 3096 35176
rect 10134 35164 10140 35176
rect 10192 35164 10198 35216
rect 12526 35164 12532 35216
rect 12584 35204 12590 35216
rect 12912 35204 12940 35235
rect 16390 35232 16396 35244
rect 16448 35232 16454 35284
rect 16853 35275 16911 35281
rect 16853 35241 16865 35275
rect 16899 35272 16911 35275
rect 17770 35272 17776 35284
rect 16899 35244 17776 35272
rect 16899 35241 16911 35244
rect 16853 35235 16911 35241
rect 17770 35232 17776 35244
rect 17828 35232 17834 35284
rect 18233 35275 18291 35281
rect 18233 35241 18245 35275
rect 18279 35272 18291 35275
rect 20622 35272 20628 35284
rect 18279 35244 20628 35272
rect 18279 35241 18291 35244
rect 18233 35235 18291 35241
rect 20622 35232 20628 35244
rect 20680 35232 20686 35284
rect 26053 35275 26111 35281
rect 26053 35241 26065 35275
rect 26099 35272 26111 35275
rect 26786 35272 26792 35284
rect 26099 35244 26792 35272
rect 26099 35241 26111 35244
rect 26053 35235 26111 35241
rect 26786 35232 26792 35244
rect 26844 35232 26850 35284
rect 32125 35275 32183 35281
rect 32125 35241 32137 35275
rect 32171 35272 32183 35275
rect 32214 35272 32220 35284
rect 32171 35244 32220 35272
rect 32171 35241 32183 35244
rect 32125 35235 32183 35241
rect 32214 35232 32220 35244
rect 32272 35232 32278 35284
rect 13814 35204 13820 35216
rect 12584 35176 12940 35204
rect 13096 35176 13820 35204
rect 12584 35164 12590 35176
rect 5994 35136 6000 35148
rect 3988 35108 6000 35136
rect 3988 35077 4016 35108
rect 5994 35096 6000 35108
rect 6052 35096 6058 35148
rect 6089 35139 6147 35145
rect 6089 35105 6101 35139
rect 6135 35136 6147 35139
rect 7009 35139 7067 35145
rect 7009 35136 7021 35139
rect 6135 35108 7021 35136
rect 6135 35105 6147 35108
rect 6089 35099 6147 35105
rect 7009 35105 7021 35108
rect 7055 35105 7067 35139
rect 9122 35136 9128 35148
rect 9083 35108 9128 35136
rect 7009 35099 7067 35105
rect 9122 35096 9128 35108
rect 9180 35096 9186 35148
rect 9306 35136 9312 35148
rect 9267 35108 9312 35136
rect 9306 35096 9312 35108
rect 9364 35096 9370 35148
rect 10505 35139 10563 35145
rect 10505 35105 10517 35139
rect 10551 35105 10563 35139
rect 11974 35136 11980 35148
rect 11935 35108 11980 35136
rect 10505 35099 10563 35105
rect 3053 35071 3111 35077
rect 3053 35037 3065 35071
rect 3099 35037 3111 35071
rect 3053 35031 3111 35037
rect 3973 35071 4031 35077
rect 3973 35037 3985 35071
rect 4019 35037 4031 35071
rect 3973 35031 4031 35037
rect 6273 35071 6331 35077
rect 6273 35037 6285 35071
rect 6319 35037 6331 35071
rect 6730 35068 6736 35080
rect 6691 35040 6736 35068
rect 6273 35031 6331 35037
rect 4338 34960 4344 35012
rect 4396 35000 4402 35012
rect 4433 35003 4491 35009
rect 4433 35000 4445 35003
rect 4396 34972 4445 35000
rect 4396 34960 4402 34972
rect 4433 34969 4445 34972
rect 4479 34969 4491 35003
rect 4433 34963 4491 34969
rect 4706 34960 4712 35012
rect 4764 35000 4770 35012
rect 6288 35000 6316 35031
rect 6730 35028 6736 35040
rect 6788 35028 6794 35080
rect 8110 35028 8116 35080
rect 8168 35068 8174 35080
rect 8205 35071 8263 35077
rect 8205 35068 8217 35071
rect 8168 35040 8217 35068
rect 8168 35028 8174 35040
rect 8205 35037 8217 35040
rect 8251 35037 8263 35071
rect 8205 35031 8263 35037
rect 10520 35000 10548 35099
rect 11974 35096 11980 35108
rect 12032 35096 12038 35148
rect 13096 35145 13124 35176
rect 13814 35164 13820 35176
rect 13872 35204 13878 35216
rect 14642 35204 14648 35216
rect 13872 35176 14648 35204
rect 13872 35164 13878 35176
rect 14642 35164 14648 35176
rect 14700 35164 14706 35216
rect 13081 35139 13139 35145
rect 13081 35136 13093 35139
rect 12636 35108 13093 35136
rect 12253 35071 12311 35077
rect 12253 35037 12265 35071
rect 12299 35068 12311 35071
rect 12434 35068 12440 35080
rect 12299 35040 12440 35068
rect 12299 35037 12311 35040
rect 12253 35031 12311 35037
rect 12434 35028 12440 35040
rect 12492 35028 12498 35080
rect 4764 34972 6316 35000
rect 10428 34972 10548 35000
rect 4764 34960 4770 34972
rect 4062 34892 4068 34944
rect 4120 34932 4126 34944
rect 10428 34932 10456 34972
rect 11790 34960 11796 35012
rect 11848 35000 11854 35012
rect 12636 35000 12664 35108
rect 13081 35105 13093 35108
rect 13127 35105 13139 35139
rect 14090 35136 14096 35148
rect 14051 35108 14096 35136
rect 13081 35099 13139 35105
rect 14090 35096 14096 35108
rect 14148 35096 14154 35148
rect 15194 35136 15200 35148
rect 15155 35108 15200 35136
rect 15194 35096 15200 35108
rect 15252 35096 15258 35148
rect 17954 35136 17960 35148
rect 16592 35108 17816 35136
rect 17915 35108 17960 35136
rect 16592 35080 16620 35108
rect 12802 35028 12808 35080
rect 12860 35068 12866 35080
rect 12897 35071 12955 35077
rect 12897 35068 12909 35071
rect 12860 35040 12909 35068
rect 12860 35028 12866 35040
rect 12897 35037 12909 35040
rect 12943 35037 12955 35071
rect 16574 35068 16580 35080
rect 16535 35040 16580 35068
rect 12897 35031 12955 35037
rect 16574 35028 16580 35040
rect 16632 35028 16638 35080
rect 16666 35028 16672 35080
rect 16724 35068 16730 35080
rect 16724 35040 16769 35068
rect 16724 35028 16730 35040
rect 16850 35028 16856 35080
rect 16908 35068 16914 35080
rect 17788 35068 17816 35108
rect 17954 35096 17960 35108
rect 18012 35096 18018 35148
rect 21910 35136 21916 35148
rect 21871 35108 21916 35136
rect 21910 35096 21916 35108
rect 21968 35096 21974 35148
rect 23750 35136 23756 35148
rect 23711 35108 23756 35136
rect 23750 35096 23756 35108
rect 23808 35136 23814 35148
rect 24578 35136 24584 35148
rect 23808 35108 24584 35136
rect 23808 35096 23814 35108
rect 24578 35096 24584 35108
rect 24636 35096 24642 35148
rect 24673 35139 24731 35145
rect 24673 35105 24685 35139
rect 24719 35136 24731 35139
rect 24762 35136 24768 35148
rect 24719 35108 24768 35136
rect 24719 35105 24731 35108
rect 24673 35099 24731 35105
rect 24762 35096 24768 35108
rect 24820 35096 24826 35148
rect 26142 35096 26148 35148
rect 26200 35136 26206 35148
rect 26697 35139 26755 35145
rect 26697 35136 26709 35139
rect 26200 35108 26709 35136
rect 26200 35096 26206 35108
rect 26697 35105 26709 35108
rect 26743 35105 26755 35139
rect 28350 35136 28356 35148
rect 28311 35108 28356 35136
rect 26697 35099 26755 35105
rect 28350 35096 28356 35108
rect 28408 35096 28414 35148
rect 29546 35136 29552 35148
rect 29507 35108 29552 35136
rect 29546 35096 29552 35108
rect 29604 35096 29610 35148
rect 17862 35068 17868 35080
rect 16908 35040 16953 35068
rect 17775 35040 17868 35068
rect 16908 35028 16914 35040
rect 17862 35028 17868 35040
rect 17920 35068 17926 35080
rect 18049 35071 18107 35077
rect 18049 35068 18061 35071
rect 17920 35040 18061 35068
rect 17920 35028 17926 35040
rect 18049 35037 18061 35040
rect 18095 35068 18107 35071
rect 18782 35068 18788 35080
rect 18095 35040 18788 35068
rect 18095 35037 18107 35040
rect 18049 35031 18107 35037
rect 18782 35028 18788 35040
rect 18840 35028 18846 35080
rect 23474 35028 23480 35080
rect 23532 35068 23538 35080
rect 24397 35071 24455 35077
rect 24397 35068 24409 35071
rect 23532 35040 24409 35068
rect 23532 35028 23538 35040
rect 24397 35037 24409 35040
rect 24443 35037 24455 35071
rect 25866 35068 25872 35080
rect 25827 35040 25872 35068
rect 24397 35031 24455 35037
rect 25866 35028 25872 35040
rect 25924 35028 25930 35080
rect 31938 35068 31944 35080
rect 31899 35040 31944 35068
rect 31938 35028 31944 35040
rect 31996 35028 32002 35080
rect 11848 34972 12664 35000
rect 11848 34960 11854 34972
rect 12710 34960 12716 35012
rect 12768 35000 12774 35012
rect 13173 35003 13231 35009
rect 13173 35000 13185 35003
rect 12768 34972 13185 35000
rect 12768 34960 12774 34972
rect 13173 34969 13185 34972
rect 13219 34969 13231 35003
rect 13173 34963 13231 34969
rect 13538 34960 13544 35012
rect 13596 35000 13602 35012
rect 14277 35003 14335 35009
rect 14277 35000 14289 35003
rect 13596 34972 14289 35000
rect 13596 34960 13602 34972
rect 14277 34969 14289 34972
rect 14323 34969 14335 35003
rect 14277 34963 14335 34969
rect 17310 34960 17316 35012
rect 17368 35000 17374 35012
rect 17773 35003 17831 35009
rect 17773 35000 17785 35003
rect 17368 34972 17785 35000
rect 17368 34960 17374 34972
rect 17773 34969 17785 34972
rect 17819 34969 17831 35003
rect 17773 34963 17831 34969
rect 21174 34960 21180 35012
rect 21232 35000 21238 35012
rect 22097 35003 22155 35009
rect 22097 35000 22109 35003
rect 21232 34972 22109 35000
rect 21232 34960 21238 34972
rect 22097 34969 22109 34972
rect 22143 34969 22155 35003
rect 26878 35000 26884 35012
rect 26839 34972 26884 35000
rect 22097 34963 22155 34969
rect 26878 34960 26884 34972
rect 26936 34960 26942 35012
rect 29822 35009 29828 35012
rect 29816 34963 29828 35009
rect 29880 35000 29886 35012
rect 29880 34972 29916 35000
rect 29822 34960 29828 34963
rect 29880 34960 29886 34972
rect 18230 34932 18236 34944
rect 4120 34904 18236 34932
rect 4120 34892 4126 34904
rect 18230 34892 18236 34904
rect 18288 34892 18294 34944
rect 30098 34892 30104 34944
rect 30156 34932 30162 34944
rect 30929 34935 30987 34941
rect 30929 34932 30941 34935
rect 30156 34904 30941 34932
rect 30156 34892 30162 34904
rect 30929 34901 30941 34904
rect 30975 34901 30987 34935
rect 30929 34895 30987 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 6730 34728 6736 34740
rect 6691 34700 6736 34728
rect 6730 34688 6736 34700
rect 6788 34688 6794 34740
rect 8110 34728 8116 34740
rect 8071 34700 8116 34728
rect 8110 34688 8116 34700
rect 8168 34688 8174 34740
rect 11514 34728 11520 34740
rect 11475 34700 11520 34728
rect 11514 34688 11520 34700
rect 11572 34688 11578 34740
rect 12434 34688 12440 34740
rect 12492 34728 12498 34740
rect 13357 34731 13415 34737
rect 12492 34700 12537 34728
rect 12492 34688 12498 34700
rect 13357 34697 13369 34731
rect 13403 34697 13415 34731
rect 13357 34691 13415 34697
rect 3329 34663 3387 34669
rect 3329 34629 3341 34663
rect 3375 34660 3387 34663
rect 3878 34660 3884 34672
rect 3375 34632 3884 34660
rect 3375 34629 3387 34632
rect 3329 34623 3387 34629
rect 3878 34620 3884 34632
rect 3936 34620 3942 34672
rect 7193 34663 7251 34669
rect 7193 34629 7205 34663
rect 7239 34660 7251 34663
rect 7653 34663 7711 34669
rect 7653 34660 7665 34663
rect 7239 34632 7665 34660
rect 7239 34629 7251 34632
rect 7193 34623 7251 34629
rect 7653 34629 7665 34632
rect 7699 34660 7711 34663
rect 8018 34660 8024 34672
rect 7699 34632 8024 34660
rect 7699 34629 7711 34632
rect 7653 34623 7711 34629
rect 8018 34620 8024 34632
rect 8076 34620 8082 34672
rect 12802 34660 12808 34672
rect 11716 34632 12434 34660
rect 3142 34592 3148 34604
rect 3103 34564 3148 34592
rect 3142 34552 3148 34564
rect 3200 34552 3206 34604
rect 6917 34595 6975 34601
rect 6917 34561 6929 34595
rect 6963 34592 6975 34595
rect 7466 34592 7472 34604
rect 6963 34564 7472 34592
rect 6963 34561 6975 34564
rect 6917 34555 6975 34561
rect 7466 34552 7472 34564
rect 7524 34592 7530 34604
rect 11716 34601 11744 34632
rect 7929 34595 7987 34601
rect 7929 34592 7941 34595
rect 7524 34564 7941 34592
rect 7524 34552 7530 34564
rect 7929 34561 7941 34564
rect 7975 34561 7987 34595
rect 7929 34555 7987 34561
rect 11701 34595 11759 34601
rect 11701 34561 11713 34595
rect 11747 34561 11759 34595
rect 11701 34555 11759 34561
rect 11790 34552 11796 34604
rect 11848 34592 11854 34604
rect 11848 34564 11893 34592
rect 11848 34552 11854 34564
rect 11974 34552 11980 34604
rect 12032 34592 12038 34604
rect 12406 34592 12434 34632
rect 12636 34632 12808 34660
rect 12636 34601 12664 34632
rect 12802 34620 12808 34632
rect 12860 34660 12866 34672
rect 13372 34660 13400 34691
rect 15930 34688 15936 34740
rect 15988 34728 15994 34740
rect 16669 34731 16727 34737
rect 16669 34728 16681 34731
rect 15988 34700 16681 34728
rect 15988 34688 15994 34700
rect 16669 34697 16681 34700
rect 16715 34697 16727 34731
rect 16669 34691 16727 34697
rect 16850 34688 16856 34740
rect 16908 34688 16914 34740
rect 18046 34688 18052 34740
rect 18104 34728 18110 34740
rect 18966 34728 18972 34740
rect 18104 34700 18149 34728
rect 18927 34700 18972 34728
rect 18104 34688 18110 34700
rect 18966 34688 18972 34700
rect 19024 34688 19030 34740
rect 21174 34728 21180 34740
rect 21135 34700 21180 34728
rect 21174 34688 21180 34700
rect 21232 34688 21238 34740
rect 29822 34728 29828 34740
rect 29783 34700 29828 34728
rect 29822 34688 29828 34700
rect 29880 34688 29886 34740
rect 30282 34728 30288 34740
rect 30243 34700 30288 34728
rect 30282 34688 30288 34700
rect 30340 34688 30346 34740
rect 12860 34632 13400 34660
rect 16868 34660 16896 34688
rect 16868 34632 17172 34660
rect 12860 34620 12866 34632
rect 12621 34595 12679 34601
rect 12621 34592 12633 34595
rect 12032 34564 12077 34592
rect 12406 34564 12633 34592
rect 12032 34552 12038 34564
rect 12621 34561 12633 34564
rect 12667 34561 12679 34595
rect 12894 34592 12900 34604
rect 12855 34564 12900 34592
rect 12621 34555 12679 34561
rect 12894 34552 12900 34564
rect 12952 34552 12958 34604
rect 13538 34592 13544 34604
rect 13451 34564 13544 34592
rect 13538 34552 13544 34564
rect 13596 34592 13602 34604
rect 15930 34592 15936 34604
rect 13596 34564 15936 34592
rect 13596 34552 13602 34564
rect 15930 34552 15936 34564
rect 15988 34552 15994 34604
rect 16114 34552 16120 34604
rect 16172 34592 16178 34604
rect 16574 34592 16580 34604
rect 16172 34564 16580 34592
rect 16172 34552 16178 34564
rect 16574 34552 16580 34564
rect 16632 34592 16638 34604
rect 17144 34601 17172 34632
rect 32122 34620 32128 34672
rect 32180 34660 32186 34672
rect 34790 34660 34796 34672
rect 32180 34632 34796 34660
rect 32180 34620 32186 34632
rect 16853 34595 16911 34601
rect 16853 34592 16865 34595
rect 16632 34564 16865 34592
rect 16632 34552 16638 34564
rect 16853 34561 16865 34564
rect 16899 34561 16911 34595
rect 16853 34555 16911 34561
rect 17129 34595 17187 34601
rect 17129 34561 17141 34595
rect 17175 34592 17187 34595
rect 17589 34595 17647 34601
rect 17589 34592 17601 34595
rect 17175 34564 17601 34592
rect 17175 34561 17187 34564
rect 17129 34555 17187 34561
rect 17589 34561 17601 34564
rect 17635 34592 17647 34595
rect 17635 34564 17816 34592
rect 17635 34561 17647 34564
rect 17589 34555 17647 34561
rect 4338 34524 4344 34536
rect 4299 34496 4344 34524
rect 4338 34484 4344 34496
rect 4396 34524 4402 34536
rect 4614 34524 4620 34536
rect 4396 34496 4620 34524
rect 4396 34484 4402 34496
rect 4614 34484 4620 34496
rect 4672 34484 4678 34536
rect 7101 34527 7159 34533
rect 7101 34493 7113 34527
rect 7147 34524 7159 34527
rect 7837 34527 7895 34533
rect 7837 34524 7849 34527
rect 7147 34496 7849 34524
rect 7147 34493 7159 34496
rect 7101 34487 7159 34493
rect 7837 34493 7849 34496
rect 7883 34493 7895 34527
rect 7837 34487 7895 34493
rect 4062 34416 4068 34468
rect 4120 34456 4126 34468
rect 4356 34456 4384 34484
rect 7852 34456 7880 34487
rect 11882 34484 11888 34536
rect 11940 34524 11946 34536
rect 12713 34527 12771 34533
rect 12713 34524 12725 34527
rect 11940 34496 12725 34524
rect 11940 34484 11946 34496
rect 12713 34493 12725 34496
rect 12759 34524 12771 34527
rect 16666 34524 16672 34536
rect 12759 34496 16672 34524
rect 12759 34493 12771 34496
rect 12713 34487 12771 34493
rect 16666 34484 16672 34496
rect 16724 34524 16730 34536
rect 16942 34524 16948 34536
rect 16724 34496 16948 34524
rect 16724 34484 16730 34496
rect 16942 34484 16948 34496
rect 17000 34484 17006 34536
rect 17678 34524 17684 34536
rect 17639 34496 17684 34524
rect 17678 34484 17684 34496
rect 17736 34484 17742 34536
rect 17788 34524 17816 34564
rect 17862 34552 17868 34604
rect 17920 34601 17926 34604
rect 17920 34595 17939 34601
rect 17927 34561 17939 34595
rect 18509 34595 18567 34601
rect 18509 34592 18521 34595
rect 17920 34555 17939 34561
rect 18248 34564 18521 34592
rect 17920 34552 17926 34555
rect 18046 34524 18052 34536
rect 17788 34496 18052 34524
rect 18046 34484 18052 34496
rect 18104 34484 18110 34536
rect 18138 34484 18144 34536
rect 18196 34524 18202 34536
rect 18248 34524 18276 34564
rect 18509 34561 18521 34564
rect 18555 34561 18567 34595
rect 18782 34592 18788 34604
rect 18743 34564 18788 34592
rect 18509 34555 18567 34561
rect 18782 34552 18788 34564
rect 18840 34552 18846 34604
rect 20162 34552 20168 34604
rect 20220 34592 20226 34604
rect 20993 34595 21051 34601
rect 20993 34592 21005 34595
rect 20220 34564 21005 34592
rect 20220 34552 20226 34564
rect 20993 34561 21005 34564
rect 21039 34561 21051 34595
rect 24302 34592 24308 34604
rect 24263 34564 24308 34592
rect 20993 34555 21051 34561
rect 24302 34552 24308 34564
rect 24360 34552 24366 34604
rect 29638 34592 29644 34604
rect 29599 34564 29644 34592
rect 29638 34552 29644 34564
rect 29696 34552 29702 34604
rect 30466 34592 30472 34604
rect 30427 34564 30472 34592
rect 30466 34552 30472 34564
rect 30524 34552 30530 34604
rect 32968 34601 32996 34632
rect 34790 34620 34796 34632
rect 34848 34620 34854 34672
rect 33226 34601 33232 34604
rect 32953 34595 33011 34601
rect 32953 34561 32965 34595
rect 32999 34561 33011 34595
rect 32953 34555 33011 34561
rect 33220 34555 33232 34601
rect 33284 34592 33290 34604
rect 33284 34564 33320 34592
rect 33226 34552 33232 34555
rect 33284 34552 33290 34564
rect 18598 34524 18604 34536
rect 18196 34496 18276 34524
rect 18559 34496 18604 34524
rect 18196 34484 18202 34496
rect 18598 34484 18604 34496
rect 18656 34484 18662 34536
rect 21818 34524 21824 34536
rect 21779 34496 21824 34524
rect 21818 34484 21824 34496
rect 21876 34484 21882 34536
rect 22002 34524 22008 34536
rect 21963 34496 22008 34524
rect 22002 34484 22008 34496
rect 22060 34484 22066 34536
rect 22281 34527 22339 34533
rect 22281 34493 22293 34527
rect 22327 34493 22339 34527
rect 24486 34524 24492 34536
rect 24447 34496 24492 34524
rect 22281 34487 22339 34493
rect 7926 34456 7932 34468
rect 4120 34428 4384 34456
rect 4448 34428 7788 34456
rect 7852 34428 7932 34456
rect 4120 34416 4126 34428
rect 2685 34391 2743 34397
rect 2685 34357 2697 34391
rect 2731 34388 2743 34391
rect 2774 34388 2780 34400
rect 2731 34360 2780 34388
rect 2731 34357 2743 34360
rect 2685 34351 2743 34357
rect 2774 34348 2780 34360
rect 2832 34348 2838 34400
rect 3694 34348 3700 34400
rect 3752 34388 3758 34400
rect 4448 34388 4476 34428
rect 3752 34360 4476 34388
rect 5629 34391 5687 34397
rect 3752 34348 3758 34360
rect 5629 34357 5641 34391
rect 5675 34388 5687 34391
rect 6270 34388 6276 34400
rect 5675 34360 6276 34388
rect 5675 34357 5687 34360
rect 5629 34351 5687 34357
rect 6270 34348 6276 34360
rect 6328 34348 6334 34400
rect 7193 34391 7251 34397
rect 7193 34357 7205 34391
rect 7239 34388 7251 34391
rect 7650 34388 7656 34400
rect 7239 34360 7656 34388
rect 7239 34357 7251 34360
rect 7193 34351 7251 34357
rect 7650 34348 7656 34360
rect 7708 34348 7714 34400
rect 7760 34388 7788 34428
rect 7926 34416 7932 34428
rect 7984 34416 7990 34468
rect 14458 34456 14464 34468
rect 8036 34428 14464 34456
rect 8036 34388 8064 34428
rect 14458 34416 14464 34428
rect 14516 34416 14522 34468
rect 18414 34416 18420 34468
rect 18472 34456 18478 34468
rect 22296 34456 22324 34487
rect 24486 34484 24492 34496
rect 24544 34484 24550 34536
rect 24578 34484 24584 34536
rect 24636 34524 24642 34536
rect 24765 34527 24823 34533
rect 24765 34524 24777 34527
rect 24636 34496 24777 34524
rect 24636 34484 24642 34496
rect 24765 34493 24777 34496
rect 24811 34493 24823 34527
rect 24765 34487 24823 34493
rect 23658 34456 23664 34468
rect 18472 34428 23664 34456
rect 18472 34416 18478 34428
rect 23658 34416 23664 34428
rect 23716 34416 23722 34468
rect 7760 34360 8064 34388
rect 11977 34391 12035 34397
rect 11977 34357 11989 34391
rect 12023 34388 12035 34391
rect 12526 34388 12532 34400
rect 12023 34360 12532 34388
rect 12023 34357 12035 34360
rect 11977 34351 12035 34357
rect 12526 34348 12532 34360
rect 12584 34388 12590 34400
rect 12621 34391 12679 34397
rect 12621 34388 12633 34391
rect 12584 34360 12633 34388
rect 12584 34348 12590 34360
rect 12621 34357 12633 34360
rect 12667 34357 12679 34391
rect 16114 34388 16120 34400
rect 16075 34360 16120 34388
rect 12621 34351 12679 34357
rect 16114 34348 16120 34360
rect 16172 34348 16178 34400
rect 17126 34388 17132 34400
rect 17039 34360 17132 34388
rect 17126 34348 17132 34360
rect 17184 34388 17190 34400
rect 17770 34388 17776 34400
rect 17184 34360 17776 34388
rect 17184 34348 17190 34360
rect 17770 34348 17776 34360
rect 17828 34388 17834 34400
rect 17865 34391 17923 34397
rect 17865 34388 17877 34391
rect 17828 34360 17877 34388
rect 17828 34348 17834 34360
rect 17865 34357 17877 34360
rect 17911 34388 17923 34391
rect 18509 34391 18567 34397
rect 18509 34388 18521 34391
rect 17911 34360 18521 34388
rect 17911 34357 17923 34360
rect 17865 34351 17923 34357
rect 18509 34357 18521 34360
rect 18555 34357 18567 34391
rect 18509 34351 18567 34357
rect 19334 34348 19340 34400
rect 19392 34388 19398 34400
rect 19429 34391 19487 34397
rect 19429 34388 19441 34391
rect 19392 34360 19441 34388
rect 19392 34348 19398 34360
rect 19429 34357 19441 34360
rect 19475 34357 19487 34391
rect 34330 34388 34336 34400
rect 34291 34360 34336 34388
rect 19429 34351 19487 34357
rect 34330 34348 34336 34360
rect 34388 34348 34394 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 5994 34144 6000 34196
rect 6052 34184 6058 34196
rect 7285 34187 7343 34193
rect 7285 34184 7297 34187
rect 6052 34156 7297 34184
rect 6052 34144 6058 34156
rect 7285 34153 7297 34156
rect 7331 34153 7343 34187
rect 7742 34184 7748 34196
rect 7703 34156 7748 34184
rect 7285 34147 7343 34153
rect 7742 34144 7748 34156
rect 7800 34144 7806 34196
rect 12526 34144 12532 34196
rect 12584 34184 12590 34196
rect 13081 34187 13139 34193
rect 13081 34184 13093 34187
rect 12584 34156 13093 34184
rect 12584 34144 12590 34156
rect 13081 34153 13093 34156
rect 13127 34153 13139 34187
rect 13081 34147 13139 34153
rect 15657 34187 15715 34193
rect 15657 34153 15669 34187
rect 15703 34184 15715 34187
rect 17313 34187 17371 34193
rect 17313 34184 17325 34187
rect 15703 34156 17325 34184
rect 15703 34153 15715 34156
rect 15657 34147 15715 34153
rect 17313 34153 17325 34156
rect 17359 34184 17371 34187
rect 18233 34187 18291 34193
rect 18233 34184 18245 34187
rect 17359 34156 18245 34184
rect 17359 34153 17371 34156
rect 17313 34147 17371 34153
rect 18233 34153 18245 34156
rect 18279 34184 18291 34187
rect 18598 34184 18604 34196
rect 18279 34156 18604 34184
rect 18279 34153 18291 34156
rect 18233 34147 18291 34153
rect 18598 34144 18604 34156
rect 18656 34184 18662 34196
rect 19245 34187 19303 34193
rect 19245 34184 19257 34187
rect 18656 34156 19257 34184
rect 18656 34144 18662 34156
rect 19245 34153 19257 34156
rect 19291 34153 19303 34187
rect 21818 34184 21824 34196
rect 21779 34156 21824 34184
rect 19245 34147 19303 34153
rect 21818 34144 21824 34156
rect 21876 34144 21882 34196
rect 23106 34144 23112 34196
rect 23164 34184 23170 34196
rect 23201 34187 23259 34193
rect 23201 34184 23213 34187
rect 23164 34156 23213 34184
rect 23164 34144 23170 34156
rect 23201 34153 23213 34156
rect 23247 34153 23259 34187
rect 23201 34147 23259 34153
rect 29638 34144 29644 34196
rect 29696 34184 29702 34196
rect 29733 34187 29791 34193
rect 29733 34184 29745 34187
rect 29696 34156 29745 34184
rect 29696 34144 29702 34156
rect 29733 34153 29745 34156
rect 29779 34153 29791 34187
rect 29733 34147 29791 34153
rect 30466 34144 30472 34196
rect 30524 34184 30530 34196
rect 30561 34187 30619 34193
rect 30561 34184 30573 34187
rect 30524 34156 30573 34184
rect 30524 34144 30530 34156
rect 30561 34153 30573 34156
rect 30607 34153 30619 34187
rect 30561 34147 30619 34153
rect 31849 34187 31907 34193
rect 31849 34153 31861 34187
rect 31895 34184 31907 34187
rect 31938 34184 31944 34196
rect 31895 34156 31944 34184
rect 31895 34153 31907 34156
rect 31849 34147 31907 34153
rect 31938 34144 31944 34156
rect 31996 34144 32002 34196
rect 32861 34187 32919 34193
rect 32861 34153 32873 34187
rect 32907 34184 32919 34187
rect 33226 34184 33232 34196
rect 32907 34156 33232 34184
rect 32907 34153 32919 34156
rect 32861 34147 32919 34153
rect 33226 34144 33232 34156
rect 33284 34144 33290 34196
rect 16301 34119 16359 34125
rect 16301 34085 16313 34119
rect 16347 34116 16359 34119
rect 17126 34116 17132 34128
rect 16347 34088 17132 34116
rect 16347 34085 16359 34088
rect 16301 34079 16359 34085
rect 17126 34076 17132 34088
rect 17184 34076 17190 34128
rect 18693 34119 18751 34125
rect 18693 34085 18705 34119
rect 18739 34116 18751 34119
rect 20901 34119 20959 34125
rect 18739 34088 20760 34116
rect 18739 34085 18751 34088
rect 18693 34079 18751 34085
rect 4614 34048 4620 34060
rect 4575 34020 4620 34048
rect 4614 34008 4620 34020
rect 4672 34008 4678 34060
rect 6270 34048 6276 34060
rect 6231 34020 6276 34048
rect 6270 34008 6276 34020
rect 6328 34008 6334 34060
rect 7653 34051 7711 34057
rect 7653 34017 7665 34051
rect 7699 34048 7711 34051
rect 7926 34048 7932 34060
rect 7699 34020 7932 34048
rect 7699 34017 7711 34020
rect 7653 34011 7711 34017
rect 7926 34008 7932 34020
rect 7984 34008 7990 34060
rect 16206 34008 16212 34060
rect 16264 34048 16270 34060
rect 17405 34051 17463 34057
rect 17405 34048 17417 34051
rect 16264 34020 17417 34048
rect 16264 34008 16270 34020
rect 17405 34017 17417 34020
rect 17451 34017 17463 34051
rect 17405 34011 17463 34017
rect 17954 34008 17960 34060
rect 18012 34048 18018 34060
rect 18325 34051 18383 34057
rect 18325 34048 18337 34051
rect 18012 34020 18337 34048
rect 18012 34008 18018 34020
rect 18325 34017 18337 34020
rect 18371 34017 18383 34051
rect 18325 34011 18383 34017
rect 18782 34008 18788 34060
rect 18840 34048 18846 34060
rect 19337 34051 19395 34057
rect 19337 34048 19349 34051
rect 18840 34020 19349 34048
rect 18840 34008 18846 34020
rect 19337 34017 19349 34020
rect 19383 34017 19395 34051
rect 20732 34048 20760 34088
rect 20901 34085 20913 34119
rect 20947 34116 20959 34119
rect 22002 34116 22008 34128
rect 20947 34088 22008 34116
rect 20947 34085 20959 34088
rect 20901 34079 20959 34085
rect 22002 34076 22008 34088
rect 22060 34076 22066 34128
rect 20732 34020 22094 34048
rect 19337 34011 19395 34017
rect 1394 33980 1400 33992
rect 1355 33952 1400 33980
rect 1394 33940 1400 33952
rect 1452 33980 1458 33992
rect 2041 33983 2099 33989
rect 2041 33980 2053 33983
rect 1452 33952 2053 33980
rect 1452 33940 1458 33952
rect 2041 33949 2053 33952
rect 2087 33949 2099 33983
rect 7466 33980 7472 33992
rect 7427 33952 7472 33980
rect 2041 33943 2099 33949
rect 7466 33940 7472 33952
rect 7524 33940 7530 33992
rect 11333 33983 11391 33989
rect 11333 33949 11345 33983
rect 11379 33949 11391 33983
rect 12342 33980 12348 33992
rect 12303 33952 12348 33980
rect 11333 33943 11391 33949
rect 6086 33912 6092 33924
rect 6047 33884 6092 33912
rect 6086 33872 6092 33884
rect 6144 33872 6150 33924
rect 7745 33915 7803 33921
rect 7745 33881 7757 33915
rect 7791 33912 7803 33915
rect 8018 33912 8024 33924
rect 7791 33884 8024 33912
rect 7791 33881 7803 33884
rect 7745 33875 7803 33881
rect 8018 33872 8024 33884
rect 8076 33872 8082 33924
rect 1581 33847 1639 33853
rect 1581 33813 1593 33847
rect 1627 33844 1639 33847
rect 2682 33844 2688 33856
rect 1627 33816 2688 33844
rect 1627 33813 1639 33816
rect 1581 33807 1639 33813
rect 2682 33804 2688 33816
rect 2740 33804 2746 33856
rect 11146 33844 11152 33856
rect 11107 33816 11152 33844
rect 11146 33804 11152 33816
rect 11204 33804 11210 33856
rect 11348 33844 11376 33943
rect 12342 33940 12348 33952
rect 12400 33940 12406 33992
rect 12621 33983 12679 33989
rect 12621 33949 12633 33983
rect 12667 33980 12679 33983
rect 13265 33983 13323 33989
rect 13265 33980 13277 33983
rect 12667 33952 13277 33980
rect 12667 33949 12679 33952
rect 12621 33943 12679 33949
rect 13265 33949 13277 33952
rect 13311 33980 13323 33983
rect 15473 33983 15531 33989
rect 15473 33980 15485 33983
rect 13311 33952 15485 33980
rect 13311 33949 13323 33952
rect 13265 33943 13323 33949
rect 15473 33949 15485 33952
rect 15519 33980 15531 33983
rect 15654 33980 15660 33992
rect 15519 33952 15660 33980
rect 15519 33949 15531 33952
rect 15473 33943 15531 33949
rect 15654 33940 15660 33952
rect 15712 33980 15718 33992
rect 16117 33983 16175 33989
rect 16117 33980 16129 33983
rect 15712 33952 16129 33980
rect 15712 33940 15718 33952
rect 16117 33949 16129 33952
rect 16163 33949 16175 33983
rect 16117 33943 16175 33949
rect 17218 33940 17224 33992
rect 17276 33980 17282 33992
rect 17589 33983 17647 33989
rect 17589 33980 17601 33983
rect 17276 33952 17601 33980
rect 17276 33940 17282 33952
rect 17589 33949 17601 33952
rect 17635 33980 17647 33983
rect 18509 33983 18567 33989
rect 18509 33980 18521 33983
rect 17635 33952 18521 33980
rect 17635 33949 17647 33952
rect 17589 33943 17647 33949
rect 18509 33949 18521 33952
rect 18555 33980 18567 33983
rect 19521 33983 19579 33989
rect 19521 33980 19533 33983
rect 18555 33952 19533 33980
rect 18555 33949 18567 33952
rect 18509 33943 18567 33949
rect 19521 33949 19533 33952
rect 19567 33949 19579 33983
rect 20717 33983 20775 33989
rect 20717 33980 20729 33983
rect 19521 33943 19579 33949
rect 19628 33952 20729 33980
rect 12710 33872 12716 33924
rect 12768 33912 12774 33924
rect 17310 33912 17316 33924
rect 12768 33884 17316 33912
rect 12768 33872 12774 33884
rect 17310 33872 17316 33884
rect 17368 33912 17374 33924
rect 18233 33915 18291 33921
rect 18233 33912 18245 33915
rect 17368 33884 18245 33912
rect 17368 33872 17374 33884
rect 18233 33881 18245 33884
rect 18279 33881 18291 33915
rect 18233 33875 18291 33881
rect 19245 33915 19303 33921
rect 19245 33881 19257 33915
rect 19291 33912 19303 33915
rect 19334 33912 19340 33924
rect 19291 33884 19340 33912
rect 19291 33881 19303 33884
rect 19245 33875 19303 33881
rect 19334 33872 19340 33884
rect 19392 33872 19398 33924
rect 13262 33844 13268 33856
rect 11348 33816 13268 33844
rect 13262 33804 13268 33816
rect 13320 33844 13326 33856
rect 13538 33844 13544 33856
rect 13320 33816 13544 33844
rect 13320 33804 13326 33816
rect 13538 33804 13544 33816
rect 13596 33804 13602 33856
rect 16666 33804 16672 33856
rect 16724 33844 16730 33856
rect 16761 33847 16819 33853
rect 16761 33844 16773 33847
rect 16724 33816 16773 33844
rect 16724 33804 16730 33816
rect 16761 33813 16773 33816
rect 16807 33813 16819 33847
rect 16761 33807 16819 33813
rect 17773 33847 17831 33853
rect 17773 33813 17785 33847
rect 17819 33844 17831 33847
rect 19628 33844 19656 33952
rect 20717 33949 20729 33952
rect 20763 33949 20775 33983
rect 20717 33943 20775 33949
rect 22066 33912 22094 34020
rect 24486 34008 24492 34060
rect 24544 34048 24550 34060
rect 24857 34051 24915 34057
rect 24857 34048 24869 34051
rect 24544 34020 24869 34048
rect 24544 34008 24550 34020
rect 24857 34017 24869 34020
rect 24903 34017 24915 34051
rect 24857 34011 24915 34017
rect 26878 34008 26884 34060
rect 26936 34048 26942 34060
rect 27617 34051 27675 34057
rect 27617 34048 27629 34051
rect 26936 34020 27629 34048
rect 26936 34008 26942 34020
rect 27617 34017 27629 34020
rect 27663 34017 27675 34051
rect 27617 34011 27675 34017
rect 30101 34051 30159 34057
rect 30101 34017 30113 34051
rect 30147 34048 30159 34051
rect 30929 34051 30987 34057
rect 30929 34048 30941 34051
rect 30147 34020 30941 34048
rect 30147 34017 30159 34020
rect 30101 34011 30159 34017
rect 30929 34017 30941 34020
rect 30975 34048 30987 34051
rect 31481 34051 31539 34057
rect 31481 34048 31493 34051
rect 30975 34020 31493 34048
rect 30975 34017 30987 34020
rect 30929 34011 30987 34017
rect 31481 34017 31493 34020
rect 31527 34048 31539 34051
rect 31570 34048 31576 34060
rect 31527 34020 31576 34048
rect 31527 34017 31539 34020
rect 31481 34011 31539 34017
rect 31570 34008 31576 34020
rect 31628 34008 31634 34060
rect 24394 33940 24400 33992
rect 24452 33980 24458 33992
rect 24581 33983 24639 33989
rect 24581 33980 24593 33983
rect 24452 33952 24593 33980
rect 24452 33940 24458 33952
rect 24581 33949 24593 33952
rect 24627 33949 24639 33983
rect 26050 33980 26056 33992
rect 26011 33952 26056 33980
rect 24581 33943 24639 33949
rect 26050 33940 26056 33952
rect 26108 33940 26114 33992
rect 26329 33983 26387 33989
rect 26329 33949 26341 33983
rect 26375 33980 26387 33983
rect 27154 33980 27160 33992
rect 26375 33952 27160 33980
rect 26375 33949 26387 33952
rect 26329 33943 26387 33949
rect 27154 33940 27160 33952
rect 27212 33940 27218 33992
rect 27341 33983 27399 33989
rect 27341 33949 27353 33983
rect 27387 33949 27399 33983
rect 27341 33943 27399 33949
rect 25866 33912 25872 33924
rect 19720 33884 21036 33912
rect 22066 33884 25872 33912
rect 19720 33853 19748 33884
rect 17819 33816 19656 33844
rect 19705 33847 19763 33853
rect 17819 33813 17831 33816
rect 17773 33807 17831 33813
rect 19705 33813 19717 33847
rect 19751 33813 19763 33847
rect 21008 33844 21036 33884
rect 25866 33872 25872 33884
rect 25924 33872 25930 33924
rect 23474 33844 23480 33856
rect 21008 33816 23480 33844
rect 19705 33807 19763 33813
rect 23474 33804 23480 33816
rect 23532 33804 23538 33856
rect 23566 33804 23572 33856
rect 23624 33844 23630 33856
rect 27356 33844 27384 33943
rect 28994 33940 29000 33992
rect 29052 33980 29058 33992
rect 29917 33983 29975 33989
rect 29917 33980 29929 33983
rect 29052 33952 29929 33980
rect 29052 33940 29058 33952
rect 29917 33949 29929 33952
rect 29963 33949 29975 33983
rect 30742 33980 30748 33992
rect 30703 33952 30748 33980
rect 29917 33943 29975 33949
rect 30742 33940 30748 33952
rect 30800 33940 30806 33992
rect 31662 33980 31668 33992
rect 31623 33952 31668 33980
rect 31662 33940 31668 33952
rect 31720 33940 31726 33992
rect 32490 33940 32496 33992
rect 32548 33980 32554 33992
rect 32677 33983 32735 33989
rect 32677 33980 32689 33983
rect 32548 33952 32689 33980
rect 32548 33940 32554 33952
rect 32677 33949 32689 33952
rect 32723 33949 32735 33983
rect 32677 33943 32735 33949
rect 37461 33983 37519 33989
rect 37461 33949 37473 33983
rect 37507 33980 37519 33983
rect 38102 33980 38108 33992
rect 37507 33952 38108 33980
rect 37507 33949 37519 33952
rect 37461 33943 37519 33949
rect 38102 33940 38108 33952
rect 38160 33940 38166 33992
rect 23624 33816 27384 33844
rect 23624 33804 23630 33816
rect 37734 33804 37740 33856
rect 37792 33844 37798 33856
rect 37921 33847 37979 33853
rect 37921 33844 37933 33847
rect 37792 33816 37933 33844
rect 37792 33804 37798 33816
rect 37921 33813 37933 33816
rect 37967 33813 37979 33847
rect 37921 33807 37979 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 10413 33643 10471 33649
rect 10413 33609 10425 33643
rect 10459 33640 10471 33643
rect 11974 33640 11980 33652
rect 10459 33612 11980 33640
rect 10459 33609 10471 33612
rect 10413 33603 10471 33609
rect 4614 33572 4620 33584
rect 4575 33544 4620 33572
rect 4614 33532 4620 33544
rect 4672 33532 4678 33584
rect 8018 33572 8024 33584
rect 7931 33544 8024 33572
rect 8018 33532 8024 33544
rect 8076 33572 8082 33584
rect 10428 33572 10456 33603
rect 11974 33600 11980 33612
rect 12032 33600 12038 33652
rect 16117 33643 16175 33649
rect 16117 33609 16129 33643
rect 16163 33640 16175 33643
rect 16206 33640 16212 33652
rect 16163 33612 16212 33640
rect 16163 33609 16175 33612
rect 16117 33603 16175 33609
rect 16206 33600 16212 33612
rect 16264 33600 16270 33652
rect 19797 33643 19855 33649
rect 19797 33609 19809 33643
rect 19843 33640 19855 33643
rect 20162 33640 20168 33652
rect 19843 33612 20168 33640
rect 19843 33609 19855 33612
rect 19797 33603 19855 33609
rect 20162 33600 20168 33612
rect 20220 33600 20226 33652
rect 32490 33640 32496 33652
rect 32451 33612 32496 33640
rect 32490 33600 32496 33612
rect 32548 33600 32554 33652
rect 8076 33544 10456 33572
rect 18616 33544 19656 33572
rect 8076 33532 8082 33544
rect 7466 33464 7472 33516
rect 7524 33504 7530 33516
rect 7745 33507 7803 33513
rect 7745 33504 7757 33507
rect 7524 33476 7757 33504
rect 7524 33464 7530 33476
rect 7745 33473 7757 33476
rect 7791 33504 7803 33507
rect 10229 33507 10287 33513
rect 7791 33476 8248 33504
rect 7791 33473 7803 33476
rect 7745 33467 7803 33473
rect 2774 33396 2780 33448
rect 2832 33436 2838 33448
rect 2958 33436 2964 33448
rect 2832 33408 2877 33436
rect 2919 33408 2964 33436
rect 2832 33396 2838 33408
rect 2958 33396 2964 33408
rect 3016 33396 3022 33448
rect 7926 33436 7932 33448
rect 7887 33408 7932 33436
rect 7926 33396 7932 33408
rect 7984 33396 7990 33448
rect 8220 33436 8248 33476
rect 10229 33473 10241 33507
rect 10275 33504 10287 33507
rect 10502 33504 10508 33516
rect 10275 33476 10508 33504
rect 10275 33473 10287 33476
rect 10229 33467 10287 33473
rect 10502 33464 10508 33476
rect 10560 33464 10566 33516
rect 12437 33507 12495 33513
rect 12437 33473 12449 33507
rect 12483 33504 12495 33507
rect 12710 33504 12716 33516
rect 12483 33476 12716 33504
rect 12483 33473 12495 33476
rect 12437 33467 12495 33473
rect 12710 33464 12716 33476
rect 12768 33464 12774 33516
rect 16666 33504 16672 33516
rect 16627 33476 16672 33504
rect 16666 33464 16672 33476
rect 16724 33504 16730 33516
rect 16724 33476 17172 33504
rect 16724 33464 16730 33476
rect 11146 33436 11152 33448
rect 8220 33408 11152 33436
rect 11146 33396 11152 33408
rect 11204 33396 11210 33448
rect 12161 33439 12219 33445
rect 12161 33436 12173 33439
rect 11624 33408 12173 33436
rect 7742 33328 7748 33380
rect 7800 33368 7806 33380
rect 11054 33368 11060 33380
rect 7800 33340 11060 33368
rect 7800 33328 7806 33340
rect 7098 33300 7104 33312
rect 7059 33272 7104 33300
rect 7098 33260 7104 33272
rect 7156 33260 7162 33312
rect 7558 33300 7564 33312
rect 7519 33272 7564 33300
rect 7558 33260 7564 33272
rect 7616 33260 7622 33312
rect 8036 33309 8064 33340
rect 11054 33328 11060 33340
rect 11112 33328 11118 33380
rect 8021 33303 8079 33309
rect 8021 33269 8033 33303
rect 8067 33269 8079 33303
rect 8021 33263 8079 33269
rect 10502 33260 10508 33312
rect 10560 33300 10566 33312
rect 11624 33309 11652 33408
rect 12161 33405 12173 33408
rect 12207 33405 12219 33439
rect 16942 33436 16948 33448
rect 16903 33408 16948 33436
rect 12161 33399 12219 33405
rect 16942 33396 16948 33408
rect 17000 33396 17006 33448
rect 17144 33436 17172 33476
rect 17218 33464 17224 33516
rect 17276 33504 17282 33516
rect 18616 33513 18644 33544
rect 18601 33507 18659 33513
rect 18601 33504 18613 33507
rect 17276 33476 18613 33504
rect 17276 33464 17282 33476
rect 18601 33473 18613 33476
rect 18647 33473 18659 33507
rect 18601 33467 18659 33473
rect 18690 33464 18696 33516
rect 18748 33504 18754 33516
rect 18877 33507 18935 33513
rect 18748 33476 18793 33504
rect 18748 33464 18754 33476
rect 18877 33473 18889 33507
rect 18923 33504 18935 33507
rect 19334 33504 19340 33516
rect 18923 33476 19340 33504
rect 18923 33473 18935 33476
rect 18877 33467 18935 33473
rect 19334 33464 19340 33476
rect 19392 33504 19398 33516
rect 19628 33513 19656 33544
rect 19613 33507 19671 33513
rect 19392 33476 19564 33504
rect 19392 33464 19398 33476
rect 18138 33436 18144 33448
rect 17144 33408 18144 33436
rect 18138 33396 18144 33408
rect 18196 33396 18202 33448
rect 18708 33436 18736 33464
rect 19429 33439 19487 33445
rect 19429 33436 19441 33439
rect 18708 33408 19441 33436
rect 19429 33405 19441 33408
rect 19475 33405 19487 33439
rect 19536 33436 19564 33476
rect 19613 33473 19625 33507
rect 19659 33473 19671 33507
rect 32306 33504 32312 33516
rect 32267 33476 32312 33504
rect 19613 33467 19671 33473
rect 32306 33464 32312 33476
rect 32364 33464 32370 33516
rect 24486 33436 24492 33448
rect 19536 33408 20024 33436
rect 24447 33408 24492 33436
rect 19429 33399 19487 33405
rect 19996 33312 20024 33408
rect 24486 33396 24492 33408
rect 24544 33396 24550 33448
rect 24670 33436 24676 33448
rect 24631 33408 24676 33436
rect 24670 33396 24676 33408
rect 24728 33396 24734 33448
rect 25590 33436 25596 33448
rect 25551 33408 25596 33436
rect 25590 33396 25596 33408
rect 25648 33396 25654 33448
rect 31570 33396 31576 33448
rect 31628 33436 31634 33448
rect 32125 33439 32183 33445
rect 32125 33436 32137 33439
rect 31628 33408 32137 33436
rect 31628 33396 31634 33408
rect 32125 33405 32137 33408
rect 32171 33405 32183 33439
rect 32125 33399 32183 33405
rect 10873 33303 10931 33309
rect 10873 33300 10885 33303
rect 10560 33272 10885 33300
rect 10560 33260 10566 33272
rect 10873 33269 10885 33272
rect 10919 33300 10931 33303
rect 11609 33303 11667 33309
rect 11609 33300 11621 33303
rect 10919 33272 11621 33300
rect 10919 33269 10931 33272
rect 10873 33263 10931 33269
rect 11609 33269 11621 33272
rect 11655 33269 11667 33303
rect 18414 33300 18420 33312
rect 18375 33272 18420 33300
rect 11609 33263 11667 33269
rect 18414 33260 18420 33272
rect 18472 33260 18478 33312
rect 18598 33300 18604 33312
rect 18559 33272 18604 33300
rect 18598 33260 18604 33272
rect 18656 33300 18662 33312
rect 19337 33303 19395 33309
rect 19337 33300 19349 33303
rect 18656 33272 19349 33300
rect 18656 33260 18662 33272
rect 19337 33269 19349 33272
rect 19383 33269 19395 33303
rect 19337 33263 19395 33269
rect 19978 33260 19984 33312
rect 20036 33300 20042 33312
rect 20257 33303 20315 33309
rect 20257 33300 20269 33303
rect 20036 33272 20269 33300
rect 20036 33260 20042 33272
rect 20257 33269 20269 33272
rect 20303 33269 20315 33303
rect 27154 33300 27160 33312
rect 27115 33272 27160 33300
rect 20257 33263 20315 33269
rect 27154 33260 27160 33272
rect 27212 33260 27218 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 11054 33056 11060 33108
rect 11112 33096 11118 33108
rect 11885 33099 11943 33105
rect 11885 33096 11897 33099
rect 11112 33068 11897 33096
rect 11112 33056 11118 33068
rect 11885 33065 11897 33068
rect 11931 33096 11943 33099
rect 12342 33096 12348 33108
rect 11931 33068 12348 33096
rect 11931 33065 11943 33068
rect 11885 33059 11943 33065
rect 12342 33056 12348 33068
rect 12400 33056 12406 33108
rect 17218 33096 17224 33108
rect 17179 33068 17224 33096
rect 17218 33056 17224 33068
rect 17276 33056 17282 33108
rect 18325 33099 18383 33105
rect 18325 33065 18337 33099
rect 18371 33096 18383 33099
rect 18690 33096 18696 33108
rect 18371 33068 18696 33096
rect 18371 33065 18383 33068
rect 18325 33059 18383 33065
rect 18690 33056 18696 33068
rect 18748 33056 18754 33108
rect 24486 33056 24492 33108
rect 24544 33096 24550 33108
rect 24581 33099 24639 33105
rect 24581 33096 24593 33099
rect 24544 33068 24593 33096
rect 24544 33056 24550 33068
rect 24581 33065 24593 33068
rect 24627 33065 24639 33099
rect 24581 33059 24639 33065
rect 2958 32920 2964 32972
rect 3016 32960 3022 32972
rect 4065 32963 4123 32969
rect 4065 32960 4077 32963
rect 3016 32932 4077 32960
rect 3016 32920 3022 32932
rect 4065 32929 4077 32932
rect 4111 32929 4123 32963
rect 4065 32923 4123 32929
rect 11793 32963 11851 32969
rect 11793 32929 11805 32963
rect 11839 32960 11851 32963
rect 11882 32960 11888 32972
rect 11839 32932 11888 32960
rect 11839 32929 11851 32932
rect 11793 32923 11851 32929
rect 11882 32920 11888 32932
rect 11940 32920 11946 32972
rect 14550 32920 14556 32972
rect 14608 32960 14614 32972
rect 14921 32963 14979 32969
rect 14921 32960 14933 32963
rect 14608 32932 14933 32960
rect 14608 32920 14614 32932
rect 14921 32929 14933 32932
rect 14967 32960 14979 32963
rect 15381 32963 15439 32969
rect 15381 32960 15393 32963
rect 14967 32932 15393 32960
rect 14967 32929 14979 32932
rect 14921 32923 14979 32929
rect 15381 32929 15393 32932
rect 15427 32929 15439 32963
rect 15381 32923 15439 32929
rect 17954 32920 17960 32972
rect 18012 32960 18018 32972
rect 18322 32960 18328 32972
rect 18012 32932 18328 32960
rect 18012 32920 18018 32932
rect 18322 32920 18328 32932
rect 18380 32920 18386 32972
rect 22833 32963 22891 32969
rect 22833 32929 22845 32963
rect 22879 32960 22891 32963
rect 23290 32960 23296 32972
rect 22879 32932 23296 32960
rect 22879 32929 22891 32932
rect 22833 32923 22891 32929
rect 23290 32920 23296 32932
rect 23348 32920 23354 32972
rect 25590 32960 25596 32972
rect 25551 32932 25596 32960
rect 25590 32920 25596 32932
rect 25648 32920 25654 32972
rect 27154 32920 27160 32972
rect 27212 32960 27218 32972
rect 27433 32963 27491 32969
rect 27433 32960 27445 32963
rect 27212 32932 27445 32960
rect 27212 32920 27218 32932
rect 27433 32929 27445 32932
rect 27479 32929 27491 32963
rect 27433 32923 27491 32929
rect 3786 32892 3792 32904
rect 3747 32864 3792 32892
rect 3786 32852 3792 32864
rect 3844 32852 3850 32904
rect 7558 32852 7564 32904
rect 7616 32892 7622 32904
rect 7745 32895 7803 32901
rect 7745 32892 7757 32895
rect 7616 32864 7757 32892
rect 7616 32852 7622 32864
rect 7745 32861 7757 32864
rect 7791 32861 7803 32895
rect 7745 32855 7803 32861
rect 11146 32852 11152 32904
rect 11204 32892 11210 32904
rect 11609 32895 11667 32901
rect 11609 32892 11621 32895
rect 11204 32864 11621 32892
rect 11204 32852 11210 32864
rect 11609 32861 11621 32864
rect 11655 32861 11667 32895
rect 11609 32855 11667 32861
rect 12434 32852 12440 32904
rect 12492 32892 12498 32904
rect 14642 32892 14648 32904
rect 12492 32864 12537 32892
rect 14603 32864 14648 32892
rect 12492 32852 12498 32864
rect 14642 32852 14648 32864
rect 14700 32852 14706 32904
rect 15930 32852 15936 32904
rect 15988 32892 15994 32904
rect 17037 32895 17095 32901
rect 17037 32892 17049 32895
rect 15988 32864 17049 32892
rect 15988 32852 15994 32864
rect 17037 32861 17049 32864
rect 17083 32861 17095 32895
rect 18138 32892 18144 32904
rect 18099 32864 18144 32892
rect 17037 32855 17095 32861
rect 18138 32852 18144 32864
rect 18196 32892 18202 32904
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18196 32864 19257 32892
rect 18196 32852 18202 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 22554 32892 22560 32904
rect 22515 32864 22560 32892
rect 19245 32855 19303 32861
rect 22554 32852 22560 32864
rect 22612 32852 22618 32904
rect 11885 32827 11943 32833
rect 11885 32793 11897 32827
rect 11931 32824 11943 32827
rect 27246 32824 27252 32836
rect 11931 32796 12434 32824
rect 27207 32796 27252 32824
rect 11931 32793 11943 32796
rect 11885 32787 11943 32793
rect 7374 32716 7380 32768
rect 7432 32756 7438 32768
rect 7561 32759 7619 32765
rect 7561 32756 7573 32759
rect 7432 32728 7573 32756
rect 7432 32716 7438 32728
rect 7561 32725 7573 32728
rect 7607 32725 7619 32759
rect 7561 32719 7619 32725
rect 11425 32759 11483 32765
rect 11425 32725 11437 32759
rect 11471 32756 11483 32759
rect 11514 32756 11520 32768
rect 11471 32728 11520 32756
rect 11471 32725 11483 32728
rect 11425 32719 11483 32725
rect 11514 32716 11520 32728
rect 11572 32716 11578 32768
rect 12406 32756 12434 32796
rect 27246 32784 27252 32796
rect 27304 32784 27310 32836
rect 12894 32756 12900 32768
rect 12406 32728 12900 32756
rect 12894 32716 12900 32728
rect 12952 32756 12958 32768
rect 17034 32756 17040 32768
rect 12952 32728 17040 32756
rect 12952 32716 12958 32728
rect 17034 32716 17040 32728
rect 17092 32716 17098 32768
rect 19889 32759 19947 32765
rect 19889 32725 19901 32759
rect 19935 32756 19947 32759
rect 19978 32756 19984 32768
rect 19935 32728 19984 32756
rect 19935 32725 19947 32728
rect 19889 32719 19947 32725
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 25593 32555 25651 32561
rect 25593 32521 25605 32555
rect 25639 32552 25651 32555
rect 27246 32552 27252 32564
rect 25639 32524 27252 32552
rect 25639 32521 25651 32524
rect 25593 32515 25651 32521
rect 27246 32512 27252 32524
rect 27304 32512 27310 32564
rect 4709 32487 4767 32493
rect 4709 32453 4721 32487
rect 4755 32484 4767 32487
rect 5258 32484 5264 32496
rect 4755 32456 5264 32484
rect 4755 32453 4767 32456
rect 4709 32447 4767 32453
rect 5258 32444 5264 32456
rect 5316 32444 5322 32496
rect 7374 32484 7380 32496
rect 7335 32456 7380 32484
rect 7374 32444 7380 32456
rect 7432 32444 7438 32496
rect 12621 32487 12679 32493
rect 12621 32453 12633 32487
rect 12667 32484 12679 32487
rect 15194 32484 15200 32496
rect 12667 32456 15200 32484
rect 12667 32453 12679 32456
rect 12621 32447 12679 32453
rect 15194 32444 15200 32456
rect 15252 32444 15258 32496
rect 1394 32416 1400 32428
rect 1355 32388 1400 32416
rect 1394 32376 1400 32388
rect 1452 32416 1458 32428
rect 2041 32419 2099 32425
rect 2041 32416 2053 32419
rect 1452 32388 2053 32416
rect 1452 32376 1458 32388
rect 2041 32385 2053 32388
rect 2087 32385 2099 32419
rect 2041 32379 2099 32385
rect 7098 32376 7104 32428
rect 7156 32416 7162 32428
rect 7193 32419 7251 32425
rect 7193 32416 7205 32419
rect 7156 32388 7205 32416
rect 7156 32376 7162 32388
rect 7193 32385 7205 32388
rect 7239 32385 7251 32419
rect 14274 32416 14280 32428
rect 14235 32388 14280 32416
rect 7193 32379 7251 32385
rect 14274 32376 14280 32388
rect 14332 32376 14338 32428
rect 17957 32419 18015 32425
rect 17957 32385 17969 32419
rect 18003 32416 18015 32419
rect 18046 32416 18052 32428
rect 18003 32388 18052 32416
rect 18003 32385 18015 32388
rect 17957 32379 18015 32385
rect 18046 32376 18052 32388
rect 18104 32376 18110 32428
rect 18693 32419 18751 32425
rect 18693 32385 18705 32419
rect 18739 32416 18751 32419
rect 18782 32416 18788 32428
rect 18739 32388 18788 32416
rect 18739 32385 18751 32388
rect 18693 32379 18751 32385
rect 18782 32376 18788 32388
rect 18840 32376 18846 32428
rect 23661 32419 23719 32425
rect 23661 32385 23673 32419
rect 23707 32416 23719 32419
rect 24670 32416 24676 32428
rect 23707 32388 24676 32416
rect 23707 32385 23719 32388
rect 23661 32379 23719 32385
rect 24670 32376 24676 32388
rect 24728 32376 24734 32428
rect 25406 32416 25412 32428
rect 25367 32388 25412 32416
rect 25406 32376 25412 32388
rect 25464 32376 25470 32428
rect 2866 32348 2872 32360
rect 2827 32320 2872 32348
rect 2866 32308 2872 32320
rect 2924 32308 2930 32360
rect 3050 32348 3056 32360
rect 3011 32320 3056 32348
rect 3050 32308 3056 32320
rect 3108 32308 3114 32360
rect 9030 32348 9036 32360
rect 8991 32320 9036 32348
rect 9030 32308 9036 32320
rect 9088 32308 9094 32360
rect 12434 32308 12440 32360
rect 12492 32348 12498 32360
rect 18233 32351 18291 32357
rect 12492 32320 12537 32348
rect 12492 32308 12498 32320
rect 18233 32317 18245 32351
rect 18279 32348 18291 32351
rect 19334 32348 19340 32360
rect 18279 32320 19340 32348
rect 18279 32317 18291 32320
rect 18233 32311 18291 32317
rect 19334 32308 19340 32320
rect 19392 32308 19398 32360
rect 22094 32308 22100 32360
rect 22152 32348 22158 32360
rect 23385 32351 23443 32357
rect 23385 32348 23397 32351
rect 22152 32320 23397 32348
rect 22152 32308 22158 32320
rect 23385 32317 23397 32320
rect 23431 32317 23443 32351
rect 23385 32311 23443 32317
rect 1578 32212 1584 32224
rect 1539 32184 1584 32212
rect 1578 32172 1584 32184
rect 1636 32172 1642 32224
rect 5353 32215 5411 32221
rect 5353 32181 5365 32215
rect 5399 32212 5411 32215
rect 5810 32212 5816 32224
rect 5399 32184 5816 32212
rect 5399 32181 5411 32184
rect 5353 32175 5411 32181
rect 5810 32172 5816 32184
rect 5868 32172 5874 32224
rect 18874 32212 18880 32224
rect 18835 32184 18880 32212
rect 18874 32172 18880 32184
rect 18932 32172 18938 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 2866 32008 2872 32020
rect 2827 31980 2872 32008
rect 2866 31968 2872 31980
rect 2924 31968 2930 32020
rect 18509 32011 18567 32017
rect 18509 31977 18521 32011
rect 18555 32008 18567 32011
rect 18598 32008 18604 32020
rect 18555 31980 18604 32008
rect 18555 31977 18567 31980
rect 18509 31971 18567 31977
rect 18598 31968 18604 31980
rect 18656 31968 18662 32020
rect 24394 32008 24400 32020
rect 24355 31980 24400 32008
rect 24394 31968 24400 31980
rect 24452 31968 24458 32020
rect 24486 31968 24492 32020
rect 24544 32008 24550 32020
rect 24581 32011 24639 32017
rect 24581 32008 24593 32011
rect 24544 31980 24593 32008
rect 24544 31968 24550 31980
rect 24581 31977 24593 31980
rect 24627 31977 24639 32011
rect 24581 31971 24639 31977
rect 16390 31900 16396 31952
rect 16448 31940 16454 31952
rect 18230 31940 18236 31952
rect 16448 31912 18236 31940
rect 16448 31900 16454 31912
rect 18230 31900 18236 31912
rect 18288 31900 18294 31952
rect 37642 31940 37648 31952
rect 37603 31912 37648 31940
rect 37642 31900 37648 31912
rect 37700 31900 37706 31952
rect 4154 31832 4160 31884
rect 4212 31872 4218 31884
rect 5258 31872 5264 31884
rect 4212 31844 5264 31872
rect 4212 31832 4218 31844
rect 5258 31832 5264 31844
rect 5316 31832 5322 31884
rect 5810 31872 5816 31884
rect 5771 31844 5816 31872
rect 5810 31832 5816 31844
rect 5868 31832 5874 31884
rect 6086 31832 6092 31884
rect 6144 31872 6150 31884
rect 6917 31875 6975 31881
rect 6917 31872 6929 31875
rect 6144 31844 6929 31872
rect 6144 31832 6150 31844
rect 6917 31841 6929 31844
rect 6963 31841 6975 31875
rect 11514 31872 11520 31884
rect 11475 31844 11520 31872
rect 6917 31835 6975 31841
rect 11514 31832 11520 31844
rect 11572 31832 11578 31884
rect 16574 31872 16580 31884
rect 16535 31844 16580 31872
rect 16574 31832 16580 31844
rect 16632 31832 16638 31884
rect 29822 31832 29828 31884
rect 29880 31872 29886 31884
rect 30193 31875 30251 31881
rect 30193 31872 30205 31875
rect 29880 31844 30205 31872
rect 29880 31832 29886 31844
rect 30193 31841 30205 31844
rect 30239 31872 30251 31875
rect 32401 31875 32459 31881
rect 32401 31872 32413 31875
rect 30239 31844 32413 31872
rect 30239 31841 30251 31844
rect 30193 31835 30251 31841
rect 32401 31841 32413 31844
rect 32447 31872 32459 31875
rect 33594 31872 33600 31884
rect 32447 31844 33600 31872
rect 32447 31841 32459 31844
rect 32401 31835 32459 31841
rect 33594 31832 33600 31844
rect 33652 31832 33658 31884
rect 7193 31807 7251 31813
rect 7193 31773 7205 31807
rect 7239 31804 7251 31807
rect 9858 31804 9864 31816
rect 7239 31776 9864 31804
rect 7239 31773 7251 31776
rect 7193 31767 7251 31773
rect 9858 31764 9864 31776
rect 9916 31764 9922 31816
rect 11330 31764 11336 31816
rect 11388 31804 11394 31816
rect 11793 31807 11851 31813
rect 11793 31804 11805 31807
rect 11388 31776 11805 31804
rect 11388 31764 11394 31776
rect 11793 31773 11805 31776
rect 11839 31773 11851 31807
rect 11793 31767 11851 31773
rect 12434 31764 12440 31816
rect 12492 31804 12498 31816
rect 12805 31807 12863 31813
rect 12805 31804 12817 31807
rect 12492 31776 12817 31804
rect 12492 31764 12498 31776
rect 12805 31773 12817 31776
rect 12851 31773 12863 31807
rect 12805 31767 12863 31773
rect 13078 31764 13084 31816
rect 13136 31804 13142 31816
rect 14093 31807 14151 31813
rect 14093 31804 14105 31807
rect 13136 31776 14105 31804
rect 13136 31764 13142 31776
rect 14093 31773 14105 31776
rect 14139 31773 14151 31807
rect 14093 31767 14151 31773
rect 15657 31807 15715 31813
rect 15657 31773 15669 31807
rect 15703 31804 15715 31807
rect 16117 31807 16175 31813
rect 16117 31804 16129 31807
rect 15703 31776 16129 31804
rect 15703 31773 15715 31776
rect 15657 31767 15715 31773
rect 16117 31773 16129 31776
rect 16163 31773 16175 31807
rect 16117 31767 16175 31773
rect 18414 31764 18420 31816
rect 18472 31804 18478 31816
rect 18601 31807 18659 31813
rect 18601 31804 18613 31807
rect 18472 31776 18613 31804
rect 18472 31764 18478 31776
rect 18601 31773 18613 31776
rect 18647 31773 18659 31807
rect 18601 31767 18659 31773
rect 19429 31807 19487 31813
rect 19429 31773 19441 31807
rect 19475 31804 19487 31807
rect 20070 31804 20076 31816
rect 19475 31776 20076 31804
rect 19475 31773 19487 31776
rect 19429 31767 19487 31773
rect 20070 31764 20076 31776
rect 20128 31764 20134 31816
rect 24578 31804 24584 31816
rect 24539 31776 24584 31804
rect 24578 31764 24584 31776
rect 24636 31764 24642 31816
rect 24673 31807 24731 31813
rect 24673 31773 24685 31807
rect 24719 31773 24731 31807
rect 24673 31767 24731 31773
rect 5534 31696 5540 31748
rect 5592 31736 5598 31748
rect 5629 31739 5687 31745
rect 5629 31736 5641 31739
rect 5592 31708 5641 31736
rect 5592 31696 5598 31708
rect 5629 31705 5641 31708
rect 5675 31705 5687 31739
rect 5629 31699 5687 31705
rect 7926 31696 7932 31748
rect 7984 31736 7990 31748
rect 14734 31736 14740 31748
rect 7984 31708 14740 31736
rect 7984 31696 7990 31708
rect 14734 31696 14740 31708
rect 14792 31696 14798 31748
rect 16298 31736 16304 31748
rect 16259 31708 16304 31736
rect 16298 31696 16304 31708
rect 16356 31696 16362 31748
rect 24486 31696 24492 31748
rect 24544 31736 24550 31748
rect 24688 31736 24716 31767
rect 35250 31764 35256 31816
rect 35308 31804 35314 31816
rect 36265 31807 36323 31813
rect 36265 31804 36277 31807
rect 35308 31776 36277 31804
rect 35308 31764 35314 31776
rect 36265 31773 36277 31776
rect 36311 31773 36323 31807
rect 36265 31767 36323 31773
rect 24857 31739 24915 31745
rect 24857 31736 24869 31739
rect 24544 31708 24716 31736
rect 24780 31708 24869 31736
rect 24544 31696 24550 31708
rect 12986 31668 12992 31680
rect 12947 31640 12992 31668
rect 12986 31628 12992 31640
rect 13044 31628 13050 31680
rect 22830 31628 22836 31680
rect 22888 31668 22894 31680
rect 23753 31671 23811 31677
rect 23753 31668 23765 31671
rect 22888 31640 23765 31668
rect 22888 31628 22894 31640
rect 23753 31637 23765 31640
rect 23799 31668 23811 31671
rect 24780 31668 24808 31708
rect 24857 31705 24869 31708
rect 24903 31705 24915 31739
rect 29914 31736 29920 31748
rect 29875 31708 29920 31736
rect 24857 31699 24915 31705
rect 29914 31696 29920 31708
rect 29972 31696 29978 31748
rect 32125 31739 32183 31745
rect 32125 31705 32137 31739
rect 32171 31736 32183 31739
rect 33134 31736 33140 31748
rect 32171 31708 33140 31736
rect 32171 31705 32183 31708
rect 32125 31699 32183 31705
rect 33134 31696 33140 31708
rect 33192 31696 33198 31748
rect 33318 31736 33324 31748
rect 33231 31708 33324 31736
rect 33318 31696 33324 31708
rect 33376 31736 33382 31748
rect 34054 31736 34060 31748
rect 33376 31708 34060 31736
rect 33376 31696 33382 31708
rect 34054 31696 34060 31708
rect 34112 31736 34118 31748
rect 34330 31736 34336 31748
rect 34112 31708 34336 31736
rect 34112 31696 34118 31708
rect 34330 31696 34336 31708
rect 34388 31696 34394 31748
rect 36170 31696 36176 31748
rect 36228 31736 36234 31748
rect 36510 31739 36568 31745
rect 36510 31736 36522 31739
rect 36228 31708 36522 31736
rect 36228 31696 36234 31708
rect 36510 31705 36522 31708
rect 36556 31705 36568 31739
rect 36510 31699 36568 31705
rect 25409 31671 25467 31677
rect 25409 31668 25421 31671
rect 23799 31640 25421 31668
rect 23799 31637 23811 31640
rect 23753 31631 23811 31637
rect 25409 31637 25421 31640
rect 25455 31668 25467 31671
rect 25590 31668 25596 31680
rect 25455 31640 25596 31668
rect 25455 31637 25467 31640
rect 25409 31631 25467 31637
rect 25590 31628 25596 31640
rect 25648 31628 25654 31680
rect 29546 31668 29552 31680
rect 29507 31640 29552 31668
rect 29546 31628 29552 31640
rect 29604 31628 29610 31680
rect 30006 31628 30012 31680
rect 30064 31668 30070 31680
rect 30837 31671 30895 31677
rect 30064 31640 30109 31668
rect 30064 31628 30070 31640
rect 30837 31637 30849 31671
rect 30883 31668 30895 31671
rect 31386 31668 31392 31680
rect 30883 31640 31392 31668
rect 30883 31637 30895 31640
rect 30837 31631 30895 31637
rect 31386 31628 31392 31640
rect 31444 31628 31450 31680
rect 31754 31668 31760 31680
rect 31715 31640 31760 31668
rect 31754 31628 31760 31640
rect 31812 31628 31818 31680
rect 32214 31628 32220 31680
rect 32272 31668 32278 31680
rect 32272 31640 32317 31668
rect 32272 31628 32278 31640
rect 32398 31628 32404 31680
rect 32456 31668 32462 31680
rect 32953 31671 33011 31677
rect 32953 31668 32965 31671
rect 32456 31640 32965 31668
rect 32456 31628 32462 31640
rect 32953 31637 32965 31640
rect 32999 31637 33011 31671
rect 32953 31631 33011 31637
rect 33410 31628 33416 31680
rect 33468 31668 33474 31680
rect 33468 31640 33513 31668
rect 33468 31628 33474 31640
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 3050 31424 3056 31476
rect 3108 31464 3114 31476
rect 3697 31467 3755 31473
rect 3697 31464 3709 31467
rect 3108 31436 3709 31464
rect 3108 31424 3114 31436
rect 3697 31433 3709 31436
rect 3743 31433 3755 31467
rect 22281 31467 22339 31473
rect 3697 31427 3755 31433
rect 6886 31436 22232 31464
rect 1578 31356 1584 31408
rect 1636 31396 1642 31408
rect 2501 31399 2559 31405
rect 2501 31396 2513 31399
rect 1636 31368 2513 31396
rect 1636 31356 1642 31368
rect 2501 31365 2513 31368
rect 2547 31365 2559 31399
rect 2501 31359 2559 31365
rect 3602 31356 3608 31408
rect 3660 31396 3666 31408
rect 6886 31396 6914 31436
rect 3660 31368 6914 31396
rect 3660 31356 3666 31368
rect 9030 31356 9036 31408
rect 9088 31396 9094 31408
rect 9125 31399 9183 31405
rect 9125 31396 9137 31399
rect 9088 31368 9137 31396
rect 9088 31356 9094 31368
rect 9125 31365 9137 31368
rect 9171 31365 9183 31399
rect 9125 31359 9183 31365
rect 10965 31399 11023 31405
rect 10965 31365 10977 31399
rect 11011 31396 11023 31399
rect 11885 31399 11943 31405
rect 11885 31396 11897 31399
rect 11011 31368 11897 31396
rect 11011 31365 11023 31368
rect 10965 31359 11023 31365
rect 11885 31365 11897 31368
rect 11931 31396 11943 31399
rect 12066 31396 12072 31408
rect 11931 31368 12072 31396
rect 11931 31365 11943 31368
rect 11885 31359 11943 31365
rect 12066 31356 12072 31368
rect 12124 31396 12130 31408
rect 12986 31396 12992 31408
rect 12124 31368 12296 31396
rect 12947 31368 12992 31396
rect 12124 31356 12130 31368
rect 1394 31328 1400 31340
rect 1355 31300 1400 31328
rect 1394 31288 1400 31300
rect 1452 31288 1458 31340
rect 3878 31328 3884 31340
rect 3839 31300 3884 31328
rect 3878 31288 3884 31300
rect 3936 31288 3942 31340
rect 4525 31331 4583 31337
rect 4525 31297 4537 31331
rect 4571 31328 4583 31331
rect 4798 31328 4804 31340
rect 4571 31300 4804 31328
rect 4571 31297 4583 31300
rect 4525 31291 4583 31297
rect 4798 31288 4804 31300
rect 4856 31288 4862 31340
rect 5534 31328 5540 31340
rect 5495 31300 5540 31328
rect 5534 31288 5540 31300
rect 5592 31288 5598 31340
rect 12158 31328 12164 31340
rect 12119 31300 12164 31328
rect 12158 31288 12164 31300
rect 12216 31288 12222 31340
rect 2869 31263 2927 31269
rect 2869 31229 2881 31263
rect 2915 31229 2927 31263
rect 5810 31260 5816 31272
rect 5771 31232 5816 31260
rect 2869 31223 2927 31229
rect 1581 31195 1639 31201
rect 1581 31161 1593 31195
rect 1627 31192 1639 31195
rect 2884 31192 2912 31223
rect 5810 31220 5816 31232
rect 5868 31220 5874 31272
rect 6825 31263 6883 31269
rect 6825 31229 6837 31263
rect 6871 31260 6883 31263
rect 7285 31263 7343 31269
rect 7285 31260 7297 31263
rect 6871 31232 7297 31260
rect 6871 31229 6883 31232
rect 6825 31223 6883 31229
rect 7285 31229 7297 31232
rect 7331 31229 7343 31263
rect 7466 31260 7472 31272
rect 7427 31232 7472 31260
rect 7285 31223 7343 31229
rect 7466 31220 7472 31232
rect 7524 31220 7530 31272
rect 12069 31263 12127 31269
rect 12069 31229 12081 31263
rect 12115 31229 12127 31263
rect 12069 31223 12127 31229
rect 1627 31164 2912 31192
rect 1627 31161 1639 31164
rect 1581 31155 1639 31161
rect 4062 31152 4068 31204
rect 4120 31192 4126 31204
rect 8294 31192 8300 31204
rect 4120 31164 8300 31192
rect 4120 31152 4126 31164
rect 8294 31152 8300 31164
rect 8352 31192 8358 31204
rect 9030 31192 9036 31204
rect 8352 31164 9036 31192
rect 8352 31152 8358 31164
rect 9030 31152 9036 31164
rect 9088 31152 9094 31204
rect 12084 31192 12112 31223
rect 12158 31192 12164 31204
rect 12084 31164 12164 31192
rect 12158 31152 12164 31164
rect 12216 31152 12222 31204
rect 12268 31192 12296 31368
rect 12986 31356 12992 31368
rect 13044 31356 13050 31408
rect 14645 31399 14703 31405
rect 14645 31365 14657 31399
rect 14691 31396 14703 31399
rect 16574 31396 16580 31408
rect 14691 31368 16580 31396
rect 14691 31365 14703 31368
rect 14645 31359 14703 31365
rect 16574 31356 16580 31368
rect 16632 31356 16638 31408
rect 17034 31396 17040 31408
rect 16995 31368 17040 31396
rect 17034 31356 17040 31368
rect 17092 31356 17098 31408
rect 17954 31356 17960 31408
rect 18012 31396 18018 31408
rect 18049 31399 18107 31405
rect 18049 31396 18061 31399
rect 18012 31368 18061 31396
rect 18012 31356 18018 31368
rect 18049 31365 18061 31368
rect 18095 31365 18107 31399
rect 18049 31359 18107 31365
rect 18874 31356 18880 31408
rect 18932 31396 18938 31408
rect 19705 31399 19763 31405
rect 19705 31396 19717 31399
rect 18932 31368 19717 31396
rect 18932 31356 18938 31368
rect 19705 31365 19717 31368
rect 19751 31365 19763 31399
rect 22204 31396 22232 31436
rect 22281 31433 22293 31467
rect 22327 31464 22339 31467
rect 23566 31464 23572 31476
rect 22327 31436 23572 31464
rect 22327 31433 22339 31436
rect 22281 31427 22339 31433
rect 23566 31424 23572 31436
rect 23624 31424 23630 31476
rect 26050 31464 26056 31476
rect 26011 31436 26056 31464
rect 26050 31424 26056 31436
rect 26108 31424 26114 31476
rect 31573 31467 31631 31473
rect 31573 31433 31585 31467
rect 31619 31464 31631 31467
rect 31662 31464 31668 31476
rect 31619 31436 31668 31464
rect 31619 31433 31631 31436
rect 31573 31427 31631 31433
rect 31662 31424 31668 31436
rect 31720 31424 31726 31476
rect 32214 31424 32220 31476
rect 32272 31464 32278 31476
rect 32493 31467 32551 31473
rect 32493 31464 32505 31467
rect 32272 31436 32505 31464
rect 32272 31424 32278 31436
rect 32493 31433 32505 31436
rect 32539 31433 32551 31467
rect 32493 31427 32551 31433
rect 32861 31467 32919 31473
rect 32861 31433 32873 31467
rect 32907 31464 32919 31467
rect 33318 31464 33324 31476
rect 32907 31436 33324 31464
rect 32907 31433 32919 31436
rect 32861 31427 32919 31433
rect 33318 31424 33324 31436
rect 33376 31424 33382 31476
rect 34517 31467 34575 31473
rect 34517 31433 34529 31467
rect 34563 31433 34575 31467
rect 34517 31427 34575 31433
rect 23750 31396 23756 31408
rect 22204 31368 23756 31396
rect 19705 31359 19763 31365
rect 23750 31356 23756 31368
rect 23808 31356 23814 31408
rect 24486 31356 24492 31408
rect 24544 31396 24550 31408
rect 30561 31399 30619 31405
rect 24544 31368 25728 31396
rect 24544 31356 24550 31368
rect 17221 31331 17279 31337
rect 17221 31297 17233 31331
rect 17267 31297 17279 31331
rect 17221 31291 17279 31297
rect 19889 31331 19947 31337
rect 19889 31297 19901 31331
rect 19935 31328 19947 31331
rect 20070 31328 20076 31340
rect 19935 31300 20076 31328
rect 19935 31297 19947 31300
rect 19889 31291 19947 31297
rect 12805 31263 12863 31269
rect 12805 31229 12817 31263
rect 12851 31260 12863 31263
rect 13078 31260 13084 31272
rect 12851 31232 13084 31260
rect 12851 31229 12863 31232
rect 12805 31223 12863 31229
rect 13078 31220 13084 31232
rect 13136 31220 13142 31272
rect 17236 31260 17264 31291
rect 20070 31288 20076 31300
rect 20128 31288 20134 31340
rect 21542 31288 21548 31340
rect 21600 31328 21606 31340
rect 21821 31331 21879 31337
rect 21821 31328 21833 31331
rect 21600 31300 21833 31328
rect 21600 31288 21606 31300
rect 21821 31297 21833 31300
rect 21867 31297 21879 31331
rect 21821 31291 21879 31297
rect 22097 31331 22155 31337
rect 22097 31297 22109 31331
rect 22143 31328 22155 31331
rect 22186 31328 22192 31340
rect 22143 31300 22192 31328
rect 22143 31297 22155 31300
rect 22097 31291 22155 31297
rect 22186 31288 22192 31300
rect 22244 31288 22250 31340
rect 25590 31328 25596 31340
rect 25551 31300 25596 31328
rect 25590 31288 25596 31300
rect 25648 31288 25654 31340
rect 19334 31260 19340 31272
rect 17236 31232 19340 31260
rect 19334 31220 19340 31232
rect 19392 31220 19398 31272
rect 21910 31260 21916 31272
rect 21871 31232 21916 31260
rect 21910 31220 21916 31232
rect 21968 31220 21974 31272
rect 23290 31260 23296 31272
rect 23251 31232 23296 31260
rect 23290 31220 23296 31232
rect 23348 31220 23354 31272
rect 23477 31263 23535 31269
rect 23477 31229 23489 31263
rect 23523 31229 23535 31263
rect 23750 31260 23756 31272
rect 23711 31232 23756 31260
rect 23477 31223 23535 31229
rect 22830 31192 22836 31204
rect 12268 31164 22836 31192
rect 22830 31152 22836 31164
rect 22888 31152 22894 31204
rect 22922 31152 22928 31204
rect 22980 31192 22986 31204
rect 23492 31192 23520 31223
rect 23750 31220 23756 31232
rect 23808 31260 23814 31272
rect 25038 31260 25044 31272
rect 23808 31232 25044 31260
rect 23808 31220 23814 31232
rect 25038 31220 25044 31232
rect 25096 31220 25102 31272
rect 25700 31269 25728 31368
rect 30561 31365 30573 31399
rect 30607 31396 30619 31399
rect 31205 31399 31263 31405
rect 30607 31368 31156 31396
rect 30607 31365 30619 31368
rect 30561 31359 30619 31365
rect 25869 31331 25927 31337
rect 25869 31328 25881 31331
rect 25792 31300 25881 31328
rect 25685 31263 25743 31269
rect 25685 31229 25697 31263
rect 25731 31229 25743 31263
rect 25685 31223 25743 31229
rect 22980 31164 23520 31192
rect 22980 31152 22986 31164
rect 24578 31152 24584 31204
rect 24636 31192 24642 31204
rect 25792 31192 25820 31300
rect 25869 31297 25881 31300
rect 25915 31297 25927 31331
rect 25869 31291 25927 31297
rect 29549 31331 29607 31337
rect 29549 31297 29561 31331
rect 29595 31328 29607 31331
rect 30098 31328 30104 31340
rect 29595 31300 30104 31328
rect 29595 31297 29607 31300
rect 29549 31291 29607 31297
rect 30098 31288 30104 31300
rect 30156 31288 30162 31340
rect 31021 31331 31079 31337
rect 31021 31297 31033 31331
rect 31067 31297 31079 31331
rect 31128 31328 31156 31368
rect 31205 31365 31217 31399
rect 31251 31396 31263 31399
rect 31754 31396 31760 31408
rect 31251 31368 31760 31396
rect 31251 31365 31263 31368
rect 31205 31359 31263 31365
rect 31754 31356 31760 31368
rect 31812 31356 31818 31408
rect 34532 31396 34560 31427
rect 35498 31399 35556 31405
rect 35498 31396 35510 31399
rect 34532 31368 35510 31396
rect 35498 31365 35510 31368
rect 35544 31365 35556 31399
rect 35498 31359 35556 31365
rect 31294 31328 31300 31340
rect 31128 31300 31300 31328
rect 31021 31291 31079 31297
rect 29638 31260 29644 31272
rect 29599 31232 29644 31260
rect 29638 31220 29644 31232
rect 29696 31220 29702 31272
rect 29822 31260 29828 31272
rect 29783 31232 29828 31260
rect 29822 31220 29828 31232
rect 29880 31220 29886 31272
rect 31036 31260 31064 31291
rect 31294 31288 31300 31300
rect 31352 31288 31358 31340
rect 31386 31288 31392 31340
rect 31444 31328 31450 31340
rect 34330 31328 34336 31340
rect 31444 31300 31489 31328
rect 34291 31300 34336 31328
rect 31444 31288 31450 31300
rect 34330 31288 34336 31300
rect 34388 31288 34394 31340
rect 32490 31260 32496 31272
rect 31036 31232 32496 31260
rect 32490 31220 32496 31232
rect 32548 31220 32554 31272
rect 32953 31263 33011 31269
rect 32953 31229 32965 31263
rect 32999 31229 33011 31263
rect 33134 31260 33140 31272
rect 33095 31232 33140 31260
rect 32953 31223 33011 31229
rect 24636 31164 25820 31192
rect 24636 31152 24642 31164
rect 29914 31152 29920 31204
rect 29972 31192 29978 31204
rect 32968 31192 32996 31223
rect 33134 31220 33140 31232
rect 33192 31220 33198 31272
rect 34790 31220 34796 31272
rect 34848 31260 34854 31272
rect 35250 31260 35256 31272
rect 34848 31232 35256 31260
rect 34848 31220 34854 31232
rect 35250 31220 35256 31232
rect 35308 31220 35314 31272
rect 29972 31164 32996 31192
rect 29972 31152 29978 31164
rect 2682 31133 2688 31136
rect 2666 31127 2688 31133
rect 2666 31093 2678 31127
rect 2666 31087 2688 31093
rect 2682 31084 2688 31087
rect 2740 31084 2746 31136
rect 2774 31084 2780 31136
rect 2832 31124 2838 31136
rect 3145 31127 3203 31133
rect 2832 31096 2877 31124
rect 2832 31084 2838 31096
rect 3145 31093 3157 31127
rect 3191 31124 3203 31127
rect 3602 31124 3608 31136
rect 3191 31096 3608 31124
rect 3191 31093 3203 31096
rect 3145 31087 3203 31093
rect 3602 31084 3608 31096
rect 3660 31084 3666 31136
rect 3970 31084 3976 31136
rect 4028 31124 4034 31136
rect 4341 31127 4399 31133
rect 4341 31124 4353 31127
rect 4028 31096 4353 31124
rect 4028 31084 4034 31096
rect 4341 31093 4353 31096
rect 4387 31093 4399 31127
rect 11974 31124 11980 31136
rect 11935 31096 11980 31124
rect 4341 31087 4399 31093
rect 11974 31084 11980 31096
rect 12032 31084 12038 31136
rect 12345 31127 12403 31133
rect 12345 31093 12357 31127
rect 12391 31124 12403 31127
rect 15378 31124 15384 31136
rect 12391 31096 15384 31124
rect 12391 31093 12403 31096
rect 12345 31087 12403 31093
rect 15378 31084 15384 31096
rect 15436 31084 15442 31136
rect 21634 31084 21640 31136
rect 21692 31124 21698 31136
rect 21821 31127 21879 31133
rect 21821 31124 21833 31127
rect 21692 31096 21833 31124
rect 21692 31084 21698 31096
rect 21821 31093 21833 31096
rect 21867 31093 21879 31127
rect 21821 31087 21879 31093
rect 24394 31084 24400 31136
rect 24452 31124 24458 31136
rect 25593 31127 25651 31133
rect 25593 31124 25605 31127
rect 24452 31096 25605 31124
rect 24452 31084 24458 31096
rect 25593 31093 25605 31096
rect 25639 31093 25651 31127
rect 25593 31087 25651 31093
rect 28626 31084 28632 31136
rect 28684 31124 28690 31136
rect 29181 31127 29239 31133
rect 29181 31124 29193 31127
rect 28684 31096 29193 31124
rect 28684 31084 28690 31096
rect 29181 31093 29193 31096
rect 29227 31093 29239 31127
rect 29181 31087 29239 31093
rect 36538 31084 36544 31136
rect 36596 31124 36602 31136
rect 36633 31127 36691 31133
rect 36633 31124 36645 31127
rect 36596 31096 36645 31124
rect 36596 31084 36602 31096
rect 36633 31093 36645 31096
rect 36679 31093 36691 31127
rect 36633 31087 36691 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 7466 30920 7472 30932
rect 7427 30892 7472 30920
rect 7466 30880 7472 30892
rect 7524 30880 7530 30932
rect 8389 30923 8447 30929
rect 7852 30892 8064 30920
rect 1394 30852 1400 30864
rect 1355 30824 1400 30852
rect 1394 30812 1400 30824
rect 1452 30812 1458 30864
rect 5810 30812 5816 30864
rect 5868 30852 5874 30864
rect 7852 30852 7880 30892
rect 5868 30824 7880 30852
rect 7929 30855 7987 30861
rect 5868 30812 5874 30824
rect 7929 30821 7941 30855
rect 7975 30821 7987 30855
rect 8036 30852 8064 30892
rect 8389 30889 8401 30923
rect 8435 30920 8447 30923
rect 9401 30923 9459 30929
rect 9401 30920 9413 30923
rect 8435 30892 9413 30920
rect 8435 30889 8447 30892
rect 8389 30883 8447 30889
rect 9401 30889 9413 30892
rect 9447 30889 9459 30923
rect 9858 30920 9864 30932
rect 9819 30892 9864 30920
rect 9401 30883 9459 30889
rect 8941 30855 8999 30861
rect 8941 30852 8953 30855
rect 8036 30824 8953 30852
rect 7929 30815 7987 30821
rect 8941 30821 8953 30824
rect 8987 30821 8999 30855
rect 9416 30852 9444 30883
rect 9858 30880 9864 30892
rect 9916 30880 9922 30932
rect 10321 30923 10379 30929
rect 10321 30920 10333 30923
rect 9968 30892 10333 30920
rect 9968 30852 9996 30892
rect 10321 30889 10333 30892
rect 10367 30920 10379 30923
rect 15194 30920 15200 30932
rect 10367 30892 14596 30920
rect 15155 30892 15200 30920
rect 10367 30889 10379 30892
rect 10321 30883 10379 30889
rect 14568 30852 14596 30892
rect 15194 30880 15200 30892
rect 15252 30880 15258 30932
rect 19429 30923 19487 30929
rect 19429 30920 19441 30923
rect 17788 30892 19441 30920
rect 17788 30864 17816 30892
rect 19429 30889 19441 30892
rect 19475 30889 19487 30923
rect 19429 30883 19487 30889
rect 20901 30923 20959 30929
rect 20901 30889 20913 30923
rect 20947 30920 20959 30923
rect 21634 30920 21640 30932
rect 20947 30892 21640 30920
rect 20947 30889 20959 30892
rect 20901 30883 20959 30889
rect 21634 30880 21640 30892
rect 21692 30880 21698 30932
rect 22005 30923 22063 30929
rect 22005 30889 22017 30923
rect 22051 30920 22063 30923
rect 22094 30920 22100 30932
rect 22051 30892 22100 30920
rect 22051 30889 22063 30892
rect 22005 30883 22063 30889
rect 22094 30880 22100 30892
rect 22152 30880 22158 30932
rect 22922 30920 22928 30932
rect 22883 30892 22928 30920
rect 22922 30880 22928 30892
rect 22980 30880 22986 30932
rect 23290 30880 23296 30932
rect 23348 30920 23354 30932
rect 23385 30923 23443 30929
rect 23385 30920 23397 30923
rect 23348 30892 23397 30920
rect 23348 30880 23354 30892
rect 23385 30889 23397 30892
rect 23431 30889 23443 30923
rect 24394 30920 24400 30932
rect 24355 30892 24400 30920
rect 23385 30883 23443 30889
rect 24394 30880 24400 30892
rect 24452 30880 24458 30932
rect 24857 30923 24915 30929
rect 24857 30889 24869 30923
rect 24903 30920 24915 30923
rect 25406 30920 25412 30932
rect 24903 30892 25412 30920
rect 24903 30889 24915 30892
rect 24857 30883 24915 30889
rect 25406 30880 25412 30892
rect 25464 30880 25470 30932
rect 28994 30920 29000 30932
rect 28955 30892 29000 30920
rect 28994 30880 29000 30892
rect 29052 30880 29058 30932
rect 29549 30923 29607 30929
rect 29549 30889 29561 30923
rect 29595 30920 29607 30923
rect 29638 30920 29644 30932
rect 29595 30892 29644 30920
rect 29595 30889 29607 30892
rect 29549 30883 29607 30889
rect 29638 30880 29644 30892
rect 29696 30880 29702 30932
rect 30006 30880 30012 30932
rect 30064 30920 30070 30932
rect 30745 30923 30803 30929
rect 30745 30920 30757 30923
rect 30064 30892 30757 30920
rect 30064 30880 30070 30892
rect 30745 30889 30757 30892
rect 30791 30889 30803 30923
rect 30745 30883 30803 30889
rect 31941 30923 31999 30929
rect 31941 30889 31953 30923
rect 31987 30920 31999 30923
rect 32306 30920 32312 30932
rect 31987 30892 32312 30920
rect 31987 30889 31999 30892
rect 31941 30883 31999 30889
rect 32306 30880 32312 30892
rect 32364 30880 32370 30932
rect 33045 30923 33103 30929
rect 33045 30889 33057 30923
rect 33091 30920 33103 30923
rect 33410 30920 33416 30932
rect 33091 30892 33416 30920
rect 33091 30889 33103 30892
rect 33045 30883 33103 30889
rect 33410 30880 33416 30892
rect 33468 30880 33474 30932
rect 35621 30923 35679 30929
rect 35621 30889 35633 30923
rect 35667 30920 35679 30923
rect 36170 30920 36176 30932
rect 35667 30892 36176 30920
rect 35667 30889 35679 30892
rect 35621 30883 35679 30889
rect 36170 30880 36176 30892
rect 36228 30880 36234 30932
rect 17770 30852 17776 30864
rect 9416 30824 9996 30852
rect 10060 30824 12434 30852
rect 14568 30824 17776 30852
rect 8941 30815 8999 30821
rect 3970 30784 3976 30796
rect 3931 30756 3976 30784
rect 3970 30744 3976 30756
rect 4028 30744 4034 30796
rect 4062 30744 4068 30796
rect 4120 30784 4126 30796
rect 4249 30787 4307 30793
rect 4249 30784 4261 30787
rect 4120 30756 4261 30784
rect 4120 30744 4126 30756
rect 4249 30753 4261 30756
rect 4295 30753 4307 30787
rect 4249 30747 4307 30753
rect 3237 30719 3295 30725
rect 3237 30685 3249 30719
rect 3283 30716 3295 30719
rect 3789 30719 3847 30725
rect 3789 30716 3801 30719
rect 3283 30688 3801 30716
rect 3283 30685 3295 30688
rect 3237 30679 3295 30685
rect 3789 30685 3801 30688
rect 3835 30685 3847 30719
rect 3789 30679 3847 30685
rect 7285 30719 7343 30725
rect 7285 30685 7297 30719
rect 7331 30716 7343 30719
rect 7944 30716 7972 30815
rect 10060 30784 10088 30824
rect 8128 30756 10088 30784
rect 8128 30725 8156 30756
rect 9140 30725 9168 30756
rect 7331 30688 7972 30716
rect 8113 30719 8171 30725
rect 7331 30685 7343 30688
rect 7285 30679 7343 30685
rect 8113 30685 8125 30719
rect 8159 30685 8171 30719
rect 8113 30679 8171 30685
rect 8205 30719 8263 30725
rect 8205 30685 8217 30719
rect 8251 30685 8263 30719
rect 8205 30679 8263 30685
rect 9125 30719 9183 30725
rect 9125 30685 9137 30719
rect 9171 30685 9183 30719
rect 9125 30679 9183 30685
rect 9217 30719 9275 30725
rect 9217 30685 9229 30719
rect 9263 30716 9275 30719
rect 9306 30716 9312 30728
rect 9263 30688 9312 30716
rect 9263 30685 9275 30688
rect 9217 30679 9275 30685
rect 8220 30580 8248 30679
rect 9306 30676 9312 30688
rect 9364 30676 9370 30728
rect 10060 30725 10088 30756
rect 10229 30787 10287 30793
rect 10229 30753 10241 30787
rect 10275 30784 10287 30787
rect 11330 30784 11336 30796
rect 10275 30756 10456 30784
rect 11291 30756 11336 30784
rect 10275 30753 10287 30756
rect 10229 30747 10287 30753
rect 10052 30719 10110 30725
rect 10052 30685 10064 30719
rect 10098 30685 10110 30719
rect 10052 30679 10110 30685
rect 8389 30651 8447 30657
rect 8389 30617 8401 30651
rect 8435 30648 8447 30651
rect 9401 30651 9459 30657
rect 9401 30648 9413 30651
rect 8435 30620 9413 30648
rect 8435 30617 8447 30620
rect 8389 30611 8447 30617
rect 9401 30617 9413 30620
rect 9447 30648 9459 30651
rect 9490 30648 9496 30660
rect 9447 30620 9496 30648
rect 9447 30617 9459 30620
rect 9401 30611 9459 30617
rect 9490 30608 9496 30620
rect 9548 30648 9554 30660
rect 10321 30651 10379 30657
rect 10321 30648 10333 30651
rect 9548 30620 10333 30648
rect 9548 30608 9554 30620
rect 10321 30617 10333 30620
rect 10367 30617 10379 30651
rect 10321 30611 10379 30617
rect 9306 30580 9312 30592
rect 8220 30552 9312 30580
rect 9306 30540 9312 30552
rect 9364 30580 9370 30592
rect 10428 30580 10456 30756
rect 11330 30744 11336 30756
rect 11388 30744 11394 30796
rect 12406 30784 12434 30824
rect 17770 30812 17776 30824
rect 17828 30812 17834 30864
rect 19245 30855 19303 30861
rect 19245 30852 19257 30855
rect 17972 30824 19257 30852
rect 14734 30784 14740 30796
rect 12406 30756 14412 30784
rect 14695 30756 14740 30784
rect 11146 30716 11152 30728
rect 11107 30688 11152 30716
rect 11146 30676 11152 30688
rect 11204 30676 11210 30728
rect 14384 30716 14412 30756
rect 14734 30744 14740 30756
rect 14792 30784 14798 30796
rect 15102 30784 15108 30796
rect 14792 30756 15108 30784
rect 14792 30744 14798 30756
rect 15102 30744 15108 30756
rect 15160 30744 15166 30796
rect 16298 30744 16304 30796
rect 16356 30784 16362 30796
rect 17972 30793 18000 30824
rect 19245 30821 19257 30824
rect 19291 30821 19303 30855
rect 19245 30815 19303 30821
rect 21085 30855 21143 30861
rect 21085 30821 21097 30855
rect 21131 30852 21143 30855
rect 22554 30852 22560 30864
rect 21131 30824 22560 30852
rect 21131 30821 21143 30824
rect 21085 30815 21143 30821
rect 22554 30812 22560 30824
rect 22612 30812 22618 30864
rect 17681 30787 17739 30793
rect 17681 30784 17693 30787
rect 16356 30756 17693 30784
rect 16356 30744 16362 30756
rect 17681 30753 17693 30756
rect 17727 30753 17739 30787
rect 17681 30747 17739 30753
rect 17957 30787 18015 30793
rect 17957 30753 17969 30787
rect 18003 30753 18015 30787
rect 17957 30747 18015 30753
rect 18693 30787 18751 30793
rect 18693 30753 18705 30787
rect 18739 30784 18751 30787
rect 19978 30784 19984 30796
rect 18739 30756 19984 30784
rect 18739 30753 18751 30756
rect 18693 30747 18751 30753
rect 19978 30744 19984 30756
rect 20036 30744 20042 30796
rect 20717 30787 20775 30793
rect 20717 30753 20729 30787
rect 20763 30784 20775 30787
rect 21637 30787 21695 30793
rect 21637 30784 21649 30787
rect 20763 30756 21649 30784
rect 20763 30753 20775 30756
rect 20717 30747 20775 30753
rect 21637 30753 21649 30756
rect 21683 30784 21695 30787
rect 21910 30784 21916 30796
rect 21683 30756 21916 30784
rect 21683 30753 21695 30756
rect 21637 30747 21695 30753
rect 15378 30716 15384 30728
rect 14384 30688 15240 30716
rect 15339 30688 15384 30716
rect 12986 30648 12992 30660
rect 12947 30620 12992 30648
rect 12986 30608 12992 30620
rect 13044 30608 13050 30660
rect 14550 30648 14556 30660
rect 14511 30620 14556 30648
rect 14550 30608 14556 30620
rect 14608 30608 14614 30660
rect 15212 30648 15240 30688
rect 15378 30676 15384 30688
rect 15436 30676 15442 30728
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 18064 30688 19441 30716
rect 18064 30660 18092 30688
rect 19429 30685 19441 30688
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 19518 30676 19524 30728
rect 19576 30716 19582 30728
rect 20732 30716 20760 30747
rect 21910 30744 21916 30756
rect 21968 30744 21974 30796
rect 24486 30784 24492 30796
rect 24447 30756 24492 30784
rect 24486 30744 24492 30756
rect 24544 30744 24550 30796
rect 30193 30787 30251 30793
rect 30193 30753 30205 30787
rect 30239 30784 30251 30787
rect 30834 30784 30840 30796
rect 30239 30756 30840 30784
rect 30239 30753 30251 30756
rect 30193 30747 30251 30753
rect 30834 30744 30840 30756
rect 30892 30784 30898 30796
rect 31297 30787 31355 30793
rect 31297 30784 31309 30787
rect 30892 30756 31309 30784
rect 30892 30744 30898 30756
rect 31297 30753 31309 30756
rect 31343 30753 31355 30787
rect 31297 30747 31355 30753
rect 33134 30744 33140 30796
rect 33192 30784 33198 30796
rect 33689 30787 33747 30793
rect 33689 30784 33701 30787
rect 33192 30756 33701 30784
rect 33192 30744 33198 30756
rect 33689 30753 33701 30756
rect 33735 30784 33747 30787
rect 36722 30784 36728 30796
rect 33735 30756 36728 30784
rect 33735 30753 33747 30756
rect 33689 30747 33747 30753
rect 36722 30744 36728 30756
rect 36780 30744 36786 30796
rect 20898 30716 20904 30728
rect 19576 30688 20760 30716
rect 20859 30688 20904 30716
rect 19576 30676 19582 30688
rect 20898 30676 20904 30688
rect 20956 30716 20962 30728
rect 21821 30719 21879 30725
rect 21821 30716 21833 30719
rect 20956 30688 21833 30716
rect 20956 30676 20962 30688
rect 21821 30685 21833 30688
rect 21867 30716 21879 30719
rect 22186 30716 22192 30728
rect 21867 30688 22192 30716
rect 21867 30685 21879 30688
rect 21821 30679 21879 30685
rect 22186 30676 22192 30688
rect 22244 30676 22250 30728
rect 22738 30716 22744 30728
rect 22699 30688 22744 30716
rect 22738 30676 22744 30688
rect 22796 30676 22802 30728
rect 24210 30676 24216 30728
rect 24268 30716 24274 30728
rect 24578 30716 24584 30728
rect 24268 30688 24584 30716
rect 24268 30676 24274 30688
rect 24578 30676 24584 30688
rect 24636 30716 24642 30728
rect 24673 30719 24731 30725
rect 24673 30716 24685 30719
rect 24636 30688 24685 30716
rect 24636 30676 24642 30688
rect 24673 30685 24685 30688
rect 24719 30685 24731 30719
rect 28442 30716 28448 30728
rect 28403 30688 28448 30716
rect 24673 30679 24731 30685
rect 28442 30676 28448 30688
rect 28500 30676 28506 30728
rect 28626 30716 28632 30728
rect 28587 30688 28632 30716
rect 28626 30676 28632 30688
rect 28684 30676 28690 30728
rect 28810 30716 28816 30728
rect 28771 30688 28816 30716
rect 28810 30676 28816 30688
rect 28868 30676 28874 30728
rect 29914 30716 29920 30728
rect 29875 30688 29920 30716
rect 29914 30676 29920 30688
rect 29972 30676 29978 30728
rect 30098 30676 30104 30728
rect 30156 30716 30162 30728
rect 31205 30719 31263 30725
rect 31205 30716 31217 30719
rect 30156 30688 31217 30716
rect 30156 30676 30162 30688
rect 31205 30685 31217 30688
rect 31251 30685 31263 30719
rect 31205 30679 31263 30685
rect 31386 30676 31392 30728
rect 31444 30716 31450 30728
rect 32125 30719 32183 30725
rect 32125 30716 32137 30719
rect 31444 30688 32137 30716
rect 31444 30676 31450 30688
rect 32125 30685 32137 30688
rect 32171 30685 32183 30719
rect 32125 30679 32183 30685
rect 32309 30719 32367 30725
rect 32309 30685 32321 30719
rect 32355 30716 32367 30719
rect 32398 30716 32404 30728
rect 32355 30688 32404 30716
rect 32355 30685 32367 30688
rect 32309 30679 32367 30685
rect 32398 30676 32404 30688
rect 32456 30676 32462 30728
rect 32490 30676 32496 30728
rect 32548 30716 32554 30728
rect 33502 30716 33508 30728
rect 32548 30688 32593 30716
rect 33463 30688 33508 30716
rect 32548 30676 32554 30688
rect 33502 30676 33508 30688
rect 33560 30676 33566 30728
rect 35434 30716 35440 30728
rect 35395 30688 35440 30716
rect 35434 30676 35440 30688
rect 35492 30676 35498 30728
rect 18046 30648 18052 30660
rect 15212 30620 18052 30648
rect 18046 30608 18052 30620
rect 18104 30608 18110 30660
rect 18509 30651 18567 30657
rect 18509 30617 18521 30651
rect 18555 30617 18567 30651
rect 18509 30611 18567 30617
rect 9364 30552 10456 30580
rect 16669 30583 16727 30589
rect 9364 30540 9370 30552
rect 16669 30549 16681 30583
rect 16715 30580 16727 30583
rect 18524 30580 18552 30611
rect 19334 30608 19340 30660
rect 19392 30648 19398 30660
rect 19705 30651 19763 30657
rect 19705 30648 19717 30651
rect 19392 30620 19717 30648
rect 19392 30608 19398 30620
rect 19705 30617 19717 30620
rect 19751 30648 19763 30651
rect 20254 30648 20260 30660
rect 19751 30620 20260 30648
rect 19751 30617 19763 30620
rect 19705 30611 19763 30617
rect 20254 30608 20260 30620
rect 20312 30648 20318 30660
rect 20625 30651 20683 30657
rect 20625 30648 20637 30651
rect 20312 30620 20637 30648
rect 20312 30608 20318 30620
rect 20625 30617 20637 30620
rect 20671 30648 20683 30651
rect 21542 30648 21548 30660
rect 20671 30620 21548 30648
rect 20671 30617 20683 30620
rect 20625 30611 20683 30617
rect 21542 30608 21548 30620
rect 21600 30608 21606 30660
rect 22830 30608 22836 30660
rect 22888 30648 22894 30660
rect 24397 30651 24455 30657
rect 24397 30648 24409 30651
rect 22888 30620 24409 30648
rect 22888 30608 22894 30620
rect 24397 30617 24409 30620
rect 24443 30648 24455 30651
rect 25317 30651 25375 30657
rect 25317 30648 25329 30651
rect 24443 30620 25329 30648
rect 24443 30617 24455 30620
rect 24397 30611 24455 30617
rect 25317 30617 25329 30620
rect 25363 30617 25375 30651
rect 25317 30611 25375 30617
rect 28721 30651 28779 30657
rect 28721 30617 28733 30651
rect 28767 30617 28779 30651
rect 28721 30611 28779 30617
rect 19242 30580 19248 30592
rect 16715 30552 19248 30580
rect 16715 30549 16727 30552
rect 16669 30543 16727 30549
rect 19242 30540 19248 30552
rect 19300 30580 19306 30592
rect 20070 30580 20076 30592
rect 19300 30552 20076 30580
rect 19300 30540 19306 30552
rect 20070 30540 20076 30552
rect 20128 30540 20134 30592
rect 27982 30580 27988 30592
rect 27943 30552 27988 30580
rect 27982 30540 27988 30552
rect 28040 30580 28046 30592
rect 28736 30580 28764 30611
rect 31846 30608 31852 30660
rect 31904 30648 31910 30660
rect 32217 30651 32275 30657
rect 32217 30648 32229 30651
rect 31904 30620 32229 30648
rect 31904 30608 31910 30620
rect 32217 30617 32229 30620
rect 32263 30617 32275 30651
rect 33520 30648 33548 30676
rect 32217 30611 32275 30617
rect 32324 30620 33548 30648
rect 28040 30552 28764 30580
rect 28040 30540 28046 30552
rect 29638 30540 29644 30592
rect 29696 30580 29702 30592
rect 30009 30583 30067 30589
rect 30009 30580 30021 30583
rect 29696 30552 30021 30580
rect 29696 30540 29702 30552
rect 30009 30549 30021 30552
rect 30055 30549 30067 30583
rect 31110 30580 31116 30592
rect 31023 30552 31116 30580
rect 30009 30543 30067 30549
rect 31110 30540 31116 30552
rect 31168 30580 31174 30592
rect 32324 30580 32352 30620
rect 33410 30580 33416 30592
rect 31168 30552 32352 30580
rect 33371 30552 33416 30580
rect 31168 30540 31174 30552
rect 33410 30540 33416 30552
rect 33468 30540 33474 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 3878 30376 3884 30388
rect 3839 30348 3884 30376
rect 3878 30336 3884 30348
rect 3936 30336 3942 30388
rect 4798 30376 4804 30388
rect 4759 30348 4804 30376
rect 4798 30336 4804 30348
rect 4856 30336 4862 30388
rect 19978 30336 19984 30388
rect 20036 30376 20042 30388
rect 20530 30376 20536 30388
rect 20036 30348 20536 30376
rect 20036 30336 20042 30348
rect 20530 30336 20536 30348
rect 20588 30336 20594 30388
rect 28442 30336 28448 30388
rect 28500 30376 28506 30388
rect 32398 30376 32404 30388
rect 28500 30348 32404 30376
rect 28500 30336 28506 30348
rect 4341 30311 4399 30317
rect 4341 30277 4353 30311
rect 4387 30308 4399 30311
rect 4706 30308 4712 30320
rect 4387 30280 4712 30308
rect 4387 30277 4399 30280
rect 4341 30271 4399 30277
rect 4706 30268 4712 30280
rect 4764 30308 4770 30320
rect 5261 30311 5319 30317
rect 5261 30308 5273 30311
rect 4764 30280 5273 30308
rect 4764 30268 4770 30280
rect 5261 30277 5273 30280
rect 5307 30277 5319 30311
rect 5261 30271 5319 30277
rect 11977 30311 12035 30317
rect 11977 30277 11989 30311
rect 12023 30308 12035 30311
rect 12066 30308 12072 30320
rect 12023 30280 12072 30308
rect 12023 30277 12035 30280
rect 11977 30271 12035 30277
rect 12066 30268 12072 30280
rect 12124 30268 12130 30320
rect 13909 30311 13967 30317
rect 13909 30277 13921 30311
rect 13955 30308 13967 30311
rect 15654 30308 15660 30320
rect 13955 30280 15660 30308
rect 13955 30277 13967 30280
rect 13909 30271 13967 30277
rect 15654 30268 15660 30280
rect 15712 30268 15718 30320
rect 19245 30311 19303 30317
rect 19245 30277 19257 30311
rect 19291 30308 19303 30311
rect 19334 30308 19340 30320
rect 19291 30280 19340 30308
rect 19291 30277 19303 30280
rect 19245 30271 19303 30277
rect 19334 30268 19340 30280
rect 19392 30268 19398 30320
rect 4062 30240 4068 30252
rect 3975 30212 4068 30240
rect 4062 30200 4068 30212
rect 4120 30240 4126 30252
rect 4985 30243 5043 30249
rect 4120 30212 4292 30240
rect 4120 30200 4126 30212
rect 4157 30175 4215 30181
rect 4157 30141 4169 30175
rect 4203 30141 4215 30175
rect 4264 30172 4292 30212
rect 4985 30209 4997 30243
rect 5031 30209 5043 30243
rect 4985 30203 5043 30209
rect 10965 30243 11023 30249
rect 10965 30209 10977 30243
rect 11011 30240 11023 30243
rect 11146 30240 11152 30252
rect 11011 30212 11152 30240
rect 11011 30209 11023 30212
rect 10965 30203 11023 30209
rect 5000 30172 5028 30203
rect 11146 30200 11152 30212
rect 11204 30200 11210 30252
rect 12250 30240 12256 30252
rect 12163 30212 12256 30240
rect 12250 30200 12256 30212
rect 12308 30200 12314 30252
rect 12526 30200 12532 30252
rect 12584 30240 12590 30252
rect 13357 30243 13415 30249
rect 13357 30240 13369 30243
rect 12584 30212 13369 30240
rect 12584 30200 12590 30212
rect 13357 30209 13369 30212
rect 13403 30209 13415 30243
rect 14090 30240 14096 30252
rect 14051 30212 14096 30240
rect 13357 30203 13415 30209
rect 4264 30144 5028 30172
rect 4157 30135 4215 30141
rect 4172 30104 4200 30135
rect 4798 30104 4804 30116
rect 4172 30076 4804 30104
rect 4798 30064 4804 30076
rect 4856 30064 4862 30116
rect 5000 30104 5028 30144
rect 5074 30132 5080 30184
rect 5132 30172 5138 30184
rect 8205 30175 8263 30181
rect 5132 30144 5177 30172
rect 5132 30132 5138 30144
rect 8205 30141 8217 30175
rect 8251 30172 8263 30175
rect 8294 30172 8300 30184
rect 8251 30144 8300 30172
rect 8251 30141 8263 30144
rect 8205 30135 8263 30141
rect 8294 30132 8300 30144
rect 8352 30132 8358 30184
rect 9122 30172 9128 30184
rect 9083 30144 9128 30172
rect 9122 30132 9128 30144
rect 9180 30132 9186 30184
rect 9306 30172 9312 30184
rect 9267 30144 9312 30172
rect 9306 30132 9312 30144
rect 9364 30132 9370 30184
rect 12158 30172 12164 30184
rect 12119 30144 12164 30172
rect 12158 30132 12164 30144
rect 12216 30132 12222 30184
rect 12268 30104 12296 30200
rect 13372 30172 13400 30203
rect 14090 30200 14096 30212
rect 14148 30200 14154 30252
rect 18046 30240 18052 30252
rect 18007 30212 18052 30240
rect 18046 30200 18052 30212
rect 18104 30240 18110 30252
rect 18969 30243 19027 30249
rect 18969 30240 18981 30243
rect 18104 30212 18981 30240
rect 18104 30200 18110 30212
rect 18969 30209 18981 30212
rect 19015 30209 19027 30243
rect 20438 30240 20444 30252
rect 20399 30212 20444 30240
rect 18969 30203 19027 30209
rect 20438 30200 20444 30212
rect 20496 30200 20502 30252
rect 21818 30200 21824 30252
rect 21876 30240 21882 30252
rect 22005 30243 22063 30249
rect 22005 30240 22017 30243
rect 21876 30212 22017 30240
rect 21876 30200 21882 30212
rect 22005 30209 22017 30212
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 29089 30243 29147 30249
rect 29089 30209 29101 30243
rect 29135 30240 29147 30243
rect 29196 30240 29224 30348
rect 32398 30336 32404 30348
rect 32456 30336 32462 30388
rect 29273 30311 29331 30317
rect 29273 30277 29285 30311
rect 29319 30308 29331 30311
rect 29546 30308 29552 30320
rect 29319 30280 29552 30308
rect 29319 30277 29331 30280
rect 29273 30271 29331 30277
rect 29546 30268 29552 30280
rect 29604 30268 29610 30320
rect 32493 30311 32551 30317
rect 32493 30277 32505 30311
rect 32539 30308 32551 30311
rect 34330 30308 34336 30320
rect 32539 30280 34336 30308
rect 32539 30277 32551 30280
rect 32493 30271 32551 30277
rect 34330 30268 34336 30280
rect 34388 30268 34394 30320
rect 29135 30212 29224 30240
rect 29365 30243 29423 30249
rect 29135 30209 29147 30212
rect 29089 30203 29147 30209
rect 29365 30209 29377 30243
rect 29411 30209 29423 30243
rect 29365 30203 29423 30209
rect 29457 30243 29515 30249
rect 29457 30209 29469 30243
rect 29503 30240 29515 30243
rect 30282 30240 30288 30252
rect 29503 30212 30288 30240
rect 29503 30209 29515 30212
rect 29457 30203 29515 30209
rect 18325 30175 18383 30181
rect 18325 30172 18337 30175
rect 13372 30144 18337 30172
rect 18325 30141 18337 30144
rect 18371 30172 18383 30175
rect 19153 30175 19211 30181
rect 18371 30144 19104 30172
rect 18371 30141 18383 30144
rect 18325 30135 18383 30141
rect 5000 30076 12296 30104
rect 12434 30064 12440 30116
rect 12492 30104 12498 30116
rect 18782 30104 18788 30116
rect 12492 30076 12537 30104
rect 18743 30076 18788 30104
rect 12492 30064 12498 30076
rect 18782 30064 18788 30076
rect 18840 30064 18846 30116
rect 19076 30104 19104 30144
rect 19153 30141 19165 30175
rect 19199 30172 19211 30175
rect 19334 30172 19340 30184
rect 19199 30144 19340 30172
rect 19199 30141 19211 30144
rect 19153 30135 19211 30141
rect 19334 30132 19340 30144
rect 19392 30132 19398 30184
rect 22646 30172 22652 30184
rect 22607 30144 22652 30172
rect 22646 30132 22652 30144
rect 22704 30132 22710 30184
rect 22833 30175 22891 30181
rect 22833 30141 22845 30175
rect 22879 30141 22891 30175
rect 23658 30172 23664 30184
rect 23619 30144 23664 30172
rect 22833 30135 22891 30141
rect 20346 30104 20352 30116
rect 19076 30076 20352 30104
rect 20346 30064 20352 30076
rect 20404 30064 20410 30116
rect 20625 30107 20683 30113
rect 20625 30073 20637 30107
rect 20671 30104 20683 30107
rect 21634 30104 21640 30116
rect 20671 30076 21640 30104
rect 20671 30073 20683 30076
rect 20625 30067 20683 30073
rect 21634 30064 21640 30076
rect 21692 30064 21698 30116
rect 22189 30107 22247 30113
rect 22189 30073 22201 30107
rect 22235 30104 22247 30107
rect 22848 30104 22876 30135
rect 23658 30132 23664 30144
rect 23716 30132 23722 30184
rect 29380 30172 29408 30203
rect 28736 30144 29408 30172
rect 22235 30076 22876 30104
rect 22235 30073 22247 30076
rect 22189 30067 22247 30073
rect 28736 30048 28764 30144
rect 28810 30064 28816 30116
rect 28868 30104 28874 30116
rect 29472 30104 29500 30203
rect 30282 30200 30288 30212
rect 30340 30200 30346 30252
rect 30466 30200 30472 30252
rect 30524 30240 30530 30252
rect 32309 30243 32367 30249
rect 32309 30240 32321 30243
rect 30524 30212 32321 30240
rect 30524 30200 30530 30212
rect 32309 30209 32321 30212
rect 32355 30209 32367 30243
rect 32309 30203 32367 30209
rect 35342 30200 35348 30252
rect 35400 30240 35406 30252
rect 35509 30243 35567 30249
rect 35509 30240 35521 30243
rect 35400 30212 35521 30240
rect 35400 30200 35406 30212
rect 35509 30209 35521 30212
rect 35555 30209 35567 30243
rect 35509 30203 35567 30209
rect 30745 30175 30803 30181
rect 30745 30141 30757 30175
rect 30791 30172 30803 30175
rect 30926 30172 30932 30184
rect 30791 30144 30932 30172
rect 30791 30141 30803 30144
rect 30745 30135 30803 30141
rect 30926 30132 30932 30144
rect 30984 30132 30990 30184
rect 31021 30175 31079 30181
rect 31021 30141 31033 30175
rect 31067 30141 31079 30175
rect 31021 30135 31079 30141
rect 32125 30175 32183 30181
rect 32125 30141 32137 30175
rect 32171 30141 32183 30175
rect 32125 30135 32183 30141
rect 28868 30076 29500 30104
rect 28868 30064 28874 30076
rect 30374 30064 30380 30116
rect 30432 30104 30438 30116
rect 31036 30104 31064 30135
rect 31481 30107 31539 30113
rect 31481 30104 31493 30107
rect 30432 30076 31493 30104
rect 30432 30064 30438 30076
rect 31481 30073 31493 30076
rect 31527 30073 31539 30107
rect 31481 30067 31539 30073
rect 4341 30039 4399 30045
rect 4341 30005 4353 30039
rect 4387 30036 4399 30039
rect 4614 30036 4620 30048
rect 4387 30008 4620 30036
rect 4387 30005 4399 30008
rect 4341 29999 4399 30005
rect 4614 29996 4620 30008
rect 4672 30036 4678 30048
rect 5261 30039 5319 30045
rect 5261 30036 5273 30039
rect 4672 30008 5273 30036
rect 4672 29996 4678 30008
rect 5261 30005 5273 30008
rect 5307 30036 5319 30039
rect 11974 30036 11980 30048
rect 5307 30008 11980 30036
rect 5307 30005 5319 30008
rect 5261 29999 5319 30005
rect 11974 29996 11980 30008
rect 12032 29996 12038 30048
rect 13262 30036 13268 30048
rect 13223 30008 13268 30036
rect 13262 29996 13268 30008
rect 13320 29996 13326 30048
rect 13906 29996 13912 30048
rect 13964 30036 13970 30048
rect 14550 30036 14556 30048
rect 13964 30008 14556 30036
rect 13964 29996 13970 30008
rect 14550 29996 14556 30008
rect 14608 30036 14614 30048
rect 14829 30039 14887 30045
rect 14829 30036 14841 30039
rect 14608 30008 14841 30036
rect 14608 29996 14614 30008
rect 14829 30005 14841 30008
rect 14875 30005 14887 30039
rect 14829 29999 14887 30005
rect 17770 29996 17776 30048
rect 17828 30036 17834 30048
rect 18969 30039 19027 30045
rect 18969 30036 18981 30039
rect 17828 30008 18981 30036
rect 17828 29996 17834 30008
rect 18969 30005 18981 30008
rect 19015 30005 19027 30039
rect 18969 29999 19027 30005
rect 19797 30039 19855 30045
rect 19797 30005 19809 30039
rect 19843 30036 19855 30039
rect 20070 30036 20076 30048
rect 19843 30008 20076 30036
rect 19843 30005 19855 30008
rect 19797 29999 19855 30005
rect 20070 29996 20076 30008
rect 20128 29996 20134 30048
rect 28629 30039 28687 30045
rect 28629 30005 28641 30039
rect 28675 30036 28687 30039
rect 28718 30036 28724 30048
rect 28675 30008 28724 30036
rect 28675 30005 28687 30008
rect 28629 29999 28687 30005
rect 28718 29996 28724 30008
rect 28776 29996 28782 30048
rect 29641 30039 29699 30045
rect 29641 30005 29653 30039
rect 29687 30036 29699 30039
rect 30742 30036 30748 30048
rect 29687 30008 30748 30036
rect 29687 30005 29699 30008
rect 29641 29999 29699 30005
rect 30742 29996 30748 30008
rect 30800 29996 30806 30048
rect 30926 29996 30932 30048
rect 30984 30036 30990 30048
rect 31570 30036 31576 30048
rect 30984 30008 31576 30036
rect 30984 29996 30990 30008
rect 31570 29996 31576 30008
rect 31628 30036 31634 30048
rect 32140 30036 32168 30135
rect 34790 30132 34796 30184
rect 34848 30172 34854 30184
rect 35253 30175 35311 30181
rect 35253 30172 35265 30175
rect 34848 30144 35265 30172
rect 34848 30132 34854 30144
rect 35253 30141 35265 30144
rect 35299 30141 35311 30175
rect 35253 30135 35311 30141
rect 31628 30008 32168 30036
rect 31628 29996 31634 30008
rect 33410 29996 33416 30048
rect 33468 30036 33474 30048
rect 36633 30039 36691 30045
rect 36633 30036 36645 30039
rect 33468 30008 36645 30036
rect 33468 29996 33474 30008
rect 36633 30005 36645 30008
rect 36679 30036 36691 30039
rect 37826 30036 37832 30048
rect 36679 30008 37832 30036
rect 36679 30005 36691 30008
rect 36633 29999 36691 30005
rect 37826 29996 37832 30008
rect 37884 29996 37890 30048
rect 38102 30036 38108 30048
rect 38063 30008 38108 30036
rect 38102 29996 38108 30008
rect 38160 29996 38166 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1581 29835 1639 29841
rect 1581 29801 1593 29835
rect 1627 29832 1639 29835
rect 2774 29832 2780 29844
rect 1627 29804 2780 29832
rect 1627 29801 1639 29804
rect 1581 29795 1639 29801
rect 2774 29792 2780 29804
rect 2832 29792 2838 29844
rect 3786 29792 3792 29844
rect 3844 29832 3850 29844
rect 3881 29835 3939 29841
rect 3881 29832 3893 29835
rect 3844 29804 3893 29832
rect 3844 29792 3850 29804
rect 3881 29801 3893 29804
rect 3927 29801 3939 29835
rect 3881 29795 3939 29801
rect 4341 29835 4399 29841
rect 4341 29801 4353 29835
rect 4387 29832 4399 29835
rect 4614 29832 4620 29844
rect 4387 29804 4620 29832
rect 4387 29801 4399 29804
rect 4341 29795 4399 29801
rect 4614 29792 4620 29804
rect 4672 29792 4678 29844
rect 7653 29835 7711 29841
rect 7653 29801 7665 29835
rect 7699 29832 7711 29835
rect 9306 29832 9312 29844
rect 7699 29804 9312 29832
rect 7699 29801 7711 29804
rect 7653 29795 7711 29801
rect 9306 29792 9312 29804
rect 9364 29792 9370 29844
rect 9493 29835 9551 29841
rect 9493 29801 9505 29835
rect 9539 29832 9551 29835
rect 11793 29835 11851 29841
rect 11793 29832 11805 29835
rect 9539 29804 11805 29832
rect 9539 29801 9551 29804
rect 9493 29795 9551 29801
rect 11793 29801 11805 29804
rect 11839 29832 11851 29835
rect 12066 29832 12072 29844
rect 11839 29804 12072 29832
rect 11839 29801 11851 29804
rect 11793 29795 11851 29801
rect 12066 29792 12072 29804
rect 12124 29792 12130 29844
rect 21634 29832 21640 29844
rect 21547 29804 21640 29832
rect 21634 29792 21640 29804
rect 21692 29792 21698 29844
rect 21818 29832 21824 29844
rect 21779 29804 21824 29832
rect 21818 29792 21824 29804
rect 21876 29792 21882 29844
rect 22281 29835 22339 29841
rect 22281 29801 22293 29835
rect 22327 29801 22339 29835
rect 22738 29832 22744 29844
rect 22699 29804 22744 29832
rect 22281 29795 22339 29801
rect 12158 29724 12164 29776
rect 12216 29764 12222 29776
rect 18138 29764 18144 29776
rect 12216 29736 18144 29764
rect 12216 29724 12222 29736
rect 18138 29724 18144 29736
rect 18196 29724 18202 29776
rect 21652 29764 21680 29792
rect 22296 29764 22324 29795
rect 22738 29792 22744 29804
rect 22796 29792 22802 29844
rect 30653 29835 30711 29841
rect 30653 29801 30665 29835
rect 30699 29832 30711 29835
rect 34790 29832 34796 29844
rect 30699 29804 34796 29832
rect 30699 29801 30711 29804
rect 30653 29795 30711 29801
rect 34790 29792 34796 29804
rect 34848 29792 34854 29844
rect 35069 29835 35127 29841
rect 35069 29801 35081 29835
rect 35115 29832 35127 29835
rect 35342 29832 35348 29844
rect 35115 29804 35348 29832
rect 35115 29801 35127 29804
rect 35069 29795 35127 29801
rect 35342 29792 35348 29804
rect 35400 29792 35406 29844
rect 21652 29736 22324 29764
rect 22646 29724 22652 29776
rect 22704 29764 22710 29776
rect 23201 29767 23259 29773
rect 23201 29764 23213 29767
rect 22704 29736 23213 29764
rect 22704 29724 22710 29736
rect 23201 29733 23213 29736
rect 23247 29733 23259 29767
rect 23201 29727 23259 29733
rect 31386 29724 31392 29776
rect 31444 29764 31450 29776
rect 32309 29767 32367 29773
rect 32309 29764 32321 29767
rect 31444 29736 32321 29764
rect 31444 29724 31450 29736
rect 32309 29733 32321 29736
rect 32355 29733 32367 29767
rect 37182 29764 37188 29776
rect 32309 29727 32367 29733
rect 36740 29736 37188 29764
rect 36740 29708 36768 29736
rect 37182 29724 37188 29736
rect 37240 29764 37246 29776
rect 37240 29736 37964 29764
rect 37240 29724 37246 29736
rect 4249 29699 4307 29705
rect 4249 29665 4261 29699
rect 4295 29696 4307 29699
rect 4798 29696 4804 29708
rect 4295 29668 4804 29696
rect 4295 29665 4307 29668
rect 4249 29659 4307 29665
rect 4798 29656 4804 29668
rect 4856 29656 4862 29708
rect 11974 29656 11980 29708
rect 12032 29696 12038 29708
rect 12529 29699 12587 29705
rect 12529 29696 12541 29699
rect 12032 29668 12541 29696
rect 12032 29656 12038 29668
rect 12529 29665 12541 29668
rect 12575 29665 12587 29699
rect 15654 29696 15660 29708
rect 15615 29668 15660 29696
rect 12529 29659 12587 29665
rect 15654 29656 15660 29668
rect 15712 29656 15718 29708
rect 17770 29696 17776 29708
rect 17731 29668 17776 29696
rect 17770 29656 17776 29668
rect 17828 29656 17834 29708
rect 20346 29656 20352 29708
rect 20404 29696 20410 29708
rect 21542 29696 21548 29708
rect 20404 29668 20576 29696
rect 21503 29668 21548 29696
rect 20404 29656 20410 29668
rect 1394 29628 1400 29640
rect 1355 29600 1400 29628
rect 1394 29588 1400 29600
rect 1452 29628 1458 29640
rect 2041 29631 2099 29637
rect 2041 29628 2053 29631
rect 1452 29600 2053 29628
rect 1452 29588 1458 29600
rect 2041 29597 2053 29600
rect 2087 29597 2099 29631
rect 4062 29628 4068 29640
rect 4023 29600 4068 29628
rect 2041 29591 2099 29597
rect 4062 29588 4068 29600
rect 4120 29588 4126 29640
rect 4341 29631 4399 29637
rect 4341 29597 4353 29631
rect 4387 29628 4399 29631
rect 4706 29628 4712 29640
rect 4387 29600 4712 29628
rect 4387 29597 4399 29600
rect 4341 29591 4399 29597
rect 4706 29588 4712 29600
rect 4764 29588 4770 29640
rect 12253 29631 12311 29637
rect 12253 29597 12265 29631
rect 12299 29628 12311 29631
rect 12299 29600 12434 29628
rect 12299 29597 12311 29600
rect 12253 29591 12311 29597
rect 8110 29520 8116 29572
rect 8168 29560 8174 29572
rect 9401 29563 9459 29569
rect 9401 29560 9413 29563
rect 8168 29532 9413 29560
rect 8168 29520 8174 29532
rect 9401 29529 9413 29532
rect 9447 29529 9459 29563
rect 9401 29523 9459 29529
rect 12406 29492 12434 29600
rect 14090 29588 14096 29640
rect 14148 29588 14154 29640
rect 15838 29588 15844 29640
rect 15896 29628 15902 29640
rect 15933 29631 15991 29637
rect 15933 29628 15945 29631
rect 15896 29600 15945 29628
rect 15896 29588 15902 29600
rect 15933 29597 15945 29600
rect 15979 29597 15991 29631
rect 15933 29591 15991 29597
rect 18049 29631 18107 29637
rect 18049 29597 18061 29631
rect 18095 29628 18107 29631
rect 20438 29628 20444 29640
rect 18095 29600 20444 29628
rect 18095 29597 18107 29600
rect 18049 29591 18107 29597
rect 14108 29560 14136 29588
rect 18064 29560 18092 29591
rect 20438 29588 20444 29600
rect 20496 29588 20502 29640
rect 20548 29637 20576 29668
rect 21542 29656 21548 29668
rect 21600 29696 21606 29708
rect 22373 29699 22431 29705
rect 22373 29696 22385 29699
rect 21600 29668 22385 29696
rect 21600 29656 21606 29668
rect 22373 29665 22385 29668
rect 22419 29665 22431 29699
rect 22373 29659 22431 29665
rect 28537 29699 28595 29705
rect 28537 29665 28549 29699
rect 28583 29696 28595 29699
rect 28718 29696 28724 29708
rect 28583 29668 28724 29696
rect 28583 29665 28595 29668
rect 28537 29659 28595 29665
rect 28718 29656 28724 29668
rect 28776 29656 28782 29708
rect 28997 29699 29055 29705
rect 28997 29665 29009 29699
rect 29043 29696 29055 29699
rect 29914 29696 29920 29708
rect 29043 29668 29920 29696
rect 29043 29665 29055 29668
rect 28997 29659 29055 29665
rect 29914 29656 29920 29668
rect 29972 29656 29978 29708
rect 31846 29696 31852 29708
rect 31807 29668 31852 29696
rect 31846 29656 31852 29668
rect 31904 29656 31910 29708
rect 36722 29696 36728 29708
rect 36683 29668 36728 29696
rect 36722 29656 36728 29668
rect 36780 29656 36786 29708
rect 37826 29696 37832 29708
rect 37787 29668 37832 29696
rect 37826 29656 37832 29668
rect 37884 29656 37890 29708
rect 37936 29705 37964 29736
rect 37921 29699 37979 29705
rect 37921 29665 37933 29699
rect 37967 29665 37979 29699
rect 37921 29659 37979 29665
rect 20533 29631 20591 29637
rect 20533 29597 20545 29631
rect 20579 29597 20591 29631
rect 20898 29628 20904 29640
rect 20533 29591 20591 29597
rect 20732 29600 20904 29628
rect 14108 29532 18092 29560
rect 13998 29492 14004 29504
rect 12406 29464 14004 29492
rect 13998 29452 14004 29464
rect 14056 29492 14062 29504
rect 14093 29495 14151 29501
rect 14093 29492 14105 29495
rect 14056 29464 14105 29492
rect 14056 29452 14062 29464
rect 14093 29461 14105 29464
rect 14139 29461 14151 29495
rect 14093 29455 14151 29461
rect 15197 29495 15255 29501
rect 15197 29461 15209 29495
rect 15243 29492 15255 29495
rect 15286 29492 15292 29504
rect 15243 29464 15292 29492
rect 15243 29461 15255 29464
rect 15197 29455 15255 29461
rect 15286 29452 15292 29464
rect 15344 29452 15350 29504
rect 20732 29501 20760 29600
rect 20898 29588 20904 29600
rect 20956 29628 20962 29640
rect 21637 29631 21695 29637
rect 21637 29628 21649 29631
rect 20956 29600 21649 29628
rect 20956 29588 20962 29600
rect 21637 29597 21649 29600
rect 21683 29628 21695 29631
rect 22557 29631 22615 29637
rect 22557 29628 22569 29631
rect 21683 29600 22569 29628
rect 21683 29597 21695 29600
rect 21637 29591 21695 29597
rect 22557 29597 22569 29600
rect 22603 29597 22615 29631
rect 22557 29591 22615 29597
rect 34514 29588 34520 29640
rect 34572 29628 34578 29640
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 34572 29600 34897 29628
rect 34572 29588 34578 29600
rect 34885 29597 34897 29600
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 35894 29588 35900 29640
rect 35952 29628 35958 29640
rect 36538 29628 36544 29640
rect 35952 29600 36544 29628
rect 35952 29588 35958 29600
rect 36538 29588 36544 29600
rect 36596 29588 36602 29640
rect 36633 29631 36691 29637
rect 36633 29597 36645 29631
rect 36679 29628 36691 29631
rect 37734 29628 37740 29640
rect 36679 29600 37740 29628
rect 36679 29597 36691 29600
rect 36633 29591 36691 29597
rect 37734 29588 37740 29600
rect 37792 29588 37798 29640
rect 21358 29560 21364 29572
rect 21271 29532 21364 29560
rect 21358 29520 21364 29532
rect 21416 29560 21422 29572
rect 22281 29563 22339 29569
rect 22281 29560 22293 29563
rect 21416 29532 22293 29560
rect 21416 29520 21422 29532
rect 22281 29529 22293 29532
rect 22327 29529 22339 29563
rect 28810 29560 28816 29572
rect 28771 29532 28816 29560
rect 22281 29523 22339 29529
rect 28810 29520 28816 29532
rect 28868 29520 28874 29572
rect 30742 29560 30748 29572
rect 30703 29532 30748 29560
rect 30742 29520 30748 29532
rect 30800 29520 30806 29572
rect 20717 29495 20775 29501
rect 20717 29461 20729 29495
rect 20763 29461 20775 29495
rect 20717 29455 20775 29461
rect 28994 29452 29000 29504
rect 29052 29492 29058 29504
rect 29730 29492 29736 29504
rect 29052 29464 29736 29492
rect 29052 29452 29058 29464
rect 29730 29452 29736 29464
rect 29788 29452 29794 29504
rect 36170 29492 36176 29504
rect 36131 29464 36176 29492
rect 36170 29452 36176 29464
rect 36228 29452 36234 29504
rect 37366 29492 37372 29504
rect 37327 29464 37372 29492
rect 37366 29452 37372 29464
rect 37424 29452 37430 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 9122 29248 9128 29300
rect 9180 29288 9186 29300
rect 17129 29291 17187 29297
rect 17129 29288 17141 29291
rect 9180 29260 17141 29288
rect 9180 29248 9186 29260
rect 17129 29257 17141 29260
rect 17175 29257 17187 29291
rect 18138 29288 18144 29300
rect 18099 29260 18144 29288
rect 17129 29251 17187 29257
rect 18138 29248 18144 29260
rect 18196 29248 18202 29300
rect 20254 29288 20260 29300
rect 20215 29260 20260 29288
rect 20254 29248 20260 29260
rect 20312 29248 20318 29300
rect 30466 29288 30472 29300
rect 29656 29260 30328 29288
rect 30427 29260 30472 29288
rect 13262 29180 13268 29232
rect 13320 29220 13326 29232
rect 18156 29220 18184 29248
rect 24486 29220 24492 29232
rect 13320 29192 15792 29220
rect 18156 29192 24492 29220
rect 13320 29180 13326 29192
rect 15013 29155 15071 29161
rect 15013 29121 15025 29155
rect 15059 29121 15071 29155
rect 15013 29115 15071 29121
rect 3053 29087 3111 29093
rect 3053 29053 3065 29087
rect 3099 29084 3111 29087
rect 3513 29087 3571 29093
rect 3513 29084 3525 29087
rect 3099 29056 3525 29084
rect 3099 29053 3111 29056
rect 3053 29047 3111 29053
rect 3513 29053 3525 29056
rect 3559 29053 3571 29087
rect 3694 29084 3700 29096
rect 3655 29056 3700 29084
rect 3513 29047 3571 29053
rect 3694 29044 3700 29056
rect 3752 29044 3758 29096
rect 3878 29044 3884 29096
rect 3936 29084 3942 29096
rect 4157 29087 4215 29093
rect 4157 29084 4169 29087
rect 3936 29056 4169 29084
rect 3936 29044 3942 29056
rect 4157 29053 4169 29056
rect 4203 29084 4215 29087
rect 9766 29084 9772 29096
rect 4203 29056 9772 29084
rect 4203 29053 4215 29056
rect 4157 29047 4215 29053
rect 9766 29044 9772 29056
rect 9824 29044 9830 29096
rect 12986 29084 12992 29096
rect 12947 29056 12992 29084
rect 12986 29044 12992 29056
rect 13044 29044 13050 29096
rect 13814 29084 13820 29096
rect 13775 29056 13820 29084
rect 13814 29044 13820 29056
rect 13872 29044 13878 29096
rect 14001 29087 14059 29093
rect 14001 29053 14013 29087
rect 14047 29053 14059 29087
rect 15028 29084 15056 29115
rect 15102 29112 15108 29164
rect 15160 29152 15166 29164
rect 15160 29124 15205 29152
rect 15160 29112 15166 29124
rect 15286 29112 15292 29164
rect 15344 29152 15350 29164
rect 15764 29161 15792 29192
rect 24486 29180 24492 29192
rect 24544 29180 24550 29232
rect 15749 29155 15807 29161
rect 15344 29124 15389 29152
rect 15344 29112 15350 29124
rect 15749 29121 15761 29155
rect 15795 29121 15807 29155
rect 17218 29152 17224 29164
rect 17179 29124 17224 29152
rect 15749 29115 15807 29121
rect 17218 29112 17224 29124
rect 17276 29112 17282 29164
rect 18233 29155 18291 29161
rect 18233 29121 18245 29155
rect 18279 29152 18291 29155
rect 19061 29155 19119 29161
rect 18279 29124 19012 29152
rect 18279 29121 18291 29124
rect 18233 29115 18291 29121
rect 15304 29084 15332 29112
rect 16666 29084 16672 29096
rect 15028 29056 15148 29084
rect 15304 29056 16672 29084
rect 14001 29047 14059 29053
rect 11701 29019 11759 29025
rect 11701 28985 11713 29019
rect 11747 29016 11759 29019
rect 14016 29016 14044 29047
rect 11747 28988 14044 29016
rect 15120 29016 15148 29056
rect 16666 29044 16672 29056
rect 16724 29044 16730 29096
rect 18785 29087 18843 29093
rect 18785 29053 18797 29087
rect 18831 29084 18843 29087
rect 18874 29084 18880 29096
rect 18831 29056 18880 29084
rect 18831 29053 18843 29056
rect 18785 29047 18843 29053
rect 18874 29044 18880 29056
rect 18932 29044 18938 29096
rect 18984 29084 19012 29124
rect 19061 29121 19073 29155
rect 19107 29152 19119 29155
rect 19334 29152 19340 29164
rect 19107 29124 19340 29152
rect 19107 29121 19119 29124
rect 19061 29115 19119 29121
rect 19334 29112 19340 29124
rect 19392 29112 19398 29164
rect 20073 29155 20131 29161
rect 20073 29121 20085 29155
rect 20119 29152 20131 29155
rect 20714 29152 20720 29164
rect 20119 29124 20720 29152
rect 20119 29121 20131 29124
rect 20073 29115 20131 29121
rect 20714 29112 20720 29124
rect 20772 29112 20778 29164
rect 23477 29155 23535 29161
rect 23477 29152 23489 29155
rect 23308 29124 23489 29152
rect 19426 29084 19432 29096
rect 18984 29056 19432 29084
rect 19426 29044 19432 29056
rect 19484 29044 19490 29096
rect 23308 29028 23336 29124
rect 23477 29121 23489 29124
rect 23523 29121 23535 29155
rect 24118 29152 24124 29164
rect 24079 29124 24124 29152
rect 23477 29115 23535 29121
rect 24118 29112 24124 29124
rect 24176 29112 24182 29164
rect 28813 29087 28871 29093
rect 28813 29053 28825 29087
rect 28859 29053 28871 29087
rect 28813 29047 28871 29053
rect 15930 29016 15936 29028
rect 15120 28988 15936 29016
rect 11747 28985 11759 28988
rect 11701 28979 11759 28985
rect 15930 28976 15936 28988
rect 15988 28976 15994 29028
rect 23017 29019 23075 29025
rect 23017 28985 23029 29019
rect 23063 29016 23075 29019
rect 23290 29016 23296 29028
rect 23063 28988 23296 29016
rect 23063 28985 23075 28988
rect 23017 28979 23075 28985
rect 23290 28976 23296 28988
rect 23348 28976 23354 29028
rect 24302 29016 24308 29028
rect 24263 28988 24308 29016
rect 24302 28976 24308 28988
rect 24360 28976 24366 29028
rect 28828 29016 28856 29047
rect 28902 29044 28908 29096
rect 28960 29084 28966 29096
rect 29089 29087 29147 29093
rect 29089 29084 29101 29087
rect 28960 29056 29101 29084
rect 28960 29044 28966 29056
rect 29089 29053 29101 29056
rect 29135 29053 29147 29087
rect 29089 29047 29147 29053
rect 29273 29087 29331 29093
rect 29273 29053 29285 29087
rect 29319 29084 29331 29087
rect 29656 29084 29684 29260
rect 29730 29180 29736 29232
rect 29788 29220 29794 29232
rect 30193 29223 30251 29229
rect 30193 29220 30205 29223
rect 29788 29192 30205 29220
rect 29788 29180 29794 29192
rect 30193 29189 30205 29192
rect 30239 29189 30251 29223
rect 30300 29220 30328 29260
rect 30466 29248 30472 29260
rect 30524 29248 30530 29300
rect 31110 29220 31116 29232
rect 30300 29192 31116 29220
rect 30193 29183 30251 29189
rect 31110 29180 31116 29192
rect 31168 29180 31174 29232
rect 31297 29223 31355 29229
rect 31297 29189 31309 29223
rect 31343 29220 31355 29223
rect 31386 29220 31392 29232
rect 31343 29192 31392 29220
rect 31343 29189 31355 29192
rect 31297 29183 31355 29189
rect 31386 29180 31392 29192
rect 31444 29180 31450 29232
rect 29917 29155 29975 29161
rect 29917 29121 29929 29155
rect 29963 29121 29975 29155
rect 30098 29152 30104 29164
rect 30059 29124 30104 29152
rect 29917 29115 29975 29121
rect 29319 29056 29684 29084
rect 29932 29084 29960 29115
rect 30098 29112 30104 29124
rect 30156 29112 30162 29164
rect 30282 29112 30288 29164
rect 30340 29152 30346 29164
rect 30340 29124 31524 29152
rect 30340 29112 30346 29124
rect 29932 29056 31432 29084
rect 29319 29053 29331 29056
rect 29273 29047 29331 29053
rect 31294 29016 31300 29028
rect 28828 28988 31300 29016
rect 31294 28976 31300 28988
rect 31352 28976 31358 29028
rect 8662 28948 8668 28960
rect 8623 28920 8668 28948
rect 8662 28908 8668 28920
rect 8720 28908 8726 28960
rect 9122 28908 9128 28960
rect 9180 28948 9186 28960
rect 9217 28951 9275 28957
rect 9217 28948 9229 28951
rect 9180 28920 9229 28948
rect 9180 28908 9186 28920
rect 9217 28917 9229 28920
rect 9263 28917 9275 28951
rect 14826 28948 14832 28960
rect 14787 28920 14832 28948
rect 9217 28911 9275 28917
rect 14826 28908 14832 28920
rect 14884 28908 14890 28960
rect 15289 28951 15347 28957
rect 15289 28917 15301 28951
rect 15335 28948 15347 28951
rect 15838 28948 15844 28960
rect 15335 28920 15844 28948
rect 15335 28917 15347 28920
rect 15289 28911 15347 28917
rect 15838 28908 15844 28920
rect 15896 28908 15902 28960
rect 20714 28948 20720 28960
rect 20675 28920 20720 28948
rect 20714 28908 20720 28920
rect 20772 28908 20778 28960
rect 23661 28951 23719 28957
rect 23661 28917 23673 28951
rect 23707 28948 23719 28951
rect 24210 28948 24216 28960
rect 23707 28920 24216 28948
rect 23707 28917 23719 28920
rect 23661 28911 23719 28917
rect 24210 28908 24216 28920
rect 24268 28908 24274 28960
rect 31404 28948 31432 29056
rect 31496 29025 31524 29124
rect 31481 29019 31539 29025
rect 31481 28985 31493 29019
rect 31527 29016 31539 29019
rect 32030 29016 32036 29028
rect 31527 28988 32036 29016
rect 31527 28985 31539 28988
rect 31481 28979 31539 28985
rect 32030 28976 32036 28988
rect 32088 28976 32094 29028
rect 32490 28948 32496 28960
rect 31404 28920 32496 28948
rect 32490 28908 32496 28920
rect 32548 28908 32554 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 3237 28747 3295 28753
rect 3237 28713 3249 28747
rect 3283 28744 3295 28747
rect 3694 28744 3700 28756
rect 3283 28716 3700 28744
rect 3283 28713 3295 28716
rect 3237 28707 3295 28713
rect 3694 28704 3700 28716
rect 3752 28704 3758 28756
rect 4433 28747 4491 28753
rect 4433 28713 4445 28747
rect 4479 28744 4491 28747
rect 4614 28744 4620 28756
rect 4479 28716 4620 28744
rect 4479 28713 4491 28716
rect 4433 28707 4491 28713
rect 4614 28704 4620 28716
rect 4672 28704 4678 28756
rect 15838 28744 15844 28756
rect 15799 28716 15844 28744
rect 15838 28704 15844 28716
rect 15896 28704 15902 28756
rect 24394 28744 24400 28756
rect 24355 28716 24400 28744
rect 24394 28704 24400 28716
rect 24452 28704 24458 28756
rect 30098 28704 30104 28756
rect 30156 28744 30162 28756
rect 30285 28747 30343 28753
rect 30285 28744 30297 28747
rect 30156 28716 30297 28744
rect 30156 28704 30162 28716
rect 30285 28713 30297 28716
rect 30331 28713 30343 28747
rect 30285 28707 30343 28713
rect 31113 28747 31171 28753
rect 31113 28713 31125 28747
rect 31159 28744 31171 28747
rect 31386 28744 31392 28756
rect 31159 28716 31392 28744
rect 31159 28713 31171 28716
rect 31113 28707 31171 28713
rect 31386 28704 31392 28716
rect 31444 28704 31450 28756
rect 33594 28744 33600 28756
rect 33555 28716 33600 28744
rect 33594 28704 33600 28716
rect 33652 28704 33658 28756
rect 3973 28679 4031 28685
rect 3973 28645 3985 28679
rect 4019 28645 4031 28679
rect 24412 28676 24440 28704
rect 3973 28639 4031 28645
rect 23308 28648 24440 28676
rect 1394 28540 1400 28552
rect 1355 28512 1400 28540
rect 1394 28500 1400 28512
rect 1452 28500 1458 28552
rect 2593 28543 2651 28549
rect 2593 28509 2605 28543
rect 2639 28540 2651 28543
rect 2774 28540 2780 28552
rect 2639 28512 2780 28540
rect 2639 28509 2651 28512
rect 2593 28503 2651 28509
rect 2774 28500 2780 28512
rect 2832 28500 2838 28552
rect 3053 28543 3111 28549
rect 3053 28509 3065 28543
rect 3099 28540 3111 28543
rect 3988 28540 4016 28639
rect 4341 28611 4399 28617
rect 4341 28577 4353 28611
rect 4387 28608 4399 28611
rect 4798 28608 4804 28620
rect 4387 28580 4804 28608
rect 4387 28577 4399 28580
rect 4341 28571 4399 28577
rect 4798 28568 4804 28580
rect 4856 28568 4862 28620
rect 8662 28568 8668 28620
rect 8720 28608 8726 28620
rect 8941 28611 8999 28617
rect 8941 28608 8953 28611
rect 8720 28580 8953 28608
rect 8720 28568 8726 28580
rect 8941 28577 8953 28580
rect 8987 28577 8999 28611
rect 9766 28608 9772 28620
rect 9727 28580 9772 28608
rect 8941 28571 8999 28577
rect 9766 28568 9772 28580
rect 9824 28568 9830 28620
rect 12250 28568 12256 28620
rect 12308 28608 12314 28620
rect 12989 28611 13047 28617
rect 12989 28608 13001 28611
rect 12308 28580 13001 28608
rect 12308 28568 12314 28580
rect 12989 28577 13001 28580
rect 13035 28577 13047 28611
rect 12989 28571 13047 28577
rect 13814 28568 13820 28620
rect 13872 28608 13878 28620
rect 14645 28611 14703 28617
rect 14645 28608 14657 28611
rect 13872 28580 14657 28608
rect 13872 28568 13878 28580
rect 14645 28577 14657 28580
rect 14691 28577 14703 28611
rect 14645 28571 14703 28577
rect 14826 28568 14832 28620
rect 14884 28608 14890 28620
rect 14921 28611 14979 28617
rect 14921 28608 14933 28611
rect 14884 28580 14933 28608
rect 14884 28568 14890 28580
rect 14921 28577 14933 28580
rect 14967 28577 14979 28611
rect 14921 28571 14979 28577
rect 15657 28611 15715 28617
rect 15657 28577 15669 28611
rect 15703 28608 15715 28611
rect 16574 28608 16580 28620
rect 15703 28580 16580 28608
rect 15703 28577 15715 28580
rect 15657 28571 15715 28577
rect 16574 28568 16580 28580
rect 16632 28568 16638 28620
rect 23308 28617 23336 28648
rect 23293 28611 23351 28617
rect 23293 28577 23305 28611
rect 23339 28577 23351 28611
rect 23293 28571 23351 28577
rect 24026 28568 24032 28620
rect 24084 28608 24090 28620
rect 24489 28611 24547 28617
rect 24489 28608 24501 28611
rect 24084 28580 24501 28608
rect 24084 28568 24090 28580
rect 24489 28577 24501 28580
rect 24535 28577 24547 28611
rect 24489 28571 24547 28577
rect 29733 28611 29791 28617
rect 29733 28577 29745 28611
rect 29779 28608 29791 28611
rect 29822 28608 29828 28620
rect 29779 28580 29828 28608
rect 29779 28577 29791 28580
rect 29733 28571 29791 28577
rect 29822 28568 29828 28580
rect 29880 28568 29886 28620
rect 4154 28540 4160 28552
rect 3099 28512 4016 28540
rect 4115 28512 4160 28540
rect 3099 28509 3111 28512
rect 3053 28503 3111 28509
rect 4154 28500 4160 28512
rect 4212 28500 4218 28552
rect 4433 28543 4491 28549
rect 4433 28509 4445 28543
rect 4479 28540 4491 28543
rect 4706 28540 4712 28552
rect 4479 28512 4712 28540
rect 4479 28509 4491 28512
rect 4433 28503 4491 28509
rect 4706 28500 4712 28512
rect 4764 28500 4770 28552
rect 5258 28500 5264 28552
rect 5316 28540 5322 28552
rect 5721 28543 5779 28549
rect 5721 28540 5733 28543
rect 5316 28512 5733 28540
rect 5316 28500 5322 28512
rect 5721 28509 5733 28512
rect 5767 28540 5779 28543
rect 8110 28540 8116 28552
rect 5767 28512 8116 28540
rect 5767 28509 5779 28512
rect 5721 28503 5779 28509
rect 8110 28500 8116 28512
rect 8168 28500 8174 28552
rect 13078 28500 13084 28552
rect 13136 28540 13142 28552
rect 13265 28543 13323 28549
rect 13265 28540 13277 28543
rect 13136 28512 13277 28540
rect 13136 28500 13142 28512
rect 13265 28509 13277 28512
rect 13311 28509 13323 28543
rect 13265 28503 13323 28509
rect 15841 28543 15899 28549
rect 15841 28509 15853 28543
rect 15887 28540 15899 28543
rect 15930 28540 15936 28552
rect 15887 28512 15936 28540
rect 15887 28509 15899 28512
rect 15841 28503 15899 28509
rect 15930 28500 15936 28512
rect 15988 28500 15994 28552
rect 23017 28543 23075 28549
rect 23017 28540 23029 28543
rect 22756 28512 23029 28540
rect 5537 28475 5595 28481
rect 5537 28441 5549 28475
rect 5583 28441 5595 28475
rect 5537 28435 5595 28441
rect 9125 28475 9183 28481
rect 9125 28441 9137 28475
rect 9171 28472 9183 28475
rect 9214 28472 9220 28484
rect 9171 28444 9220 28472
rect 9171 28441 9183 28444
rect 9125 28435 9183 28441
rect 1581 28407 1639 28413
rect 1581 28373 1593 28407
rect 1627 28404 1639 28407
rect 2590 28404 2596 28416
rect 1627 28376 2596 28404
rect 1627 28373 1639 28376
rect 1581 28367 1639 28373
rect 2590 28364 2596 28376
rect 2648 28364 2654 28416
rect 4982 28404 4988 28416
rect 4943 28376 4988 28404
rect 4982 28364 4988 28376
rect 5040 28404 5046 28416
rect 5552 28404 5580 28435
rect 9214 28432 9220 28444
rect 9272 28432 9278 28484
rect 15565 28475 15623 28481
rect 15565 28441 15577 28475
rect 15611 28472 15623 28475
rect 17034 28472 17040 28484
rect 15611 28444 17040 28472
rect 15611 28441 15623 28444
rect 15565 28435 15623 28441
rect 17034 28432 17040 28444
rect 17092 28432 17098 28484
rect 22756 28416 22784 28512
rect 23017 28509 23029 28512
rect 23063 28509 23075 28543
rect 23017 28503 23075 28509
rect 24210 28500 24216 28552
rect 24268 28540 24274 28552
rect 24673 28543 24731 28549
rect 24673 28540 24685 28543
rect 24268 28512 24685 28540
rect 24268 28500 24274 28512
rect 24673 28509 24685 28512
rect 24719 28509 24731 28543
rect 25498 28540 25504 28552
rect 25459 28512 25504 28540
rect 24673 28503 24731 28509
rect 25498 28500 25504 28512
rect 25556 28500 25562 28552
rect 29638 28500 29644 28552
rect 29696 28540 29702 28552
rect 29914 28540 29920 28552
rect 29696 28512 29920 28540
rect 29696 28500 29702 28512
rect 29914 28500 29920 28512
rect 29972 28540 29978 28552
rect 35894 28540 35900 28552
rect 29972 28512 35900 28540
rect 29972 28500 29978 28512
rect 35894 28500 35900 28512
rect 35952 28540 35958 28552
rect 36354 28540 36360 28552
rect 35952 28512 36360 28540
rect 35952 28500 35958 28512
rect 36354 28500 36360 28512
rect 36412 28500 36418 28552
rect 23934 28432 23940 28484
rect 23992 28472 23998 28484
rect 24397 28475 24455 28481
rect 24397 28472 24409 28475
rect 23992 28444 24409 28472
rect 23992 28432 23998 28444
rect 24397 28441 24409 28444
rect 24443 28441 24455 28475
rect 24397 28435 24455 28441
rect 33689 28475 33747 28481
rect 33689 28441 33701 28475
rect 33735 28472 33747 28475
rect 33778 28472 33784 28484
rect 33735 28444 33784 28472
rect 33735 28441 33747 28444
rect 33689 28435 33747 28441
rect 33778 28432 33784 28444
rect 33836 28432 33842 28484
rect 5040 28376 5580 28404
rect 16025 28407 16083 28413
rect 5040 28364 5046 28376
rect 16025 28373 16037 28407
rect 16071 28404 16083 28407
rect 16850 28404 16856 28416
rect 16071 28376 16856 28404
rect 16071 28373 16083 28376
rect 16025 28367 16083 28373
rect 16850 28364 16856 28376
rect 16908 28364 16914 28416
rect 22557 28407 22615 28413
rect 22557 28373 22569 28407
rect 22603 28404 22615 28407
rect 22738 28404 22744 28416
rect 22603 28376 22744 28404
rect 22603 28373 22615 28376
rect 22557 28367 22615 28373
rect 22738 28364 22744 28376
rect 22796 28364 22802 28416
rect 24854 28404 24860 28416
rect 24815 28376 24860 28404
rect 24854 28364 24860 28376
rect 24912 28364 24918 28416
rect 29638 28364 29644 28416
rect 29696 28404 29702 28416
rect 29825 28407 29883 28413
rect 29825 28404 29837 28407
rect 29696 28376 29837 28404
rect 29696 28364 29702 28376
rect 29825 28373 29837 28376
rect 29871 28373 29883 28407
rect 29825 28367 29883 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 4706 28160 4712 28212
rect 4764 28200 4770 28212
rect 5077 28203 5135 28209
rect 5077 28200 5089 28203
rect 4764 28172 5089 28200
rect 4764 28160 4770 28172
rect 5077 28169 5089 28172
rect 5123 28169 5135 28203
rect 16574 28200 16580 28212
rect 5077 28163 5135 28169
rect 15488 28172 16580 28200
rect 1394 28132 1400 28144
rect 1355 28104 1400 28132
rect 1394 28092 1400 28104
rect 1452 28092 1458 28144
rect 2774 28064 2780 28076
rect 2735 28036 2780 28064
rect 2774 28024 2780 28036
rect 2832 28024 2838 28076
rect 5258 28064 5264 28076
rect 5219 28036 5264 28064
rect 5258 28024 5264 28036
rect 5316 28024 5322 28076
rect 9122 28064 9128 28076
rect 9083 28036 9128 28064
rect 9122 28024 9128 28036
rect 9180 28024 9186 28076
rect 14918 28064 14924 28076
rect 14879 28036 14924 28064
rect 14918 28024 14924 28036
rect 14976 28024 14982 28076
rect 2958 27996 2964 28008
rect 2919 27968 2964 27996
rect 2958 27956 2964 27968
rect 3016 27956 3022 28008
rect 3234 27996 3240 28008
rect 3195 27968 3240 27996
rect 3234 27956 3240 27968
rect 3292 27996 3298 28008
rect 9306 27996 9312 28008
rect 3292 27968 6914 27996
rect 9267 27968 9312 27996
rect 3292 27956 3298 27968
rect 6886 27928 6914 27968
rect 9306 27956 9312 27968
rect 9364 27956 9370 28008
rect 9677 27999 9735 28005
rect 9677 27965 9689 27999
rect 9723 27996 9735 27999
rect 12986 27996 12992 28008
rect 9723 27968 12992 27996
rect 9723 27965 9735 27968
rect 9677 27959 9735 27965
rect 9692 27928 9720 27959
rect 12986 27956 12992 27968
rect 13044 27956 13050 28008
rect 15488 27996 15516 28172
rect 16574 28160 16580 28172
rect 16632 28160 16638 28212
rect 29638 28200 29644 28212
rect 29599 28172 29644 28200
rect 29638 28160 29644 28172
rect 29696 28160 29702 28212
rect 30006 28200 30012 28212
rect 29967 28172 30012 28200
rect 30006 28160 30012 28172
rect 30064 28160 30070 28212
rect 34149 28203 34207 28209
rect 34149 28169 34161 28203
rect 34195 28200 34207 28203
rect 35434 28200 35440 28212
rect 34195 28172 35440 28200
rect 34195 28169 34207 28172
rect 34149 28163 34207 28169
rect 35434 28160 35440 28172
rect 35492 28160 35498 28212
rect 15841 28135 15899 28141
rect 15841 28101 15853 28135
rect 15887 28132 15899 28135
rect 17034 28132 17040 28144
rect 15887 28104 17040 28132
rect 15887 28101 15899 28104
rect 15841 28095 15899 28101
rect 17034 28092 17040 28104
rect 17092 28092 17098 28144
rect 23658 28132 23664 28144
rect 23619 28104 23664 28132
rect 23658 28092 23664 28104
rect 23716 28092 23722 28144
rect 32490 28132 32496 28144
rect 32451 28104 32496 28132
rect 32490 28092 32496 28104
rect 32548 28092 32554 28144
rect 15565 28067 15623 28073
rect 15565 28033 15577 28067
rect 15611 28064 15623 28067
rect 15930 28064 15936 28076
rect 15611 28036 15936 28064
rect 15611 28033 15623 28036
rect 15565 28027 15623 28033
rect 15930 28024 15936 28036
rect 15988 28024 15994 28076
rect 16850 28064 16856 28076
rect 16811 28036 16856 28064
rect 16850 28024 16856 28036
rect 16908 28024 16914 28076
rect 25498 28024 25504 28076
rect 25556 28064 25562 28076
rect 27249 28067 27307 28073
rect 25556 28036 25601 28064
rect 25556 28024 25562 28036
rect 27249 28033 27261 28067
rect 27295 28064 27307 28067
rect 28810 28064 28816 28076
rect 27295 28036 28816 28064
rect 27295 28033 27307 28036
rect 27249 28027 27307 28033
rect 28810 28024 28816 28036
rect 28868 28024 28874 28076
rect 32214 28024 32220 28076
rect 32272 28064 32278 28076
rect 32677 28067 32735 28073
rect 32677 28064 32689 28067
rect 32272 28036 32689 28064
rect 32272 28024 32278 28036
rect 32677 28033 32689 28036
rect 32723 28033 32735 28067
rect 32677 28027 32735 28033
rect 33318 28024 33324 28076
rect 33376 28064 33382 28076
rect 33965 28067 34023 28073
rect 33965 28064 33977 28067
rect 33376 28036 33977 28064
rect 33376 28024 33382 28036
rect 33965 28033 33977 28036
rect 34011 28033 34023 28067
rect 33965 28027 34023 28033
rect 15657 27999 15715 28005
rect 15657 27996 15669 27999
rect 15488 27968 15669 27996
rect 15657 27965 15669 27968
rect 15703 27965 15715 27999
rect 15657 27959 15715 27965
rect 18874 27956 18880 28008
rect 18932 27996 18938 28008
rect 19429 27999 19487 28005
rect 19429 27996 19441 27999
rect 18932 27968 19441 27996
rect 18932 27956 18938 27968
rect 19429 27965 19441 27968
rect 19475 27965 19487 27999
rect 19429 27959 19487 27965
rect 19705 27999 19763 28005
rect 19705 27965 19717 27999
rect 19751 27996 19763 27999
rect 21634 27996 21640 28008
rect 19751 27968 21640 27996
rect 19751 27965 19763 27968
rect 19705 27959 19763 27965
rect 21634 27956 21640 27968
rect 21692 27956 21698 28008
rect 25314 27996 25320 28008
rect 25275 27968 25320 27996
rect 25314 27956 25320 27968
rect 25372 27956 25378 28008
rect 26234 27956 26240 28008
rect 26292 27996 26298 28008
rect 26973 27999 27031 28005
rect 26973 27996 26985 27999
rect 26292 27968 26985 27996
rect 26292 27956 26298 27968
rect 26973 27965 26985 27968
rect 27019 27965 27031 27999
rect 26973 27959 27031 27965
rect 29730 27956 29736 28008
rect 29788 27996 29794 28008
rect 30101 27999 30159 28005
rect 30101 27996 30113 27999
rect 29788 27968 30113 27996
rect 29788 27956 29794 27968
rect 30101 27965 30113 27968
rect 30147 27965 30159 27999
rect 30101 27959 30159 27965
rect 30285 27999 30343 28005
rect 30285 27965 30297 27999
rect 30331 27996 30343 27999
rect 30834 27996 30840 28008
rect 30331 27968 30840 27996
rect 30331 27965 30343 27968
rect 30285 27959 30343 27965
rect 30834 27956 30840 27968
rect 30892 27956 30898 28008
rect 33594 27956 33600 28008
rect 33652 27996 33658 28008
rect 33781 27999 33839 28005
rect 33781 27996 33793 27999
rect 33652 27968 33793 27996
rect 33652 27956 33658 27968
rect 33781 27965 33793 27968
rect 33827 27965 33839 27999
rect 33781 27959 33839 27965
rect 15838 27928 15844 27940
rect 6886 27900 9720 27928
rect 15580 27900 15844 27928
rect 13078 27820 13084 27872
rect 13136 27860 13142 27872
rect 13357 27863 13415 27869
rect 13357 27860 13369 27863
rect 13136 27832 13369 27860
rect 13136 27820 13142 27832
rect 13357 27829 13369 27832
rect 13403 27829 13415 27863
rect 14274 27860 14280 27872
rect 14235 27832 14280 27860
rect 13357 27823 13415 27829
rect 14274 27820 14280 27832
rect 14332 27820 14338 27872
rect 14458 27820 14464 27872
rect 14516 27860 14522 27872
rect 14737 27863 14795 27869
rect 14737 27860 14749 27863
rect 14516 27832 14749 27860
rect 14516 27820 14522 27832
rect 14737 27829 14749 27832
rect 14783 27829 14795 27863
rect 15378 27860 15384 27872
rect 15339 27832 15384 27860
rect 14737 27823 14795 27829
rect 15378 27820 15384 27832
rect 15436 27820 15442 27872
rect 15580 27869 15608 27900
rect 15838 27888 15844 27900
rect 15896 27928 15902 27940
rect 16482 27928 16488 27940
rect 15896 27900 16488 27928
rect 15896 27888 15902 27900
rect 16482 27888 16488 27900
rect 16540 27888 16546 27940
rect 15565 27863 15623 27869
rect 15565 27829 15577 27863
rect 15611 27829 15623 27863
rect 15565 27823 15623 27829
rect 15654 27820 15660 27872
rect 15712 27860 15718 27872
rect 16669 27863 16727 27869
rect 16669 27860 16681 27863
rect 15712 27832 16681 27860
rect 15712 27820 15718 27832
rect 16669 27829 16681 27832
rect 16715 27829 16727 27863
rect 20714 27860 20720 27872
rect 20675 27832 20720 27860
rect 16669 27823 16727 27829
rect 20714 27820 20720 27832
rect 20772 27820 20778 27872
rect 26142 27860 26148 27872
rect 26103 27832 26148 27860
rect 26142 27820 26148 27832
rect 26200 27820 26206 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 2958 27616 2964 27668
rect 3016 27656 3022 27668
rect 3053 27659 3111 27665
rect 3053 27656 3065 27659
rect 3016 27628 3065 27656
rect 3016 27616 3022 27628
rect 3053 27625 3065 27628
rect 3099 27625 3111 27659
rect 3053 27619 3111 27625
rect 4249 27659 4307 27665
rect 4249 27625 4261 27659
rect 4295 27656 4307 27659
rect 4614 27656 4620 27668
rect 4295 27628 4620 27656
rect 4295 27625 4307 27628
rect 4249 27619 4307 27625
rect 4614 27616 4620 27628
rect 4672 27656 4678 27668
rect 5074 27656 5080 27668
rect 4672 27628 5080 27656
rect 4672 27616 4678 27628
rect 5074 27616 5080 27628
rect 5132 27616 5138 27668
rect 16482 27616 16488 27668
rect 16540 27656 16546 27668
rect 16853 27659 16911 27665
rect 16853 27656 16865 27659
rect 16540 27628 16865 27656
rect 16540 27616 16546 27628
rect 16853 27625 16865 27628
rect 16899 27625 16911 27659
rect 16853 27619 16911 27625
rect 29730 27616 29736 27668
rect 29788 27656 29794 27668
rect 29788 27628 34652 27656
rect 29788 27616 29794 27628
rect 3789 27591 3847 27597
rect 3789 27557 3801 27591
rect 3835 27557 3847 27591
rect 3789 27551 3847 27557
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27452 3295 27455
rect 3804 27452 3832 27551
rect 9306 27548 9312 27600
rect 9364 27588 9370 27600
rect 10321 27591 10379 27597
rect 10321 27588 10333 27591
rect 9364 27560 10333 27588
rect 9364 27548 9370 27560
rect 10321 27557 10333 27560
rect 10367 27557 10379 27591
rect 10321 27551 10379 27557
rect 23845 27591 23903 27597
rect 23845 27557 23857 27591
rect 23891 27588 23903 27591
rect 25314 27588 25320 27600
rect 23891 27560 25320 27588
rect 23891 27557 23903 27560
rect 23845 27551 23903 27557
rect 25314 27548 25320 27560
rect 25372 27548 25378 27600
rect 26142 27548 26148 27600
rect 26200 27588 26206 27600
rect 33873 27591 33931 27597
rect 26200 27560 26280 27588
rect 26200 27548 26206 27560
rect 4157 27523 4215 27529
rect 4157 27489 4169 27523
rect 4203 27520 4215 27523
rect 4614 27520 4620 27532
rect 4203 27492 4620 27520
rect 4203 27489 4215 27492
rect 4157 27483 4215 27489
rect 4614 27480 4620 27492
rect 4672 27520 4678 27532
rect 4798 27520 4804 27532
rect 4672 27492 4804 27520
rect 4672 27480 4678 27492
rect 4798 27480 4804 27492
rect 4856 27480 4862 27532
rect 14274 27480 14280 27532
rect 14332 27520 14338 27532
rect 14553 27523 14611 27529
rect 14553 27520 14565 27523
rect 14332 27492 14565 27520
rect 14332 27480 14338 27492
rect 14553 27489 14565 27492
rect 14599 27489 14611 27523
rect 14553 27483 14611 27489
rect 14737 27523 14795 27529
rect 14737 27489 14749 27523
rect 14783 27520 14795 27523
rect 15654 27520 15660 27532
rect 14783 27492 15660 27520
rect 14783 27489 14795 27492
rect 14737 27483 14795 27489
rect 15654 27480 15660 27492
rect 15712 27480 15718 27532
rect 15746 27480 15752 27532
rect 15804 27520 15810 27532
rect 15804 27492 15849 27520
rect 15804 27480 15810 27492
rect 16574 27480 16580 27532
rect 16632 27520 16638 27532
rect 17037 27523 17095 27529
rect 17037 27520 17049 27523
rect 16632 27492 17049 27520
rect 16632 27480 16638 27492
rect 17037 27489 17049 27492
rect 17083 27520 17095 27523
rect 17678 27520 17684 27532
rect 17083 27492 17684 27520
rect 17083 27489 17095 27492
rect 17037 27483 17095 27489
rect 17678 27480 17684 27492
rect 17736 27480 17742 27532
rect 19981 27523 20039 27529
rect 19981 27489 19993 27523
rect 20027 27520 20039 27523
rect 24026 27520 24032 27532
rect 20027 27492 24032 27520
rect 20027 27489 20039 27492
rect 19981 27483 20039 27489
rect 24026 27480 24032 27492
rect 24084 27480 24090 27532
rect 24302 27480 24308 27532
rect 24360 27520 24366 27532
rect 26252 27529 26280 27560
rect 33873 27557 33885 27591
rect 33919 27588 33931 27591
rect 34514 27588 34520 27600
rect 33919 27560 34520 27588
rect 33919 27557 33931 27560
rect 33873 27551 33931 27557
rect 34514 27548 34520 27560
rect 34572 27548 34578 27600
rect 26053 27523 26111 27529
rect 26053 27520 26065 27523
rect 24360 27492 26065 27520
rect 24360 27480 24366 27492
rect 26053 27489 26065 27492
rect 26099 27489 26111 27523
rect 26053 27483 26111 27489
rect 26237 27523 26295 27529
rect 26237 27489 26249 27523
rect 26283 27489 26295 27523
rect 26237 27483 26295 27489
rect 26973 27523 27031 27529
rect 26973 27489 26985 27523
rect 27019 27520 27031 27523
rect 28902 27520 28908 27532
rect 27019 27492 28908 27520
rect 27019 27489 27031 27492
rect 26973 27483 27031 27489
rect 28902 27480 28908 27492
rect 28960 27480 28966 27532
rect 33505 27523 33563 27529
rect 33505 27489 33517 27523
rect 33551 27520 33563 27523
rect 33594 27520 33600 27532
rect 33551 27492 33600 27520
rect 33551 27489 33563 27492
rect 33505 27483 33563 27489
rect 33594 27480 33600 27492
rect 33652 27480 33658 27532
rect 3283 27424 3832 27452
rect 3973 27455 4031 27461
rect 3283 27421 3295 27424
rect 3237 27415 3295 27421
rect 3973 27421 3985 27455
rect 4019 27452 4031 27455
rect 4249 27455 4307 27461
rect 4019 27424 4200 27452
rect 4019 27421 4031 27424
rect 3973 27415 4031 27421
rect 4172 27396 4200 27424
rect 4249 27421 4261 27455
rect 4295 27452 4307 27455
rect 4706 27452 4712 27464
rect 4295 27424 4712 27452
rect 4295 27421 4307 27424
rect 4249 27415 4307 27421
rect 4706 27412 4712 27424
rect 4764 27412 4770 27464
rect 9030 27452 9036 27464
rect 8991 27424 9036 27452
rect 9030 27412 9036 27424
rect 9088 27412 9094 27464
rect 9214 27412 9220 27464
rect 9272 27452 9278 27464
rect 9309 27455 9367 27461
rect 9309 27452 9321 27455
rect 9272 27424 9321 27452
rect 9272 27412 9278 27424
rect 9309 27421 9321 27424
rect 9355 27421 9367 27455
rect 9309 27415 9367 27421
rect 9766 27412 9772 27464
rect 9824 27452 9830 27464
rect 10505 27455 10563 27461
rect 10505 27452 10517 27455
rect 9824 27424 10517 27452
rect 9824 27412 9830 27424
rect 10505 27421 10517 27424
rect 10551 27421 10563 27455
rect 10505 27415 10563 27421
rect 11149 27455 11207 27461
rect 11149 27421 11161 27455
rect 11195 27452 11207 27455
rect 11422 27452 11428 27464
rect 11195 27424 11428 27452
rect 11195 27421 11207 27424
rect 11149 27415 11207 27421
rect 11422 27412 11428 27424
rect 11480 27412 11486 27464
rect 15930 27412 15936 27464
rect 15988 27452 15994 27464
rect 17129 27455 17187 27461
rect 17129 27452 17141 27455
rect 15988 27424 17141 27452
rect 15988 27412 15994 27424
rect 17129 27421 17141 27424
rect 17175 27421 17187 27455
rect 17865 27455 17923 27461
rect 17865 27452 17877 27455
rect 17129 27415 17187 27421
rect 17328 27424 17877 27452
rect 4154 27344 4160 27396
rect 4212 27344 4218 27396
rect 16853 27387 16911 27393
rect 16853 27353 16865 27387
rect 16899 27384 16911 27387
rect 17034 27384 17040 27396
rect 16899 27356 17040 27384
rect 16899 27353 16911 27356
rect 16853 27347 16911 27353
rect 17034 27344 17040 27356
rect 17092 27344 17098 27396
rect 17328 27325 17356 27424
rect 17865 27421 17877 27424
rect 17911 27421 17923 27455
rect 18506 27452 18512 27464
rect 18467 27424 18512 27452
rect 17865 27415 17923 27421
rect 18506 27412 18512 27424
rect 18564 27412 18570 27464
rect 19334 27412 19340 27464
rect 19392 27452 19398 27464
rect 20441 27455 20499 27461
rect 20441 27452 20453 27455
rect 19392 27424 20453 27452
rect 19392 27412 19398 27424
rect 20441 27421 20453 27424
rect 20487 27452 20499 27455
rect 20622 27452 20628 27464
rect 20487 27424 20628 27452
rect 20487 27421 20499 27424
rect 20441 27415 20499 27421
rect 20622 27412 20628 27424
rect 20680 27412 20686 27464
rect 20717 27455 20775 27461
rect 20717 27421 20729 27455
rect 20763 27452 20775 27455
rect 21358 27452 21364 27464
rect 20763 27424 21364 27452
rect 20763 27421 20775 27424
rect 20717 27415 20775 27421
rect 21358 27412 21364 27424
rect 21416 27412 21422 27464
rect 23661 27455 23719 27461
rect 23661 27421 23673 27455
rect 23707 27452 23719 27455
rect 24854 27452 24860 27464
rect 23707 27424 24860 27452
rect 23707 27421 23719 27424
rect 23661 27415 23719 27421
rect 24854 27412 24860 27424
rect 24912 27412 24918 27464
rect 26694 27452 26700 27464
rect 26655 27424 26700 27452
rect 26694 27412 26700 27424
rect 26752 27412 26758 27464
rect 33686 27452 33692 27464
rect 33647 27424 33692 27452
rect 33686 27412 33692 27424
rect 33744 27412 33750 27464
rect 34624 27452 34652 27628
rect 35805 27523 35863 27529
rect 35805 27489 35817 27523
rect 35851 27520 35863 27523
rect 35986 27520 35992 27532
rect 35851 27492 35992 27520
rect 35851 27489 35863 27492
rect 35805 27483 35863 27489
rect 35986 27480 35992 27492
rect 36044 27480 36050 27532
rect 36998 27520 37004 27532
rect 36959 27492 37004 27520
rect 36998 27480 37004 27492
rect 37056 27480 37062 27532
rect 35529 27455 35587 27461
rect 35529 27452 35541 27455
rect 34624 27424 35541 27452
rect 35529 27421 35541 27424
rect 35575 27421 35587 27455
rect 35529 27415 35587 27421
rect 35621 27455 35679 27461
rect 35621 27421 35633 27455
rect 35667 27452 35679 27455
rect 36170 27452 36176 27464
rect 35667 27424 36176 27452
rect 35667 27421 35679 27424
rect 35621 27415 35679 27421
rect 19426 27344 19432 27396
rect 19484 27384 19490 27396
rect 19797 27387 19855 27393
rect 19797 27384 19809 27387
rect 19484 27356 19809 27384
rect 19484 27344 19490 27356
rect 19797 27353 19809 27356
rect 19843 27384 19855 27387
rect 20254 27384 20260 27396
rect 19843 27356 20260 27384
rect 19843 27353 19855 27356
rect 19797 27347 19855 27353
rect 20254 27344 20260 27356
rect 20312 27344 20318 27396
rect 24397 27387 24455 27393
rect 24397 27353 24409 27387
rect 24443 27384 24455 27387
rect 24670 27384 24676 27396
rect 24443 27356 24676 27384
rect 24443 27353 24455 27356
rect 24397 27347 24455 27353
rect 24670 27344 24676 27356
rect 24728 27384 24734 27396
rect 25038 27384 25044 27396
rect 24728 27356 25044 27384
rect 24728 27344 24734 27356
rect 25038 27344 25044 27356
rect 25096 27344 25102 27396
rect 35544 27384 35572 27415
rect 36170 27412 36176 27424
rect 36228 27412 36234 27464
rect 36725 27455 36783 27461
rect 36725 27421 36737 27455
rect 36771 27452 36783 27455
rect 37642 27452 37648 27464
rect 36771 27424 37648 27452
rect 36771 27421 36783 27424
rect 36725 27415 36783 27421
rect 37642 27412 37648 27424
rect 37700 27412 37706 27464
rect 36078 27384 36084 27396
rect 35544 27356 36084 27384
rect 36078 27344 36084 27356
rect 36136 27344 36142 27396
rect 17313 27319 17371 27325
rect 17313 27285 17325 27319
rect 17359 27285 17371 27319
rect 17313 27279 17371 27285
rect 18049 27319 18107 27325
rect 18049 27285 18061 27319
rect 18095 27316 18107 27319
rect 18690 27316 18696 27328
rect 18095 27288 18696 27316
rect 18095 27285 18107 27288
rect 18049 27279 18107 27285
rect 18690 27276 18696 27288
rect 18748 27276 18754 27328
rect 31938 27276 31944 27328
rect 31996 27316 32002 27328
rect 32033 27319 32091 27325
rect 32033 27316 32045 27319
rect 31996 27288 32045 27316
rect 31996 27276 32002 27288
rect 32033 27285 32045 27288
rect 32079 27285 32091 27319
rect 32033 27279 32091 27285
rect 33226 27276 33232 27328
rect 33284 27316 33290 27328
rect 35161 27319 35219 27325
rect 35161 27316 35173 27319
rect 33284 27288 35173 27316
rect 33284 27276 33290 27288
rect 35161 27285 35173 27288
rect 35207 27285 35219 27319
rect 35161 27279 35219 27285
rect 35618 27276 35624 27328
rect 35676 27316 35682 27328
rect 36357 27319 36415 27325
rect 36357 27316 36369 27319
rect 35676 27288 36369 27316
rect 35676 27276 35682 27288
rect 36357 27285 36369 27288
rect 36403 27285 36415 27319
rect 36357 27279 36415 27285
rect 36814 27276 36820 27328
rect 36872 27316 36878 27328
rect 36872 27288 36917 27316
rect 36872 27276 36878 27288
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 9766 27112 9772 27124
rect 9727 27084 9772 27112
rect 9766 27072 9772 27084
rect 9824 27072 9830 27124
rect 24118 27072 24124 27124
rect 24176 27112 24182 27124
rect 24397 27115 24455 27121
rect 24397 27112 24409 27115
rect 24176 27084 24409 27112
rect 24176 27072 24182 27084
rect 24397 27081 24409 27084
rect 24443 27081 24455 27115
rect 24397 27075 24455 27081
rect 31386 27072 31392 27124
rect 31444 27112 31450 27124
rect 31481 27115 31539 27121
rect 31481 27112 31493 27115
rect 31444 27084 31493 27112
rect 31444 27072 31450 27084
rect 31481 27081 31493 27084
rect 31527 27112 31539 27115
rect 31662 27112 31668 27124
rect 31527 27084 31668 27112
rect 31527 27081 31539 27084
rect 31481 27075 31539 27081
rect 31662 27072 31668 27084
rect 31720 27112 31726 27124
rect 32769 27115 32827 27121
rect 31720 27084 32628 27112
rect 31720 27072 31726 27084
rect 9309 27047 9367 27053
rect 9309 27013 9321 27047
rect 9355 27044 9367 27047
rect 9490 27044 9496 27056
rect 9355 27016 9496 27044
rect 9355 27013 9367 27016
rect 9309 27007 9367 27013
rect 9490 27004 9496 27016
rect 9548 27004 9554 27056
rect 14458 27044 14464 27056
rect 14419 27016 14464 27044
rect 14458 27004 14464 27016
rect 14516 27004 14522 27056
rect 18690 27044 18696 27056
rect 18651 27016 18696 27044
rect 18690 27004 18696 27016
rect 18748 27004 18754 27056
rect 23934 27044 23940 27056
rect 23895 27016 23940 27044
rect 23934 27004 23940 27016
rect 23992 27004 23998 27056
rect 31938 27004 31944 27056
rect 31996 27044 32002 27056
rect 32493 27047 32551 27053
rect 32493 27044 32505 27047
rect 31996 27016 32505 27044
rect 31996 27004 32002 27016
rect 32493 27013 32505 27016
rect 32539 27013 32551 27047
rect 32493 27007 32551 27013
rect 1394 26976 1400 26988
rect 1355 26948 1400 26976
rect 1394 26936 1400 26948
rect 1452 26976 1458 26988
rect 2041 26979 2099 26985
rect 2041 26976 2053 26979
rect 1452 26948 2053 26976
rect 1452 26936 1458 26948
rect 2041 26945 2053 26948
rect 2087 26945 2099 26979
rect 9582 26976 9588 26988
rect 9543 26948 9588 26976
rect 2041 26939 2099 26945
rect 9582 26936 9588 26948
rect 9640 26936 9646 26988
rect 10410 26976 10416 26988
rect 10371 26948 10416 26976
rect 10410 26936 10416 26948
rect 10468 26936 10474 26988
rect 17221 26979 17279 26985
rect 17221 26945 17233 26979
rect 17267 26976 17279 26979
rect 18046 26976 18052 26988
rect 17267 26948 18052 26976
rect 17267 26945 17279 26948
rect 17221 26939 17279 26945
rect 18046 26936 18052 26948
rect 18104 26936 18110 26988
rect 18506 26976 18512 26988
rect 18467 26948 18512 26976
rect 18506 26936 18512 26948
rect 18564 26936 18570 26988
rect 24210 26976 24216 26988
rect 24171 26948 24216 26976
rect 24210 26936 24216 26948
rect 24268 26936 24274 26988
rect 29825 26979 29883 26985
rect 29825 26945 29837 26979
rect 29871 26976 29883 26979
rect 30006 26976 30012 26988
rect 29871 26948 30012 26976
rect 29871 26945 29883 26948
rect 29825 26939 29883 26945
rect 30006 26936 30012 26948
rect 30064 26936 30070 26988
rect 32214 26976 32220 26988
rect 32175 26948 32220 26976
rect 32214 26936 32220 26948
rect 32272 26936 32278 26988
rect 32398 26976 32404 26988
rect 32359 26948 32404 26976
rect 32398 26936 32404 26948
rect 32456 26936 32462 26988
rect 32600 26985 32628 27084
rect 32769 27081 32781 27115
rect 32815 27112 32827 27115
rect 33686 27112 33692 27124
rect 32815 27084 33692 27112
rect 32815 27081 32827 27084
rect 32769 27075 32827 27081
rect 33686 27072 33692 27084
rect 33744 27072 33750 27124
rect 34054 27112 34060 27124
rect 34015 27084 34060 27112
rect 34054 27072 34060 27084
rect 34112 27072 34118 27124
rect 36725 27115 36783 27121
rect 36725 27081 36737 27115
rect 36771 27112 36783 27115
rect 36814 27112 36820 27124
rect 36771 27084 36820 27112
rect 36771 27081 36783 27084
rect 36725 27075 36783 27081
rect 36814 27072 36820 27084
rect 36872 27072 36878 27124
rect 37182 27004 37188 27056
rect 37240 27044 37246 27056
rect 37645 27047 37703 27053
rect 37645 27044 37657 27047
rect 37240 27016 37657 27044
rect 37240 27004 37246 27016
rect 37645 27013 37657 27016
rect 37691 27013 37703 27047
rect 37645 27007 37703 27013
rect 32585 26979 32643 26985
rect 32585 26945 32597 26979
rect 32631 26945 32643 26979
rect 32585 26939 32643 26945
rect 33965 26979 34023 26985
rect 33965 26945 33977 26979
rect 34011 26976 34023 26979
rect 34793 26979 34851 26985
rect 34793 26976 34805 26979
rect 34011 26948 34805 26976
rect 34011 26945 34023 26948
rect 33965 26939 34023 26945
rect 9214 26868 9220 26920
rect 9272 26908 9278 26920
rect 9398 26908 9404 26920
rect 9272 26880 9404 26908
rect 9272 26868 9278 26880
rect 9398 26868 9404 26880
rect 9456 26868 9462 26920
rect 14274 26908 14280 26920
rect 14235 26880 14280 26908
rect 14274 26868 14280 26880
rect 14332 26868 14338 26920
rect 14737 26911 14795 26917
rect 14737 26877 14749 26911
rect 14783 26908 14795 26911
rect 15746 26908 15752 26920
rect 14783 26880 15752 26908
rect 14783 26877 14795 26880
rect 14737 26871 14795 26877
rect 3970 26800 3976 26852
rect 4028 26840 4034 26852
rect 5534 26840 5540 26852
rect 4028 26812 5540 26840
rect 4028 26800 4034 26812
rect 5534 26800 5540 26812
rect 5592 26800 5598 26852
rect 11882 26800 11888 26852
rect 11940 26840 11946 26852
rect 14752 26840 14780 26871
rect 15746 26868 15752 26880
rect 15804 26868 15810 26920
rect 17497 26911 17555 26917
rect 17497 26877 17509 26911
rect 17543 26908 17555 26911
rect 17678 26908 17684 26920
rect 17543 26880 17684 26908
rect 17543 26877 17555 26880
rect 17497 26871 17555 26877
rect 17678 26868 17684 26880
rect 17736 26868 17742 26920
rect 19426 26908 19432 26920
rect 19387 26880 19432 26908
rect 19426 26868 19432 26880
rect 19484 26868 19490 26920
rect 24026 26908 24032 26920
rect 23987 26880 24032 26908
rect 24026 26868 24032 26880
rect 24084 26908 24090 26920
rect 24486 26908 24492 26920
rect 24084 26880 24492 26908
rect 24084 26868 24090 26880
rect 24486 26868 24492 26880
rect 24544 26868 24550 26920
rect 27982 26908 27988 26920
rect 27943 26880 27988 26908
rect 27982 26868 27988 26880
rect 28040 26868 28046 26920
rect 28074 26868 28080 26920
rect 28132 26908 28138 26920
rect 29641 26911 29699 26917
rect 29641 26908 29653 26911
rect 28132 26880 29653 26908
rect 28132 26868 28138 26880
rect 29641 26877 29653 26880
rect 29687 26877 29699 26911
rect 29641 26871 29699 26877
rect 11940 26812 14780 26840
rect 11940 26800 11946 26812
rect 31386 26800 31392 26852
rect 31444 26840 31450 26852
rect 34054 26840 34060 26852
rect 31444 26812 34060 26840
rect 31444 26800 31450 26812
rect 34054 26800 34060 26812
rect 34112 26800 34118 26852
rect 1578 26772 1584 26784
rect 1539 26744 1584 26772
rect 1578 26732 1584 26744
rect 1636 26732 1642 26784
rect 4706 26772 4712 26784
rect 4667 26744 4712 26772
rect 4706 26732 4712 26744
rect 4764 26732 4770 26784
rect 5166 26772 5172 26784
rect 5127 26744 5172 26772
rect 5166 26732 5172 26744
rect 5224 26732 5230 26784
rect 9398 26772 9404 26784
rect 9359 26744 9404 26772
rect 9398 26732 9404 26744
rect 9456 26732 9462 26784
rect 10597 26775 10655 26781
rect 10597 26741 10609 26775
rect 10643 26772 10655 26775
rect 11606 26772 11612 26784
rect 10643 26744 11612 26772
rect 10643 26741 10655 26744
rect 10597 26735 10655 26741
rect 11606 26732 11612 26744
rect 11664 26732 11670 26784
rect 24213 26775 24271 26781
rect 24213 26741 24225 26775
rect 24259 26772 24271 26775
rect 24394 26772 24400 26784
rect 24259 26744 24400 26772
rect 24259 26741 24271 26744
rect 24213 26735 24271 26741
rect 24394 26732 24400 26744
rect 24452 26732 24458 26784
rect 33502 26732 33508 26784
rect 33560 26772 33566 26784
rect 33597 26775 33655 26781
rect 33597 26772 33609 26775
rect 33560 26744 33609 26772
rect 33560 26732 33566 26744
rect 33597 26741 33609 26744
rect 33643 26741 33655 26775
rect 34164 26772 34192 26948
rect 34793 26945 34805 26948
rect 34839 26945 34851 26979
rect 34793 26939 34851 26945
rect 36357 26979 36415 26985
rect 36357 26945 36369 26979
rect 36403 26976 36415 26979
rect 36446 26976 36452 26988
rect 36403 26948 36452 26976
rect 36403 26945 36415 26948
rect 36357 26939 36415 26945
rect 36446 26936 36452 26948
rect 36504 26936 36510 26988
rect 37090 26936 37096 26988
rect 37148 26976 37154 26988
rect 37829 26979 37887 26985
rect 37829 26976 37841 26979
rect 37148 26948 37841 26976
rect 37148 26936 37154 26948
rect 37829 26945 37841 26948
rect 37875 26945 37887 26979
rect 37829 26939 37887 26945
rect 34241 26911 34299 26917
rect 34241 26877 34253 26911
rect 34287 26908 34299 26911
rect 34287 26880 35894 26908
rect 34287 26877 34299 26880
rect 34241 26871 34299 26877
rect 35866 26840 35894 26880
rect 35986 26868 35992 26920
rect 36044 26908 36050 26920
rect 36081 26911 36139 26917
rect 36081 26908 36093 26911
rect 36044 26880 36093 26908
rect 36044 26868 36050 26880
rect 36081 26877 36093 26880
rect 36127 26877 36139 26911
rect 36081 26871 36139 26877
rect 36170 26868 36176 26920
rect 36228 26908 36234 26920
rect 36265 26911 36323 26917
rect 36265 26908 36277 26911
rect 36228 26880 36277 26908
rect 36228 26868 36234 26880
rect 36265 26877 36277 26880
rect 36311 26877 36323 26911
rect 36265 26871 36323 26877
rect 37182 26840 37188 26852
rect 35866 26812 37188 26840
rect 37182 26800 37188 26812
rect 37240 26800 37246 26852
rect 35894 26772 35900 26784
rect 34164 26744 35900 26772
rect 33597 26735 33655 26741
rect 35894 26732 35900 26744
rect 35952 26732 35958 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 4525 26571 4583 26577
rect 4525 26537 4537 26571
rect 4571 26568 4583 26571
rect 4614 26568 4620 26580
rect 4571 26540 4620 26568
rect 4571 26537 4583 26540
rect 4525 26531 4583 26537
rect 4614 26528 4620 26540
rect 4672 26528 4678 26580
rect 11882 26568 11888 26580
rect 6886 26540 11888 26568
rect 5534 26460 5540 26512
rect 5592 26500 5598 26512
rect 6886 26500 6914 26540
rect 11882 26528 11888 26540
rect 11940 26528 11946 26580
rect 14274 26528 14280 26580
rect 14332 26568 14338 26580
rect 14369 26571 14427 26577
rect 14369 26568 14381 26571
rect 14332 26540 14381 26568
rect 14332 26528 14338 26540
rect 14369 26537 14381 26540
rect 14415 26537 14427 26571
rect 14369 26531 14427 26537
rect 14918 26528 14924 26580
rect 14976 26568 14982 26580
rect 16117 26571 16175 26577
rect 16117 26568 16129 26571
rect 14976 26540 16129 26568
rect 14976 26528 14982 26540
rect 16117 26537 16129 26540
rect 16163 26537 16175 26571
rect 16482 26568 16488 26580
rect 16443 26540 16488 26568
rect 16117 26531 16175 26537
rect 16482 26528 16488 26540
rect 16540 26528 16546 26580
rect 18046 26568 18052 26580
rect 18007 26540 18052 26568
rect 18046 26528 18052 26540
rect 18104 26568 18110 26580
rect 18414 26568 18420 26580
rect 18104 26540 18420 26568
rect 18104 26528 18110 26540
rect 18414 26528 18420 26540
rect 18472 26528 18478 26580
rect 32398 26528 32404 26580
rect 32456 26568 32462 26580
rect 33045 26571 33103 26577
rect 33045 26568 33057 26571
rect 32456 26540 33057 26568
rect 32456 26528 32462 26540
rect 33045 26537 33057 26540
rect 33091 26537 33103 26571
rect 36446 26568 36452 26580
rect 36407 26540 36452 26568
rect 33045 26531 33103 26537
rect 36446 26528 36452 26540
rect 36504 26528 36510 26580
rect 5592 26472 6914 26500
rect 5592 26460 5598 26472
rect 5166 26432 5172 26444
rect 5127 26404 5172 26432
rect 5166 26392 5172 26404
rect 5224 26392 5230 26444
rect 6825 26435 6883 26441
rect 6825 26401 6837 26435
rect 6871 26401 6883 26435
rect 11422 26432 11428 26444
rect 11383 26404 11428 26432
rect 6825 26395 6883 26401
rect 4709 26367 4767 26373
rect 4709 26333 4721 26367
rect 4755 26333 4767 26367
rect 4709 26327 4767 26333
rect 4724 26296 4752 26327
rect 5350 26296 5356 26308
rect 4724 26268 5212 26296
rect 5311 26268 5356 26296
rect 5184 26228 5212 26268
rect 5350 26256 5356 26268
rect 5408 26256 5414 26308
rect 5626 26256 5632 26308
rect 5684 26296 5690 26308
rect 6840 26296 6868 26395
rect 11422 26392 11428 26404
rect 11480 26392 11486 26444
rect 11606 26432 11612 26444
rect 11567 26404 11612 26432
rect 11606 26392 11612 26404
rect 11664 26392 11670 26444
rect 11900 26441 11928 26528
rect 29546 26460 29552 26512
rect 29604 26500 29610 26512
rect 30282 26500 30288 26512
rect 29604 26472 30288 26500
rect 29604 26460 29610 26472
rect 30282 26460 30288 26472
rect 30340 26500 30346 26512
rect 31846 26500 31852 26512
rect 30340 26472 31852 26500
rect 30340 26460 30346 26472
rect 31846 26460 31852 26472
rect 31904 26460 31910 26512
rect 32585 26503 32643 26509
rect 32585 26469 32597 26503
rect 32631 26469 32643 26503
rect 32585 26463 32643 26469
rect 11885 26435 11943 26441
rect 11885 26401 11897 26435
rect 11931 26401 11943 26435
rect 11885 26395 11943 26401
rect 14829 26435 14887 26441
rect 14829 26401 14841 26435
rect 14875 26432 14887 26435
rect 15378 26432 15384 26444
rect 14875 26404 15384 26432
rect 14875 26401 14887 26404
rect 14829 26395 14887 26401
rect 15378 26392 15384 26404
rect 15436 26392 15442 26444
rect 19426 26432 19432 26444
rect 16500 26404 19432 26432
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26364 8447 26367
rect 9125 26367 9183 26373
rect 9125 26364 9137 26367
rect 8435 26336 9137 26364
rect 8435 26333 8447 26336
rect 8389 26327 8447 26333
rect 9125 26333 9137 26336
rect 9171 26333 9183 26367
rect 9125 26327 9183 26333
rect 14090 26324 14096 26376
rect 14148 26364 14154 26376
rect 15105 26367 15163 26373
rect 15105 26364 15117 26367
rect 14148 26336 15117 26364
rect 14148 26324 14154 26336
rect 15105 26333 15117 26336
rect 15151 26333 15163 26367
rect 15105 26327 15163 26333
rect 15930 26324 15936 26376
rect 15988 26364 15994 26376
rect 16261 26367 16319 26373
rect 16261 26364 16273 26367
rect 15988 26336 16273 26364
rect 15988 26324 15994 26336
rect 16261 26333 16273 26336
rect 16307 26333 16319 26367
rect 16390 26364 16396 26376
rect 16351 26336 16396 26364
rect 16261 26327 16319 26333
rect 16390 26324 16396 26336
rect 16448 26324 16454 26376
rect 9306 26296 9312 26308
rect 5684 26268 9168 26296
rect 9267 26268 9312 26296
rect 5684 26256 5690 26268
rect 5442 26228 5448 26240
rect 5184 26200 5448 26228
rect 5442 26188 5448 26200
rect 5500 26188 5506 26240
rect 9140 26228 9168 26268
rect 9306 26256 9312 26268
rect 9364 26256 9370 26308
rect 10965 26299 11023 26305
rect 10965 26296 10977 26299
rect 9416 26268 10977 26296
rect 9416 26228 9444 26268
rect 10965 26265 10977 26268
rect 11011 26296 11023 26299
rect 16500 26296 16528 26404
rect 19426 26392 19432 26404
rect 19484 26432 19490 26444
rect 19705 26435 19763 26441
rect 19705 26432 19717 26435
rect 19484 26404 19717 26432
rect 19484 26392 19490 26404
rect 19705 26401 19717 26404
rect 19751 26401 19763 26435
rect 19705 26395 19763 26401
rect 27985 26435 28043 26441
rect 27985 26401 27997 26435
rect 28031 26432 28043 26435
rect 30926 26432 30932 26444
rect 28031 26404 30932 26432
rect 28031 26401 28043 26404
rect 27985 26395 28043 26401
rect 30926 26392 30932 26404
rect 30984 26392 30990 26444
rect 31386 26432 31392 26444
rect 31347 26404 31392 26432
rect 31386 26392 31392 26404
rect 31444 26392 31450 26444
rect 32214 26392 32220 26444
rect 32272 26392 32278 26444
rect 32600 26432 32628 26463
rect 33134 26460 33140 26512
rect 33192 26500 33198 26512
rect 35253 26503 35311 26509
rect 35253 26500 35265 26503
rect 33192 26472 35265 26500
rect 33192 26460 33198 26472
rect 35253 26469 35265 26472
rect 35299 26469 35311 26503
rect 38010 26500 38016 26512
rect 37971 26472 38016 26500
rect 35253 26463 35311 26469
rect 38010 26460 38016 26472
rect 38068 26460 38074 26512
rect 33318 26432 33324 26444
rect 32600 26404 33324 26432
rect 33318 26392 33324 26404
rect 33376 26392 33382 26444
rect 33502 26432 33508 26444
rect 33463 26404 33508 26432
rect 33502 26392 33508 26404
rect 33560 26392 33566 26444
rect 33689 26435 33747 26441
rect 33689 26401 33701 26435
rect 33735 26432 33747 26435
rect 33778 26432 33784 26444
rect 33735 26404 33784 26432
rect 33735 26401 33747 26404
rect 33689 26395 33747 26401
rect 33778 26392 33784 26404
rect 33836 26432 33842 26444
rect 35897 26435 35955 26441
rect 35897 26432 35909 26435
rect 33836 26404 35909 26432
rect 33836 26392 33842 26404
rect 35897 26401 35909 26404
rect 35943 26432 35955 26435
rect 35986 26432 35992 26444
rect 35943 26404 35992 26432
rect 35943 26401 35955 26404
rect 35897 26395 35955 26401
rect 35986 26392 35992 26404
rect 36044 26392 36050 26444
rect 36630 26392 36636 26444
rect 36688 26432 36694 26444
rect 37090 26432 37096 26444
rect 36688 26404 37096 26432
rect 36688 26392 36694 26404
rect 37090 26392 37096 26404
rect 37148 26392 37154 26444
rect 16577 26367 16635 26373
rect 16577 26333 16589 26367
rect 16623 26364 16635 26367
rect 16666 26364 16672 26376
rect 16623 26336 16672 26364
rect 16623 26333 16635 26336
rect 16577 26327 16635 26333
rect 16666 26324 16672 26336
rect 16724 26364 16730 26376
rect 17037 26367 17095 26373
rect 17037 26364 17049 26367
rect 16724 26336 17049 26364
rect 16724 26324 16730 26336
rect 17037 26333 17049 26336
rect 17083 26333 17095 26367
rect 17037 26327 17095 26333
rect 18693 26367 18751 26373
rect 18693 26333 18705 26367
rect 18739 26364 18751 26367
rect 19245 26367 19303 26373
rect 19245 26364 19257 26367
rect 18739 26336 19257 26364
rect 18739 26333 18751 26336
rect 18693 26327 18751 26333
rect 19245 26333 19257 26336
rect 19291 26333 19303 26367
rect 27706 26364 27712 26376
rect 27667 26336 27712 26364
rect 19245 26327 19303 26333
rect 27706 26324 27712 26336
rect 27764 26324 27770 26376
rect 29546 26364 29552 26376
rect 29507 26336 29552 26364
rect 29546 26324 29552 26336
rect 29604 26324 29610 26376
rect 32030 26364 32036 26376
rect 31991 26336 32036 26364
rect 32030 26324 32036 26336
rect 32088 26324 32094 26376
rect 32232 26364 32260 26392
rect 32309 26367 32367 26373
rect 32309 26364 32321 26367
rect 32232 26336 32321 26364
rect 32309 26333 32321 26336
rect 32355 26333 32367 26367
rect 32309 26327 32367 26333
rect 32401 26367 32459 26373
rect 32401 26333 32413 26367
rect 32447 26364 32459 26367
rect 35618 26364 35624 26376
rect 32447 26336 35624 26364
rect 32447 26333 32459 26336
rect 32401 26327 32459 26333
rect 19426 26296 19432 26308
rect 11011 26268 16528 26296
rect 19387 26268 19432 26296
rect 11011 26265 11023 26268
rect 10965 26259 11023 26265
rect 19426 26256 19432 26268
rect 19484 26256 19490 26308
rect 25682 26256 25688 26308
rect 25740 26296 25746 26308
rect 25961 26299 26019 26305
rect 25961 26296 25973 26299
rect 25740 26268 25973 26296
rect 25740 26256 25746 26268
rect 25961 26265 25973 26268
rect 26007 26265 26019 26299
rect 25961 26259 26019 26265
rect 26697 26299 26755 26305
rect 26697 26265 26709 26299
rect 26743 26296 26755 26299
rect 26878 26296 26884 26308
rect 26743 26268 26884 26296
rect 26743 26265 26755 26268
rect 26697 26259 26755 26265
rect 26878 26256 26884 26268
rect 26936 26256 26942 26308
rect 30006 26256 30012 26308
rect 30064 26296 30070 26308
rect 31205 26299 31263 26305
rect 31205 26296 31217 26299
rect 30064 26268 31217 26296
rect 30064 26256 30070 26268
rect 31205 26265 31217 26268
rect 31251 26265 31263 26299
rect 32214 26296 32220 26308
rect 32175 26268 32220 26296
rect 31205 26259 31263 26265
rect 32214 26256 32220 26268
rect 32272 26256 32278 26308
rect 32324 26296 32352 26327
rect 35618 26324 35624 26336
rect 35676 26324 35682 26376
rect 35713 26367 35771 26373
rect 35713 26333 35725 26367
rect 35759 26364 35771 26367
rect 37366 26364 37372 26376
rect 35759 26336 37372 26364
rect 35759 26333 35771 26336
rect 35713 26327 35771 26333
rect 37366 26324 37372 26336
rect 37424 26324 37430 26376
rect 37642 26324 37648 26376
rect 37700 26364 37706 26376
rect 37829 26367 37887 26373
rect 37829 26364 37841 26367
rect 37700 26336 37841 26364
rect 37700 26324 37706 26336
rect 37829 26333 37841 26336
rect 37875 26333 37887 26367
rect 37829 26327 37887 26333
rect 32674 26296 32680 26308
rect 32324 26268 32680 26296
rect 32674 26256 32680 26268
rect 32732 26256 32738 26308
rect 33410 26296 33416 26308
rect 33371 26268 33416 26296
rect 33410 26256 33416 26268
rect 33468 26256 33474 26308
rect 36909 26299 36967 26305
rect 36909 26296 36921 26299
rect 35912 26268 36921 26296
rect 35912 26240 35940 26268
rect 36909 26265 36921 26268
rect 36955 26265 36967 26299
rect 36909 26259 36967 26265
rect 9140 26200 9444 26228
rect 35621 26231 35679 26237
rect 35621 26197 35633 26231
rect 35667 26228 35679 26231
rect 35894 26228 35900 26240
rect 35667 26200 35900 26228
rect 35667 26197 35679 26200
rect 35621 26191 35679 26197
rect 35894 26188 35900 26200
rect 35952 26188 35958 26240
rect 36078 26188 36084 26240
rect 36136 26228 36142 26240
rect 36817 26231 36875 26237
rect 36817 26228 36829 26231
rect 36136 26200 36829 26228
rect 36136 26188 36142 26200
rect 36817 26197 36829 26200
rect 36863 26197 36875 26231
rect 36817 26191 36875 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 2869 26027 2927 26033
rect 2869 25993 2881 26027
rect 2915 26024 2927 26027
rect 2958 26024 2964 26036
rect 2915 25996 2964 26024
rect 2915 25993 2927 25996
rect 2869 25987 2927 25993
rect 2958 25984 2964 25996
rect 3016 25984 3022 26036
rect 4709 26027 4767 26033
rect 4709 25993 4721 26027
rect 4755 25993 4767 26027
rect 5350 26024 5356 26036
rect 5311 25996 5356 26024
rect 4709 25987 4767 25993
rect 4249 25959 4307 25965
rect 4249 25925 4261 25959
rect 4295 25956 4307 25959
rect 4724 25956 4752 25987
rect 5350 25984 5356 25996
rect 5408 25984 5414 26036
rect 8941 26027 8999 26033
rect 8941 25993 8953 26027
rect 8987 26024 8999 26027
rect 9030 26024 9036 26036
rect 8987 25996 9036 26024
rect 8987 25993 8999 25996
rect 8941 25987 8999 25993
rect 9030 25984 9036 25996
rect 9088 25984 9094 26036
rect 9398 25984 9404 26036
rect 9456 26024 9462 26036
rect 9766 26024 9772 26036
rect 9456 25996 9772 26024
rect 9456 25984 9462 25996
rect 9766 25984 9772 25996
rect 9824 25984 9830 26036
rect 10321 26027 10379 26033
rect 10321 25993 10333 26027
rect 10367 25993 10379 26027
rect 13998 26024 14004 26036
rect 10321 25987 10379 25993
rect 13280 25996 14004 26024
rect 9582 25956 9588 25968
rect 4295 25928 4660 25956
rect 4724 25928 6592 25956
rect 4295 25925 4307 25928
rect 4249 25919 4307 25925
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25848 1458 25900
rect 1578 25848 1584 25900
rect 1636 25888 1642 25900
rect 2409 25891 2467 25897
rect 2409 25888 2421 25891
rect 1636 25860 2421 25888
rect 1636 25848 1642 25860
rect 2409 25857 2421 25860
rect 2455 25857 2467 25891
rect 2409 25851 2467 25857
rect 2685 25891 2743 25897
rect 2685 25857 2697 25891
rect 2731 25857 2743 25891
rect 2685 25851 2743 25857
rect 2700 25820 2728 25851
rect 2866 25848 2872 25900
rect 2924 25888 2930 25900
rect 3053 25891 3111 25897
rect 3053 25888 3065 25891
rect 2924 25860 3065 25888
rect 2924 25848 2930 25860
rect 3053 25857 3065 25860
rect 3099 25857 3111 25891
rect 3053 25851 3111 25857
rect 4154 25848 4160 25900
rect 4212 25888 4218 25900
rect 4525 25891 4583 25897
rect 4525 25888 4537 25891
rect 4212 25860 4537 25888
rect 4212 25848 4218 25860
rect 4525 25857 4537 25860
rect 4571 25857 4583 25891
rect 4632 25888 4660 25928
rect 4798 25888 4804 25900
rect 4632 25860 4804 25888
rect 4525 25851 4583 25857
rect 4798 25848 4804 25860
rect 4856 25848 4862 25900
rect 5166 25888 5172 25900
rect 5127 25860 5172 25888
rect 5166 25848 5172 25860
rect 5224 25848 5230 25900
rect 6564 25897 6592 25928
rect 9140 25928 9588 25956
rect 9140 25897 9168 25928
rect 9582 25916 9588 25928
rect 9640 25956 9646 25968
rect 10042 25956 10048 25968
rect 9640 25928 10048 25956
rect 9640 25916 9646 25928
rect 10042 25916 10048 25928
rect 10100 25956 10106 25968
rect 10100 25928 10180 25956
rect 10100 25916 10106 25928
rect 6549 25891 6607 25897
rect 6549 25857 6561 25891
rect 6595 25857 6607 25891
rect 6549 25851 6607 25857
rect 9125 25891 9183 25897
rect 9125 25857 9137 25891
rect 9171 25857 9183 25891
rect 9398 25888 9404 25900
rect 9359 25860 9404 25888
rect 9125 25851 9183 25857
rect 9398 25848 9404 25860
rect 9456 25848 9462 25900
rect 9861 25891 9919 25897
rect 9861 25857 9873 25891
rect 9907 25888 9919 25891
rect 9950 25888 9956 25900
rect 9907 25860 9956 25888
rect 9907 25857 9919 25860
rect 9861 25851 9919 25857
rect 9950 25848 9956 25860
rect 10008 25848 10014 25900
rect 10152 25897 10180 25928
rect 10137 25891 10195 25897
rect 10137 25857 10149 25891
rect 10183 25857 10195 25891
rect 10336 25888 10364 25987
rect 12526 25956 12532 25968
rect 11716 25928 12532 25956
rect 11716 25897 11744 25928
rect 12526 25916 12532 25928
rect 12584 25916 12590 25968
rect 13280 25900 13308 25996
rect 13998 25984 14004 25996
rect 14056 25984 14062 26036
rect 35989 26027 36047 26033
rect 35989 25993 36001 26027
rect 36035 26024 36047 26027
rect 36170 26024 36176 26036
rect 36035 25996 36176 26024
rect 36035 25993 36047 25996
rect 35989 25987 36047 25993
rect 36170 25984 36176 25996
rect 36228 25984 36234 26036
rect 36354 26024 36360 26036
rect 36315 25996 36360 26024
rect 36354 25984 36360 25996
rect 36412 25984 36418 26036
rect 14090 25956 14096 25968
rect 14051 25928 14096 25956
rect 14090 25916 14096 25928
rect 14148 25916 14154 25968
rect 30926 25956 30932 25968
rect 30887 25928 30932 25956
rect 30926 25916 30932 25928
rect 30984 25916 30990 25968
rect 32030 25916 32036 25968
rect 32088 25956 32094 25968
rect 32585 25959 32643 25965
rect 32585 25956 32597 25959
rect 32088 25928 32597 25956
rect 32088 25916 32094 25928
rect 32585 25925 32597 25928
rect 32631 25925 32643 25959
rect 32585 25919 32643 25925
rect 33410 25916 33416 25968
rect 33468 25956 33474 25968
rect 36449 25959 36507 25965
rect 36449 25956 36461 25959
rect 33468 25928 36461 25956
rect 33468 25916 33474 25928
rect 36449 25925 36461 25928
rect 36495 25925 36507 25959
rect 36449 25919 36507 25925
rect 10965 25891 11023 25897
rect 10965 25888 10977 25891
rect 10336 25860 10977 25888
rect 10137 25851 10195 25857
rect 10965 25857 10977 25860
rect 11011 25857 11023 25891
rect 10965 25851 11023 25857
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 12345 25891 12403 25897
rect 12345 25857 12357 25891
rect 12391 25888 12403 25891
rect 13262 25888 13268 25900
rect 12391 25860 13268 25888
rect 12391 25857 12403 25860
rect 12345 25851 12403 25857
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 22281 25891 22339 25897
rect 22281 25857 22293 25891
rect 22327 25888 22339 25891
rect 24486 25888 24492 25900
rect 22327 25860 24492 25888
rect 22327 25857 22339 25860
rect 22281 25851 22339 25857
rect 24486 25848 24492 25860
rect 24544 25848 24550 25900
rect 27249 25891 27307 25897
rect 27249 25857 27261 25891
rect 27295 25888 27307 25891
rect 28074 25888 28080 25900
rect 27295 25860 28080 25888
rect 27295 25857 27307 25860
rect 27249 25851 27307 25857
rect 28074 25848 28080 25860
rect 28132 25848 28138 25900
rect 32122 25848 32128 25900
rect 32180 25888 32186 25900
rect 32401 25891 32459 25897
rect 32401 25888 32413 25891
rect 32180 25860 32413 25888
rect 32180 25848 32186 25860
rect 32401 25857 32413 25860
rect 32447 25857 32459 25891
rect 32674 25888 32680 25900
rect 32635 25860 32680 25888
rect 32401 25851 32459 25857
rect 32674 25848 32680 25860
rect 32732 25848 32738 25900
rect 32769 25891 32827 25897
rect 32769 25857 32781 25891
rect 32815 25888 32827 25891
rect 33226 25888 33232 25900
rect 32815 25860 33232 25888
rect 32815 25857 32827 25860
rect 32769 25851 32827 25857
rect 33226 25848 33232 25860
rect 33284 25848 33290 25900
rect 1596 25792 2728 25820
rect 4433 25823 4491 25829
rect 1596 25761 1624 25792
rect 4433 25789 4445 25823
rect 4479 25820 4491 25823
rect 4614 25820 4620 25832
rect 4479 25792 4620 25820
rect 4479 25789 4491 25792
rect 4433 25783 4491 25789
rect 4614 25780 4620 25792
rect 4672 25780 4678 25832
rect 4982 25780 4988 25832
rect 5040 25820 5046 25832
rect 5350 25820 5356 25832
rect 5040 25792 5356 25820
rect 5040 25780 5046 25792
rect 5350 25780 5356 25792
rect 5408 25780 5414 25832
rect 9214 25820 9220 25832
rect 9175 25792 9220 25820
rect 9214 25780 9220 25792
rect 9272 25780 9278 25832
rect 10045 25823 10103 25829
rect 10045 25789 10057 25823
rect 10091 25820 10103 25823
rect 10226 25820 10232 25832
rect 10091 25792 10232 25820
rect 10091 25789 10103 25792
rect 10045 25783 10103 25789
rect 10226 25780 10232 25792
rect 10284 25780 10290 25832
rect 13449 25823 13507 25829
rect 13449 25789 13461 25823
rect 13495 25820 13507 25823
rect 13909 25823 13967 25829
rect 13909 25820 13921 25823
rect 13495 25792 13921 25820
rect 13495 25789 13507 25792
rect 13449 25783 13507 25789
rect 13909 25789 13921 25792
rect 13955 25789 13967 25823
rect 15286 25820 15292 25832
rect 15247 25792 15292 25820
rect 13909 25783 13967 25789
rect 15286 25780 15292 25792
rect 15344 25780 15350 25832
rect 25866 25780 25872 25832
rect 25924 25820 25930 25832
rect 26973 25823 27031 25829
rect 26973 25820 26985 25823
rect 25924 25792 26985 25820
rect 25924 25780 25930 25792
rect 26973 25789 26985 25792
rect 27019 25789 27031 25823
rect 29270 25820 29276 25832
rect 29231 25792 29276 25820
rect 26973 25783 27031 25789
rect 29270 25780 29276 25792
rect 29328 25780 29334 25832
rect 31113 25823 31171 25829
rect 31113 25789 31125 25823
rect 31159 25820 31171 25823
rect 33410 25820 33416 25832
rect 31159 25792 33416 25820
rect 31159 25789 31171 25792
rect 31113 25783 31171 25789
rect 33410 25780 33416 25792
rect 33468 25780 33474 25832
rect 36630 25820 36636 25832
rect 36591 25792 36636 25820
rect 36630 25780 36636 25792
rect 36688 25780 36694 25832
rect 1581 25755 1639 25761
rect 1581 25721 1593 25755
rect 1627 25721 1639 25755
rect 5074 25752 5080 25764
rect 1581 25715 1639 25721
rect 4540 25724 5080 25752
rect 2590 25684 2596 25696
rect 2551 25656 2596 25684
rect 2590 25644 2596 25656
rect 2648 25644 2654 25696
rect 4540 25693 4568 25724
rect 5074 25712 5080 25724
rect 5132 25712 5138 25764
rect 9306 25712 9312 25764
rect 9364 25752 9370 25764
rect 10781 25755 10839 25761
rect 10781 25752 10793 25755
rect 9364 25724 10793 25752
rect 9364 25712 9370 25724
rect 10781 25721 10793 25724
rect 10827 25721 10839 25755
rect 22462 25752 22468 25764
rect 10781 25715 10839 25721
rect 10888 25724 11744 25752
rect 22423 25724 22468 25752
rect 4525 25687 4583 25693
rect 4525 25653 4537 25687
rect 4571 25653 4583 25687
rect 4525 25647 4583 25653
rect 4982 25644 4988 25696
rect 5040 25684 5046 25696
rect 6365 25687 6423 25693
rect 6365 25684 6377 25687
rect 5040 25656 6377 25684
rect 5040 25644 5046 25656
rect 6365 25653 6377 25656
rect 6411 25653 6423 25687
rect 6365 25647 6423 25653
rect 9401 25687 9459 25693
rect 9401 25653 9413 25687
rect 9447 25684 9459 25687
rect 9766 25684 9772 25696
rect 9447 25656 9772 25684
rect 9447 25653 9459 25656
rect 9401 25647 9459 25653
rect 9766 25644 9772 25656
rect 9824 25684 9830 25696
rect 10137 25687 10195 25693
rect 10137 25684 10149 25687
rect 9824 25656 10149 25684
rect 9824 25644 9830 25656
rect 10137 25653 10149 25656
rect 10183 25684 10195 25687
rect 10318 25684 10324 25696
rect 10183 25656 10324 25684
rect 10183 25653 10195 25656
rect 10137 25647 10195 25653
rect 10318 25644 10324 25656
rect 10376 25684 10382 25696
rect 10888 25684 10916 25724
rect 11716 25696 11744 25724
rect 22462 25712 22468 25724
rect 22520 25712 22526 25764
rect 29288 25752 29316 25780
rect 31938 25752 31944 25764
rect 29288 25724 31944 25752
rect 31938 25712 31944 25724
rect 31996 25712 32002 25764
rect 32122 25712 32128 25764
rect 32180 25752 32186 25764
rect 33505 25755 33563 25761
rect 33505 25752 33517 25755
rect 32180 25724 33517 25752
rect 32180 25712 32186 25724
rect 33505 25721 33517 25724
rect 33551 25721 33563 25755
rect 33505 25715 33563 25721
rect 10376 25656 10916 25684
rect 10376 25644 10382 25656
rect 10962 25644 10968 25696
rect 11020 25684 11026 25696
rect 11517 25687 11575 25693
rect 11517 25684 11529 25687
rect 11020 25656 11529 25684
rect 11020 25644 11026 25656
rect 11517 25653 11529 25656
rect 11563 25653 11575 25687
rect 11517 25647 11575 25653
rect 11698 25644 11704 25696
rect 11756 25684 11762 25696
rect 12161 25687 12219 25693
rect 12161 25684 12173 25687
rect 11756 25656 12173 25684
rect 11756 25644 11762 25656
rect 12161 25653 12173 25656
rect 12207 25653 12219 25687
rect 12161 25647 12219 25653
rect 23014 25644 23020 25696
rect 23072 25684 23078 25696
rect 23109 25687 23167 25693
rect 23109 25684 23121 25687
rect 23072 25656 23121 25684
rect 23072 25644 23078 25656
rect 23109 25653 23121 25656
rect 23155 25653 23167 25687
rect 23109 25647 23167 25653
rect 25317 25687 25375 25693
rect 25317 25653 25329 25687
rect 25363 25684 25375 25687
rect 25406 25684 25412 25696
rect 25363 25656 25412 25684
rect 25363 25653 25375 25656
rect 25317 25647 25375 25653
rect 25406 25644 25412 25656
rect 25464 25684 25470 25696
rect 25777 25687 25835 25693
rect 25777 25684 25789 25687
rect 25464 25656 25789 25684
rect 25464 25644 25470 25656
rect 25777 25653 25789 25656
rect 25823 25653 25835 25687
rect 25777 25647 25835 25653
rect 26050 25644 26056 25696
rect 26108 25684 26114 25696
rect 26329 25687 26387 25693
rect 26329 25684 26341 25687
rect 26108 25656 26341 25684
rect 26108 25644 26114 25656
rect 26329 25653 26341 25656
rect 26375 25653 26387 25687
rect 32950 25684 32956 25696
rect 32911 25656 32956 25684
rect 26329 25647 26387 25653
rect 32950 25644 32956 25656
rect 33008 25644 33014 25696
rect 35529 25687 35587 25693
rect 35529 25653 35541 25687
rect 35575 25684 35587 25687
rect 35894 25684 35900 25696
rect 35575 25656 35900 25684
rect 35575 25653 35587 25656
rect 35529 25647 35587 25653
rect 35894 25644 35900 25656
rect 35952 25684 35958 25696
rect 36262 25684 36268 25696
rect 35952 25656 36268 25684
rect 35952 25644 35958 25656
rect 36262 25644 36268 25656
rect 36320 25644 36326 25696
rect 37642 25684 37648 25696
rect 37603 25656 37648 25684
rect 37642 25644 37648 25656
rect 37700 25644 37706 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 4157 25483 4215 25489
rect 4157 25449 4169 25483
rect 4203 25449 4215 25483
rect 4157 25443 4215 25449
rect 4341 25483 4399 25489
rect 4341 25449 4353 25483
rect 4387 25480 4399 25483
rect 5166 25480 5172 25492
rect 4387 25452 5172 25480
rect 4387 25449 4399 25452
rect 4341 25443 4399 25449
rect 1394 25412 1400 25424
rect 1355 25384 1400 25412
rect 1394 25372 1400 25384
rect 1452 25372 1458 25424
rect 4172 25412 4200 25443
rect 5166 25440 5172 25452
rect 5224 25440 5230 25492
rect 10410 25440 10416 25492
rect 10468 25480 10474 25492
rect 11241 25483 11299 25489
rect 11241 25480 11253 25483
rect 10468 25452 11253 25480
rect 10468 25440 10474 25452
rect 11241 25449 11253 25452
rect 11287 25449 11299 25483
rect 11698 25480 11704 25492
rect 11659 25452 11704 25480
rect 11241 25443 11299 25449
rect 11698 25440 11704 25452
rect 11756 25440 11762 25492
rect 19426 25480 19432 25492
rect 19387 25452 19432 25480
rect 19426 25440 19432 25452
rect 19484 25440 19490 25492
rect 21818 25480 21824 25492
rect 21779 25452 21824 25480
rect 21818 25440 21824 25452
rect 21876 25440 21882 25492
rect 25685 25483 25743 25489
rect 25685 25449 25697 25483
rect 25731 25449 25743 25483
rect 25866 25480 25872 25492
rect 25827 25452 25872 25480
rect 25685 25443 25743 25449
rect 5074 25412 5080 25424
rect 4172 25384 5080 25412
rect 5074 25372 5080 25384
rect 5132 25372 5138 25424
rect 10226 25372 10232 25424
rect 10284 25412 10290 25424
rect 25700 25412 25728 25443
rect 25866 25440 25872 25452
rect 25924 25440 25930 25492
rect 26329 25483 26387 25489
rect 26329 25449 26341 25483
rect 26375 25449 26387 25483
rect 26329 25443 26387 25449
rect 26142 25412 26148 25424
rect 10284 25384 11560 25412
rect 25700 25384 26148 25412
rect 10284 25372 10290 25384
rect 4065 25347 4123 25353
rect 4065 25313 4077 25347
rect 4111 25344 4123 25347
rect 4614 25344 4620 25356
rect 4111 25316 4620 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 4614 25304 4620 25316
rect 4672 25304 4678 25356
rect 4706 25304 4712 25356
rect 4764 25344 4770 25356
rect 4801 25347 4859 25353
rect 4801 25344 4813 25347
rect 4764 25316 4813 25344
rect 4764 25304 4770 25316
rect 4801 25313 4813 25316
rect 4847 25313 4859 25347
rect 4982 25344 4988 25356
rect 4943 25316 4988 25344
rect 4801 25307 4859 25313
rect 4982 25304 4988 25316
rect 5040 25304 5046 25356
rect 5534 25344 5540 25356
rect 5495 25316 5540 25344
rect 5534 25304 5540 25316
rect 5592 25304 5598 25356
rect 9766 25344 9772 25356
rect 9727 25316 9772 25344
rect 9766 25304 9772 25316
rect 9824 25304 9830 25356
rect 10042 25304 10048 25356
rect 10100 25344 10106 25356
rect 10962 25344 10968 25356
rect 10100 25316 10968 25344
rect 10100 25304 10106 25316
rect 10962 25304 10968 25316
rect 11020 25344 11026 25356
rect 11532 25353 11560 25384
rect 26142 25372 26148 25384
rect 26200 25412 26206 25424
rect 26344 25412 26372 25443
rect 26694 25440 26700 25492
rect 26752 25480 26758 25492
rect 26789 25483 26847 25489
rect 26789 25480 26801 25483
rect 26752 25452 26801 25480
rect 26752 25440 26758 25452
rect 26789 25449 26801 25452
rect 26835 25449 26847 25483
rect 26789 25443 26847 25449
rect 32214 25440 32220 25492
rect 32272 25480 32278 25492
rect 32401 25483 32459 25489
rect 32401 25480 32413 25483
rect 32272 25452 32413 25480
rect 32272 25440 32278 25452
rect 32401 25449 32413 25452
rect 32447 25449 32459 25483
rect 32401 25443 32459 25449
rect 26200 25384 26372 25412
rect 26200 25372 26206 25384
rect 11517 25347 11575 25353
rect 11020 25316 11468 25344
rect 11020 25304 11026 25316
rect 2590 25276 2596 25288
rect 2551 25248 2596 25276
rect 2590 25236 2596 25248
rect 2648 25236 2654 25288
rect 3234 25276 3240 25288
rect 3195 25248 3240 25276
rect 3234 25236 3240 25248
rect 3292 25236 3298 25288
rect 4154 25276 4160 25288
rect 4067 25248 4160 25276
rect 4154 25236 4160 25248
rect 4212 25276 4218 25288
rect 11440 25285 11468 25316
rect 11517 25313 11529 25347
rect 11563 25313 11575 25347
rect 21634 25344 21640 25356
rect 21595 25316 21640 25344
rect 11517 25307 11575 25313
rect 21634 25304 21640 25316
rect 21692 25304 21698 25356
rect 24946 25304 24952 25356
rect 25004 25344 25010 25356
rect 25501 25347 25559 25353
rect 25501 25344 25513 25347
rect 25004 25316 25513 25344
rect 25004 25304 25010 25316
rect 25501 25313 25513 25316
rect 25547 25344 25559 25347
rect 26050 25344 26056 25356
rect 25547 25316 26056 25344
rect 25547 25313 25559 25316
rect 25501 25307 25559 25313
rect 26050 25304 26056 25316
rect 26108 25344 26114 25356
rect 26421 25347 26479 25353
rect 26421 25344 26433 25347
rect 26108 25316 26433 25344
rect 26108 25304 26114 25316
rect 26421 25313 26433 25316
rect 26467 25313 26479 25347
rect 26421 25307 26479 25313
rect 27985 25347 28043 25353
rect 27985 25313 27997 25347
rect 28031 25344 28043 25347
rect 30006 25344 30012 25356
rect 28031 25316 30012 25344
rect 28031 25313 28043 25316
rect 27985 25307 28043 25313
rect 30006 25304 30012 25316
rect 30064 25304 30070 25356
rect 30834 25304 30840 25356
rect 30892 25344 30898 25356
rect 31757 25347 31815 25353
rect 31757 25344 31769 25347
rect 30892 25316 31769 25344
rect 30892 25304 30898 25316
rect 31757 25313 31769 25316
rect 31803 25313 31815 25347
rect 33134 25344 33140 25356
rect 31757 25307 31815 25313
rect 33060 25316 33140 25344
rect 8389 25279 8447 25285
rect 4212 25248 4844 25276
rect 4212 25236 4218 25248
rect 3881 25211 3939 25217
rect 3881 25177 3893 25211
rect 3927 25208 3939 25211
rect 4706 25208 4712 25220
rect 3927 25180 4712 25208
rect 3927 25177 3939 25180
rect 3881 25171 3939 25177
rect 4706 25168 4712 25180
rect 4764 25168 4770 25220
rect 4816 25152 4844 25248
rect 8389 25245 8401 25279
rect 8435 25276 8447 25279
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8435 25248 8953 25276
rect 8435 25245 8447 25248
rect 8389 25239 8447 25245
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 11425 25279 11483 25285
rect 11425 25245 11437 25279
rect 11471 25245 11483 25279
rect 19242 25276 19248 25288
rect 19203 25248 19248 25276
rect 11425 25239 11483 25245
rect 19242 25236 19248 25248
rect 19300 25236 19306 25288
rect 21358 25236 21364 25288
rect 21416 25276 21422 25288
rect 21545 25279 21603 25285
rect 21545 25276 21557 25279
rect 21416 25248 21557 25276
rect 21416 25236 21422 25248
rect 21545 25245 21557 25248
rect 21591 25245 21603 25279
rect 21545 25239 21603 25245
rect 21821 25279 21879 25285
rect 21821 25245 21833 25279
rect 21867 25276 21879 25279
rect 21910 25276 21916 25288
rect 21867 25248 21916 25276
rect 21867 25245 21879 25248
rect 21821 25239 21879 25245
rect 9122 25208 9128 25220
rect 9083 25180 9128 25208
rect 9122 25168 9128 25180
rect 9180 25168 9186 25220
rect 9950 25168 9956 25220
rect 10008 25208 10014 25220
rect 11701 25211 11759 25217
rect 11701 25208 11713 25211
rect 10008 25180 11713 25208
rect 10008 25168 10014 25180
rect 11701 25177 11713 25180
rect 11747 25177 11759 25211
rect 21560 25208 21588 25239
rect 21910 25236 21916 25248
rect 21968 25236 21974 25288
rect 25682 25276 25688 25288
rect 25643 25248 25688 25276
rect 25682 25236 25688 25248
rect 25740 25276 25746 25288
rect 26605 25279 26663 25285
rect 26605 25276 26617 25279
rect 25740 25248 26617 25276
rect 25740 25236 25746 25248
rect 26605 25245 26617 25248
rect 26651 25245 26663 25279
rect 26605 25239 26663 25245
rect 26970 25236 26976 25288
rect 27028 25276 27034 25288
rect 27709 25279 27767 25285
rect 27709 25276 27721 25279
rect 27028 25248 27721 25276
rect 27028 25236 27034 25248
rect 27709 25245 27721 25248
rect 27755 25245 27767 25279
rect 30374 25276 30380 25288
rect 30287 25248 30380 25276
rect 27709 25239 27767 25245
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 30653 25279 30711 25285
rect 30653 25245 30665 25279
rect 30699 25276 30711 25279
rect 30926 25276 30932 25288
rect 30699 25248 30932 25276
rect 30699 25245 30711 25248
rect 30653 25239 30711 25245
rect 30926 25236 30932 25248
rect 30984 25236 30990 25288
rect 32033 25279 32091 25285
rect 32033 25276 32045 25279
rect 31220 25248 32045 25276
rect 21726 25208 21732 25220
rect 21560 25180 21732 25208
rect 11701 25171 11759 25177
rect 21726 25168 21732 25180
rect 21784 25208 21790 25220
rect 22557 25211 22615 25217
rect 22557 25208 22569 25211
rect 21784 25180 22569 25208
rect 21784 25168 21790 25180
rect 22557 25177 22569 25180
rect 22603 25177 22615 25211
rect 22557 25171 22615 25177
rect 22741 25211 22799 25217
rect 22741 25177 22753 25211
rect 22787 25208 22799 25211
rect 22830 25208 22836 25220
rect 22787 25180 22836 25208
rect 22787 25177 22799 25180
rect 22741 25171 22799 25177
rect 22830 25168 22836 25180
rect 22888 25208 22894 25220
rect 25406 25208 25412 25220
rect 22888 25180 25412 25208
rect 22888 25168 22894 25180
rect 25406 25168 25412 25180
rect 25464 25168 25470 25220
rect 26329 25211 26387 25217
rect 26329 25208 26341 25211
rect 26206 25180 26341 25208
rect 2774 25100 2780 25152
rect 2832 25140 2838 25152
rect 3053 25143 3111 25149
rect 3053 25140 3065 25143
rect 2832 25112 3065 25140
rect 2832 25100 2838 25112
rect 3053 25109 3065 25112
rect 3099 25109 3111 25143
rect 3053 25103 3111 25109
rect 4798 25100 4804 25152
rect 4856 25100 4862 25152
rect 22002 25140 22008 25152
rect 21963 25112 22008 25140
rect 22002 25100 22008 25112
rect 22060 25100 22066 25152
rect 24946 25140 24952 25152
rect 24907 25112 24952 25140
rect 24946 25100 24952 25112
rect 25004 25100 25010 25152
rect 25774 25100 25780 25152
rect 25832 25140 25838 25152
rect 26050 25140 26056 25152
rect 25832 25112 26056 25140
rect 25832 25100 25838 25112
rect 26050 25100 26056 25112
rect 26108 25140 26114 25152
rect 26206 25140 26234 25180
rect 26329 25177 26341 25180
rect 26375 25177 26387 25211
rect 30392 25208 30420 25236
rect 31110 25208 31116 25220
rect 30392 25180 31116 25208
rect 26329 25171 26387 25177
rect 31110 25168 31116 25180
rect 31168 25168 31174 25220
rect 26108 25112 26234 25140
rect 26108 25100 26114 25112
rect 29546 25100 29552 25152
rect 29604 25140 29610 25152
rect 29825 25143 29883 25149
rect 29825 25140 29837 25143
rect 29604 25112 29837 25140
rect 29604 25100 29610 25112
rect 29825 25109 29837 25112
rect 29871 25140 29883 25143
rect 31220 25140 31248 25248
rect 32033 25245 32045 25248
rect 32079 25276 32091 25279
rect 32122 25276 32128 25288
rect 32079 25248 32128 25276
rect 32079 25245 32091 25248
rect 32033 25239 32091 25245
rect 32122 25236 32128 25248
rect 32180 25236 32186 25288
rect 32306 25236 32312 25288
rect 32364 25276 32370 25288
rect 32674 25276 32680 25288
rect 32364 25248 32680 25276
rect 32364 25236 32370 25248
rect 32674 25236 32680 25248
rect 32732 25276 32738 25288
rect 33060 25285 33088 25316
rect 33134 25304 33140 25316
rect 33192 25304 33198 25356
rect 32861 25279 32919 25285
rect 32861 25276 32873 25279
rect 32732 25248 32873 25276
rect 32732 25236 32738 25248
rect 32861 25245 32873 25248
rect 32907 25245 32919 25279
rect 32861 25239 32919 25245
rect 33045 25279 33103 25285
rect 33045 25245 33057 25279
rect 33091 25245 33103 25279
rect 33226 25276 33232 25288
rect 33187 25248 33232 25276
rect 33045 25239 33103 25245
rect 33226 25236 33232 25248
rect 33284 25236 33290 25288
rect 33137 25211 33195 25217
rect 33137 25208 33149 25211
rect 31956 25180 33149 25208
rect 29871 25112 31248 25140
rect 29871 25109 29883 25112
rect 29825 25103 29883 25109
rect 31846 25100 31852 25152
rect 31904 25140 31910 25152
rect 31956 25149 31984 25180
rect 33137 25177 33149 25180
rect 33183 25208 33195 25211
rect 33873 25211 33931 25217
rect 33873 25208 33885 25211
rect 33183 25180 33885 25208
rect 33183 25177 33195 25180
rect 33137 25171 33195 25177
rect 33873 25177 33885 25180
rect 33919 25177 33931 25211
rect 33873 25171 33931 25177
rect 31941 25143 31999 25149
rect 31941 25140 31953 25143
rect 31904 25112 31953 25140
rect 31904 25100 31910 25112
rect 31941 25109 31953 25112
rect 31987 25109 31999 25143
rect 31941 25103 31999 25109
rect 33413 25143 33471 25149
rect 33413 25109 33425 25143
rect 33459 25140 33471 25143
rect 33502 25140 33508 25152
rect 33459 25112 33508 25140
rect 33459 25109 33471 25112
rect 33413 25103 33471 25109
rect 33502 25100 33508 25112
rect 33560 25100 33566 25152
rect 36173 25143 36231 25149
rect 36173 25109 36185 25143
rect 36219 25140 36231 25143
rect 36262 25140 36268 25152
rect 36219 25112 36268 25140
rect 36219 25109 36231 25112
rect 36173 25103 36231 25109
rect 36262 25100 36268 25112
rect 36320 25100 36326 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 9122 24896 9128 24948
rect 9180 24936 9186 24948
rect 9217 24939 9275 24945
rect 9217 24936 9229 24939
rect 9180 24908 9229 24936
rect 9180 24896 9186 24908
rect 9217 24905 9229 24908
rect 9263 24905 9275 24939
rect 26329 24939 26387 24945
rect 26329 24936 26341 24939
rect 9217 24899 9275 24905
rect 25516 24908 26341 24936
rect 2774 24868 2780 24880
rect 2735 24840 2780 24868
rect 2774 24828 2780 24840
rect 2832 24828 2838 24880
rect 9766 24828 9772 24880
rect 9824 24868 9830 24880
rect 9824 24840 14044 24868
rect 9824 24828 9830 24840
rect 2590 24800 2596 24812
rect 2551 24772 2596 24800
rect 2590 24760 2596 24772
rect 2648 24760 2654 24812
rect 5074 24760 5080 24812
rect 5132 24800 5138 24812
rect 5537 24803 5595 24809
rect 5537 24800 5549 24803
rect 5132 24772 5549 24800
rect 5132 24760 5138 24772
rect 5537 24769 5549 24772
rect 5583 24769 5595 24803
rect 5537 24763 5595 24769
rect 9401 24803 9459 24809
rect 9401 24769 9413 24803
rect 9447 24800 9459 24803
rect 10042 24800 10048 24812
rect 9447 24772 9904 24800
rect 10003 24772 10048 24800
rect 9447 24769 9459 24772
rect 9401 24763 9459 24769
rect 3050 24732 3056 24744
rect 3011 24704 3056 24732
rect 3050 24692 3056 24704
rect 3108 24692 3114 24744
rect 5813 24735 5871 24741
rect 5813 24701 5825 24735
rect 5859 24701 5871 24735
rect 5813 24695 5871 24701
rect 5828 24608 5856 24695
rect 9876 24673 9904 24772
rect 10042 24760 10048 24772
rect 10100 24760 10106 24812
rect 10134 24760 10140 24812
rect 10192 24800 10198 24812
rect 10321 24803 10379 24809
rect 10321 24800 10333 24803
rect 10192 24772 10333 24800
rect 10192 24760 10198 24772
rect 10321 24769 10333 24772
rect 10367 24769 10379 24803
rect 10321 24763 10379 24769
rect 10226 24732 10232 24744
rect 10187 24704 10232 24732
rect 10226 24692 10232 24704
rect 10284 24692 10290 24744
rect 14016 24732 14044 24840
rect 21726 24828 21732 24880
rect 21784 24868 21790 24880
rect 21821 24871 21879 24877
rect 21821 24868 21833 24871
rect 21784 24840 21833 24868
rect 21784 24828 21790 24840
rect 21821 24837 21833 24840
rect 21867 24837 21879 24871
rect 21821 24831 21879 24837
rect 21910 24828 21916 24880
rect 21968 24828 21974 24880
rect 25406 24868 25412 24880
rect 25367 24840 25412 24868
rect 25406 24828 25412 24840
rect 25464 24828 25470 24880
rect 16666 24760 16672 24812
rect 16724 24800 16730 24812
rect 17221 24803 17279 24809
rect 17221 24800 17233 24803
rect 16724 24772 17233 24800
rect 16724 24760 16730 24772
rect 17221 24769 17233 24772
rect 17267 24800 17279 24803
rect 17773 24803 17831 24809
rect 17773 24800 17785 24803
rect 17267 24772 17785 24800
rect 17267 24769 17279 24772
rect 17221 24763 17279 24769
rect 17773 24769 17785 24772
rect 17819 24800 17831 24803
rect 18325 24803 18383 24809
rect 18325 24800 18337 24803
rect 17819 24772 18337 24800
rect 17819 24769 17831 24772
rect 17773 24763 17831 24769
rect 18325 24769 18337 24772
rect 18371 24769 18383 24803
rect 18325 24763 18383 24769
rect 20162 24760 20168 24812
rect 20220 24800 20226 24812
rect 20625 24803 20683 24809
rect 20625 24800 20637 24803
rect 20220 24772 20637 24800
rect 20220 24760 20226 24772
rect 20625 24769 20637 24772
rect 20671 24800 20683 24803
rect 21928 24800 21956 24828
rect 22097 24803 22155 24809
rect 22097 24800 22109 24803
rect 20671 24772 22109 24800
rect 20671 24769 20683 24772
rect 20625 24763 20683 24769
rect 22097 24769 22109 24772
rect 22143 24769 22155 24803
rect 23014 24800 23020 24812
rect 22975 24772 23020 24800
rect 22097 24763 22155 24769
rect 23014 24760 23020 24772
rect 23072 24760 23078 24812
rect 15105 24735 15163 24741
rect 15105 24732 15117 24735
rect 14016 24704 15117 24732
rect 15105 24701 15117 24704
rect 15151 24732 15163 24735
rect 15286 24732 15292 24744
rect 15151 24704 15292 24732
rect 15151 24701 15163 24704
rect 15105 24695 15163 24701
rect 15286 24692 15292 24704
rect 15344 24692 15350 24744
rect 15654 24732 15660 24744
rect 15615 24704 15660 24732
rect 15654 24692 15660 24704
rect 15712 24692 15718 24744
rect 15838 24732 15844 24744
rect 15799 24704 15844 24732
rect 15838 24692 15844 24704
rect 15896 24692 15902 24744
rect 20346 24732 20352 24744
rect 20307 24704 20352 24732
rect 20346 24692 20352 24704
rect 20404 24692 20410 24744
rect 21634 24692 21640 24744
rect 21692 24732 21698 24744
rect 21913 24735 21971 24741
rect 21913 24732 21925 24735
rect 21692 24704 21925 24732
rect 21692 24692 21698 24704
rect 21913 24701 21925 24704
rect 21959 24701 21971 24735
rect 21913 24695 21971 24701
rect 22922 24692 22928 24744
rect 22980 24732 22986 24744
rect 23201 24735 23259 24741
rect 23201 24732 23213 24735
rect 22980 24704 23213 24732
rect 22980 24692 22986 24704
rect 23201 24701 23213 24704
rect 23247 24701 23259 24735
rect 23474 24732 23480 24744
rect 23435 24704 23480 24732
rect 23201 24695 23259 24701
rect 23474 24692 23480 24704
rect 23532 24692 23538 24744
rect 24946 24692 24952 24744
rect 25004 24732 25010 24744
rect 25516 24741 25544 24908
rect 26329 24905 26341 24908
rect 26375 24905 26387 24939
rect 26329 24899 26387 24905
rect 25700 24840 27292 24868
rect 25700 24812 25728 24840
rect 25682 24800 25688 24812
rect 25643 24772 25688 24800
rect 25682 24760 25688 24772
rect 25740 24760 25746 24812
rect 26050 24760 26056 24812
rect 26108 24800 26114 24812
rect 27264 24809 27292 24840
rect 29914 24828 29920 24880
rect 29972 24868 29978 24880
rect 29972 24840 30144 24868
rect 29972 24828 29978 24840
rect 30116 24809 30144 24840
rect 26973 24803 27031 24809
rect 26973 24800 26985 24803
rect 26108 24772 26985 24800
rect 26108 24760 26114 24772
rect 26973 24769 26985 24772
rect 27019 24769 27031 24803
rect 26973 24763 27031 24769
rect 27249 24803 27307 24809
rect 27249 24769 27261 24803
rect 27295 24769 27307 24803
rect 27249 24763 27307 24769
rect 30101 24803 30159 24809
rect 30101 24769 30113 24803
rect 30147 24769 30159 24803
rect 30650 24800 30656 24812
rect 30611 24772 30656 24800
rect 30101 24763 30159 24769
rect 30650 24760 30656 24772
rect 30708 24760 30714 24812
rect 30926 24760 30932 24812
rect 30984 24800 30990 24812
rect 33594 24800 33600 24812
rect 30984 24772 33600 24800
rect 30984 24760 30990 24772
rect 33594 24760 33600 24772
rect 33652 24760 33658 24812
rect 25501 24735 25559 24741
rect 25501 24732 25513 24735
rect 25004 24704 25513 24732
rect 25004 24692 25010 24704
rect 25501 24701 25513 24704
rect 25547 24701 25559 24735
rect 25501 24695 25559 24701
rect 25590 24692 25596 24744
rect 25648 24732 25654 24744
rect 26142 24732 26148 24744
rect 25648 24704 26148 24732
rect 25648 24692 25654 24704
rect 26142 24692 26148 24704
rect 26200 24732 26206 24744
rect 26200 24704 27016 24732
rect 26200 24692 26206 24704
rect 9861 24667 9919 24673
rect 9861 24633 9873 24667
rect 9907 24633 9919 24667
rect 22281 24667 22339 24673
rect 9861 24627 9919 24633
rect 9968 24636 22232 24664
rect 3418 24556 3424 24608
rect 3476 24596 3482 24608
rect 4890 24596 4896 24608
rect 3476 24568 4896 24596
rect 3476 24556 3482 24568
rect 4890 24556 4896 24568
rect 4948 24556 4954 24608
rect 5810 24556 5816 24608
rect 5868 24596 5874 24608
rect 6365 24599 6423 24605
rect 6365 24596 6377 24599
rect 5868 24568 6377 24596
rect 5868 24556 5874 24568
rect 6365 24565 6377 24568
rect 6411 24596 6423 24599
rect 9968 24596 9996 24636
rect 10318 24596 10324 24608
rect 6411 24568 9996 24596
rect 10279 24568 10324 24596
rect 6411 24565 6423 24568
rect 6365 24559 6423 24565
rect 10318 24556 10324 24568
rect 10376 24556 10382 24608
rect 21818 24596 21824 24608
rect 21779 24568 21824 24596
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 22204 24596 22232 24636
rect 22281 24633 22293 24667
rect 22327 24664 22339 24667
rect 26602 24664 26608 24676
rect 22327 24636 26608 24664
rect 22327 24633 22339 24636
rect 22281 24627 22339 24633
rect 26602 24624 26608 24636
rect 26660 24624 26666 24676
rect 23658 24596 23664 24608
rect 22204 24568 23664 24596
rect 23658 24556 23664 24568
rect 23716 24556 23722 24608
rect 25406 24596 25412 24608
rect 25367 24568 25412 24596
rect 25406 24556 25412 24568
rect 25464 24556 25470 24608
rect 25869 24599 25927 24605
rect 25869 24565 25881 24599
rect 25915 24596 25927 24599
rect 26234 24596 26240 24608
rect 25915 24568 26240 24596
rect 25915 24565 25927 24568
rect 25869 24559 25927 24565
rect 26234 24556 26240 24568
rect 26292 24556 26298 24608
rect 26988 24605 27016 24704
rect 27062 24692 27068 24744
rect 27120 24732 27126 24744
rect 27120 24704 27165 24732
rect 27120 24692 27126 24704
rect 28994 24692 29000 24744
rect 29052 24732 29058 24744
rect 29638 24732 29644 24744
rect 29052 24704 29644 24732
rect 29052 24692 29058 24704
rect 29638 24692 29644 24704
rect 29696 24692 29702 24744
rect 29914 24732 29920 24744
rect 29875 24704 29920 24732
rect 29914 24692 29920 24704
rect 29972 24692 29978 24744
rect 27433 24667 27491 24673
rect 27433 24633 27445 24667
rect 27479 24664 27491 24667
rect 27706 24664 27712 24676
rect 27479 24636 27712 24664
rect 27479 24633 27491 24636
rect 27433 24627 27491 24633
rect 27706 24624 27712 24636
rect 27764 24624 27770 24676
rect 31662 24624 31668 24676
rect 31720 24664 31726 24676
rect 33137 24667 33195 24673
rect 33137 24664 33149 24667
rect 31720 24636 33149 24664
rect 31720 24624 31726 24636
rect 33137 24633 33149 24636
rect 33183 24664 33195 24667
rect 33226 24664 33232 24676
rect 33183 24636 33232 24664
rect 33183 24633 33195 24636
rect 33137 24627 33195 24633
rect 33226 24624 33232 24636
rect 33284 24624 33290 24676
rect 26973 24599 27031 24605
rect 26973 24565 26985 24599
rect 27019 24565 27031 24599
rect 26973 24559 27031 24565
rect 30558 24556 30564 24608
rect 30616 24596 30622 24608
rect 30745 24599 30803 24605
rect 30745 24596 30757 24599
rect 30616 24568 30757 24596
rect 30616 24556 30622 24568
rect 30745 24565 30757 24568
rect 30791 24596 30803 24599
rect 30834 24596 30840 24608
rect 30791 24568 30840 24596
rect 30791 24565 30803 24568
rect 30745 24559 30803 24565
rect 30834 24556 30840 24568
rect 30892 24556 30898 24608
rect 31110 24556 31116 24608
rect 31168 24596 31174 24608
rect 31297 24599 31355 24605
rect 31297 24596 31309 24599
rect 31168 24568 31309 24596
rect 31168 24556 31174 24568
rect 31297 24565 31309 24568
rect 31343 24565 31355 24599
rect 31297 24559 31355 24565
rect 31846 24556 31852 24608
rect 31904 24596 31910 24608
rect 32493 24599 32551 24605
rect 32493 24596 32505 24599
rect 31904 24568 32505 24596
rect 31904 24556 31910 24568
rect 32493 24565 32505 24568
rect 32539 24565 32551 24599
rect 32493 24559 32551 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1581 24395 1639 24401
rect 1581 24361 1593 24395
rect 1627 24392 1639 24395
rect 2866 24392 2872 24404
rect 1627 24364 2872 24392
rect 1627 24361 1639 24364
rect 1581 24355 1639 24361
rect 2866 24352 2872 24364
rect 2924 24352 2930 24404
rect 3234 24352 3240 24404
rect 3292 24392 3298 24404
rect 3881 24395 3939 24401
rect 3881 24392 3893 24395
rect 3292 24364 3893 24392
rect 3292 24352 3298 24364
rect 3881 24361 3893 24364
rect 3927 24361 3939 24395
rect 3881 24355 3939 24361
rect 4341 24395 4399 24401
rect 4341 24361 4353 24395
rect 4387 24392 4399 24395
rect 5074 24392 5080 24404
rect 4387 24364 5080 24392
rect 4387 24361 4399 24364
rect 4341 24355 4399 24361
rect 5074 24352 5080 24364
rect 5132 24352 5138 24404
rect 14277 24395 14335 24401
rect 14277 24361 14289 24395
rect 14323 24392 14335 24395
rect 15838 24392 15844 24404
rect 14323 24364 15844 24392
rect 14323 24361 14335 24364
rect 14277 24355 14335 24361
rect 15838 24352 15844 24364
rect 15896 24352 15902 24404
rect 17126 24392 17132 24404
rect 16132 24364 16804 24392
rect 17087 24364 17132 24392
rect 3050 24284 3056 24336
rect 3108 24324 3114 24336
rect 9766 24324 9772 24336
rect 3108 24296 9772 24324
rect 3108 24284 3114 24296
rect 9766 24284 9772 24296
rect 9824 24284 9830 24336
rect 16132 24324 16160 24364
rect 16669 24327 16727 24333
rect 16669 24324 16681 24327
rect 10980 24296 16160 24324
rect 16224 24296 16681 24324
rect 4249 24259 4307 24265
rect 4249 24225 4261 24259
rect 4295 24256 4307 24259
rect 4614 24256 4620 24268
rect 4295 24228 4620 24256
rect 4295 24225 4307 24228
rect 4249 24219 4307 24225
rect 4614 24216 4620 24228
rect 4672 24216 4678 24268
rect 4890 24216 4896 24268
rect 4948 24256 4954 24268
rect 10980 24256 11008 24296
rect 4948 24228 11008 24256
rect 4948 24216 4954 24228
rect 15654 24216 15660 24268
rect 15712 24256 15718 24268
rect 16224 24265 16252 24296
rect 16669 24293 16681 24296
rect 16715 24293 16727 24327
rect 16776 24324 16804 24364
rect 17126 24352 17132 24364
rect 17184 24352 17190 24404
rect 18138 24392 18144 24404
rect 18099 24364 18144 24392
rect 18138 24352 18144 24364
rect 18196 24352 18202 24404
rect 18325 24395 18383 24401
rect 18325 24361 18337 24395
rect 18371 24392 18383 24395
rect 19242 24392 19248 24404
rect 18371 24364 19248 24392
rect 18371 24361 18383 24364
rect 18325 24355 18383 24361
rect 19242 24352 19248 24364
rect 19300 24352 19306 24404
rect 22922 24392 22928 24404
rect 22066 24364 22784 24392
rect 22883 24364 22928 24392
rect 22066 24324 22094 24364
rect 16776 24296 22094 24324
rect 22756 24324 22784 24364
rect 22922 24352 22928 24364
rect 22980 24352 22986 24404
rect 23845 24395 23903 24401
rect 23845 24361 23857 24395
rect 23891 24392 23903 24395
rect 25406 24392 25412 24404
rect 23891 24364 25412 24392
rect 23891 24361 23903 24364
rect 23845 24355 23903 24361
rect 25406 24352 25412 24364
rect 25464 24392 25470 24404
rect 25593 24395 25651 24401
rect 25593 24392 25605 24395
rect 25464 24364 25605 24392
rect 25464 24352 25470 24364
rect 25593 24361 25605 24364
rect 25639 24361 25651 24395
rect 25593 24355 25651 24361
rect 26053 24395 26111 24401
rect 26053 24361 26065 24395
rect 26099 24392 26111 24395
rect 26970 24392 26976 24404
rect 26099 24364 26976 24392
rect 26099 24361 26111 24364
rect 26053 24355 26111 24361
rect 26970 24352 26976 24364
rect 27028 24352 27034 24404
rect 30650 24352 30656 24404
rect 30708 24392 30714 24404
rect 36630 24392 36636 24404
rect 30708 24364 36636 24392
rect 30708 24352 30714 24364
rect 36630 24352 36636 24364
rect 36688 24352 36694 24404
rect 23474 24324 23480 24336
rect 22756 24296 23480 24324
rect 16669 24287 16727 24293
rect 23474 24284 23480 24296
rect 23532 24284 23538 24336
rect 24581 24327 24639 24333
rect 24581 24293 24593 24327
rect 24627 24293 24639 24327
rect 24581 24287 24639 24293
rect 15933 24259 15991 24265
rect 15933 24256 15945 24259
rect 15712 24228 15945 24256
rect 15712 24216 15718 24228
rect 15933 24225 15945 24228
rect 15979 24225 15991 24259
rect 15933 24219 15991 24225
rect 16209 24259 16267 24265
rect 16209 24225 16221 24259
rect 16255 24225 16267 24259
rect 16209 24219 16267 24225
rect 16390 24216 16396 24268
rect 16448 24256 16454 24268
rect 16942 24256 16948 24268
rect 16448 24228 16948 24256
rect 16448 24216 16454 24228
rect 16942 24216 16948 24228
rect 17000 24256 17006 24268
rect 17957 24259 18015 24265
rect 17957 24256 17969 24259
rect 17000 24228 17969 24256
rect 17000 24216 17006 24228
rect 17957 24225 17969 24228
rect 18003 24256 18015 24259
rect 21634 24256 21640 24268
rect 18003 24228 19334 24256
rect 18003 24225 18015 24228
rect 17957 24219 18015 24225
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24188 1458 24200
rect 2041 24191 2099 24197
rect 2041 24188 2053 24191
rect 1452 24160 2053 24188
rect 1452 24148 1458 24160
rect 2041 24157 2053 24160
rect 2087 24157 2099 24191
rect 2041 24151 2099 24157
rect 4065 24191 4123 24197
rect 4065 24157 4077 24191
rect 4111 24188 4123 24191
rect 4798 24188 4804 24200
rect 4111 24160 4804 24188
rect 4111 24157 4123 24160
rect 4065 24151 4123 24157
rect 4798 24148 4804 24160
rect 4856 24148 4862 24200
rect 4985 24191 5043 24197
rect 4985 24157 4997 24191
rect 5031 24188 5043 24191
rect 5442 24188 5448 24200
rect 5031 24160 5448 24188
rect 5031 24157 5043 24160
rect 4985 24151 5043 24157
rect 5442 24148 5448 24160
rect 5500 24148 5506 24200
rect 5629 24191 5687 24197
rect 5629 24157 5641 24191
rect 5675 24188 5687 24191
rect 6089 24191 6147 24197
rect 6089 24188 6101 24191
rect 5675 24160 6101 24188
rect 5675 24157 5687 24160
rect 5629 24151 5687 24157
rect 6089 24157 6101 24160
rect 6135 24188 6147 24191
rect 6638 24188 6644 24200
rect 6135 24160 6644 24188
rect 6135 24157 6147 24160
rect 6089 24151 6147 24157
rect 6638 24148 6644 24160
rect 6696 24148 6702 24200
rect 16850 24188 16856 24200
rect 16811 24160 16856 24188
rect 16850 24148 16856 24160
rect 16908 24148 16914 24200
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24188 18199 24191
rect 18506 24188 18512 24200
rect 18187 24160 18512 24188
rect 18187 24157 18199 24160
rect 18141 24151 18199 24157
rect 18506 24148 18512 24160
rect 18564 24148 18570 24200
rect 4341 24123 4399 24129
rect 4341 24089 4353 24123
rect 4387 24120 4399 24123
rect 4706 24120 4712 24132
rect 4387 24092 4712 24120
rect 4387 24089 4399 24092
rect 4341 24083 4399 24089
rect 4706 24080 4712 24092
rect 4764 24080 4770 24132
rect 4816 24120 4844 24148
rect 4816 24092 5488 24120
rect 4614 24012 4620 24064
rect 4672 24052 4678 24064
rect 5460 24061 5488 24092
rect 16666 24080 16672 24132
rect 16724 24120 16730 24132
rect 17129 24123 17187 24129
rect 17129 24120 17141 24123
rect 16724 24092 17141 24120
rect 16724 24080 16730 24092
rect 17129 24089 17141 24092
rect 17175 24120 17187 24123
rect 17310 24120 17316 24132
rect 17175 24092 17316 24120
rect 17175 24089 17187 24092
rect 17129 24083 17187 24089
rect 17310 24080 17316 24092
rect 17368 24120 17374 24132
rect 17865 24123 17923 24129
rect 17865 24120 17877 24123
rect 17368 24092 17877 24120
rect 17368 24080 17374 24092
rect 17865 24089 17877 24092
rect 17911 24089 17923 24123
rect 19306 24120 19334 24228
rect 19444 24228 21640 24256
rect 19444 24197 19472 24228
rect 21634 24216 21640 24228
rect 21692 24216 21698 24268
rect 21729 24259 21787 24265
rect 21729 24225 21741 24259
rect 21775 24256 21787 24259
rect 23106 24256 23112 24268
rect 21775 24228 23112 24256
rect 21775 24225 21787 24228
rect 21729 24219 21787 24225
rect 23106 24216 23112 24228
rect 23164 24216 23170 24268
rect 24596 24256 24624 24287
rect 25682 24256 25688 24268
rect 24596 24228 25688 24256
rect 25682 24216 25688 24228
rect 25740 24256 25746 24268
rect 27525 24259 27583 24265
rect 25740 24228 25912 24256
rect 25740 24216 25746 24228
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 19978 24148 19984 24200
rect 20036 24188 20042 24200
rect 20165 24191 20223 24197
rect 20165 24188 20177 24191
rect 20036 24160 20177 24188
rect 20036 24148 20042 24160
rect 20165 24157 20177 24160
rect 20211 24157 20223 24191
rect 20165 24151 20223 24157
rect 20346 24148 20352 24200
rect 20404 24188 20410 24200
rect 20441 24191 20499 24197
rect 20441 24188 20453 24191
rect 20404 24160 20453 24188
rect 20404 24148 20410 24160
rect 20441 24157 20453 24160
rect 20487 24188 20499 24191
rect 21453 24191 21511 24197
rect 21453 24188 21465 24191
rect 20487 24160 21465 24188
rect 20487 24157 20499 24160
rect 20441 24151 20499 24157
rect 21453 24157 21465 24160
rect 21499 24188 21511 24191
rect 21818 24188 21824 24200
rect 21499 24160 21824 24188
rect 21499 24157 21511 24160
rect 21453 24151 21511 24157
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 22002 24148 22008 24200
rect 22060 24188 22066 24200
rect 22741 24191 22799 24197
rect 22741 24188 22753 24191
rect 22060 24160 22753 24188
rect 22060 24148 22066 24160
rect 22741 24157 22753 24160
rect 22787 24157 22799 24191
rect 23658 24188 23664 24200
rect 23619 24160 23664 24188
rect 22741 24151 22799 24157
rect 23658 24148 23664 24160
rect 23716 24148 23722 24200
rect 24302 24148 24308 24200
rect 24360 24188 24366 24200
rect 25884 24197 25912 24228
rect 27525 24225 27537 24259
rect 27571 24256 27583 24259
rect 29914 24256 29920 24268
rect 27571 24228 29920 24256
rect 27571 24225 27583 24228
rect 27525 24219 27583 24225
rect 29914 24216 29920 24228
rect 29972 24216 29978 24268
rect 32306 24256 32312 24268
rect 32267 24228 32312 24256
rect 32306 24216 32312 24228
rect 32364 24216 32370 24268
rect 33321 24259 33379 24265
rect 33321 24225 33333 24259
rect 33367 24256 33379 24259
rect 33594 24256 33600 24268
rect 33367 24228 33600 24256
rect 33367 24225 33379 24228
rect 33321 24219 33379 24225
rect 33594 24216 33600 24228
rect 33652 24216 33658 24268
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 24360 24160 24409 24188
rect 24360 24148 24366 24160
rect 24397 24157 24409 24160
rect 24443 24188 24455 24191
rect 25041 24191 25099 24197
rect 25041 24188 25053 24191
rect 24443 24160 25053 24188
rect 24443 24157 24455 24160
rect 24397 24151 24455 24157
rect 25041 24157 25053 24160
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 25777 24191 25835 24197
rect 25777 24157 25789 24191
rect 25823 24157 25835 24191
rect 25777 24151 25835 24157
rect 25869 24191 25927 24197
rect 25869 24157 25881 24191
rect 25915 24157 25927 24191
rect 26602 24188 26608 24200
rect 26563 24160 26608 24188
rect 25869 24151 25927 24157
rect 22462 24120 22468 24132
rect 19306 24092 22468 24120
rect 17865 24083 17923 24089
rect 22462 24080 22468 24092
rect 22520 24080 22526 24132
rect 25222 24080 25228 24132
rect 25280 24120 25286 24132
rect 25593 24123 25651 24129
rect 25593 24120 25605 24123
rect 25280 24092 25605 24120
rect 25280 24080 25286 24092
rect 25593 24089 25605 24092
rect 25639 24089 25651 24123
rect 25792 24120 25820 24151
rect 26602 24148 26608 24160
rect 26660 24148 26666 24200
rect 27062 24148 27068 24200
rect 27120 24188 27126 24200
rect 27249 24191 27307 24197
rect 27249 24188 27261 24191
rect 27120 24160 27261 24188
rect 27120 24148 27126 24160
rect 27249 24157 27261 24160
rect 27295 24157 27307 24191
rect 27249 24151 27307 24157
rect 32585 24191 32643 24197
rect 32585 24157 32597 24191
rect 32631 24188 32643 24191
rect 32674 24188 32680 24200
rect 32631 24160 32680 24188
rect 32631 24157 32643 24160
rect 32585 24151 32643 24157
rect 32674 24148 32680 24160
rect 32732 24148 32738 24200
rect 33502 24188 33508 24200
rect 33463 24160 33508 24188
rect 33502 24148 33508 24160
rect 33560 24148 33566 24200
rect 26234 24120 26240 24132
rect 25792 24092 26240 24120
rect 25593 24083 25651 24089
rect 26234 24080 26240 24092
rect 26292 24120 26298 24132
rect 26970 24120 26976 24132
rect 26292 24092 26976 24120
rect 26292 24080 26298 24092
rect 26970 24080 26976 24092
rect 27028 24080 27034 24132
rect 4801 24055 4859 24061
rect 4801 24052 4813 24055
rect 4672 24024 4813 24052
rect 4672 24012 4678 24024
rect 4801 24021 4813 24024
rect 4847 24021 4859 24055
rect 4801 24015 4859 24021
rect 5445 24055 5503 24061
rect 5445 24021 5457 24055
rect 5491 24021 5503 24055
rect 19242 24052 19248 24064
rect 19203 24024 19248 24052
rect 5445 24015 5503 24021
rect 19242 24012 19248 24024
rect 19300 24012 19306 24064
rect 26789 24055 26847 24061
rect 26789 24021 26801 24055
rect 26835 24052 26847 24055
rect 29822 24052 29828 24064
rect 26835 24024 29828 24052
rect 26835 24021 26847 24024
rect 26789 24015 26847 24021
rect 29822 24012 29828 24024
rect 29880 24012 29886 24064
rect 33689 24055 33747 24061
rect 33689 24021 33701 24055
rect 33735 24052 33747 24055
rect 34330 24052 34336 24064
rect 33735 24024 34336 24052
rect 33735 24021 33747 24024
rect 33689 24015 33747 24021
rect 34330 24012 34336 24024
rect 34388 24012 34394 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 16850 23808 16856 23860
rect 16908 23848 16914 23860
rect 16908 23820 16988 23848
rect 16908 23808 16914 23820
rect 16960 23780 16988 23820
rect 17218 23808 17224 23860
rect 17276 23848 17282 23860
rect 17589 23851 17647 23857
rect 17589 23848 17601 23851
rect 17276 23820 17601 23848
rect 17276 23808 17282 23820
rect 17589 23817 17601 23820
rect 17635 23817 17647 23851
rect 17589 23811 17647 23817
rect 17788 23820 22140 23848
rect 17788 23780 17816 23820
rect 16960 23752 17816 23780
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 4982 23712 4988 23724
rect 4847 23684 4988 23712
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 4982 23672 4988 23684
rect 5040 23712 5046 23724
rect 5258 23712 5264 23724
rect 5040 23684 5264 23712
rect 5040 23672 5046 23684
rect 5258 23672 5264 23684
rect 5316 23672 5322 23724
rect 5442 23672 5448 23724
rect 5500 23712 5506 23724
rect 6730 23712 6736 23724
rect 5500 23684 6736 23712
rect 5500 23672 5506 23684
rect 6730 23672 6736 23684
rect 6788 23712 6794 23724
rect 7193 23715 7251 23721
rect 7193 23712 7205 23715
rect 6788 23684 7205 23712
rect 6788 23672 6794 23684
rect 7193 23681 7205 23684
rect 7239 23681 7251 23715
rect 7193 23675 7251 23681
rect 16850 23672 16856 23724
rect 16908 23721 16914 23724
rect 16908 23712 16918 23721
rect 17129 23715 17187 23721
rect 16908 23684 16953 23712
rect 16908 23675 16918 23684
rect 17129 23681 17141 23715
rect 17175 23712 17187 23715
rect 17310 23712 17316 23724
rect 17175 23684 17316 23712
rect 17175 23681 17187 23684
rect 17129 23675 17187 23681
rect 16908 23672 16914 23675
rect 16942 23644 16948 23656
rect 16903 23616 16948 23644
rect 16942 23604 16948 23616
rect 17000 23604 17006 23656
rect 17034 23604 17040 23656
rect 17092 23644 17098 23656
rect 17144 23644 17172 23675
rect 17310 23672 17316 23684
rect 17368 23672 17374 23724
rect 17788 23721 17816 23752
rect 18049 23783 18107 23789
rect 18049 23749 18061 23783
rect 18095 23780 18107 23783
rect 18230 23780 18236 23792
rect 18095 23752 18236 23780
rect 18095 23749 18107 23752
rect 18049 23743 18107 23749
rect 18230 23740 18236 23752
rect 18288 23780 18294 23792
rect 19242 23780 19248 23792
rect 18288 23752 19248 23780
rect 18288 23740 18294 23752
rect 19242 23740 19248 23752
rect 19300 23740 19306 23792
rect 22112 23780 22140 23820
rect 23658 23808 23664 23860
rect 23716 23848 23722 23860
rect 24029 23851 24087 23857
rect 24029 23848 24041 23851
rect 23716 23820 24041 23848
rect 23716 23808 23722 23820
rect 24029 23817 24041 23820
rect 24075 23817 24087 23851
rect 24029 23811 24087 23817
rect 25222 23808 25228 23860
rect 25280 23848 25286 23860
rect 26050 23848 26056 23860
rect 25280 23820 26056 23848
rect 25280 23808 25286 23820
rect 26050 23808 26056 23820
rect 26108 23848 26114 23860
rect 27617 23851 27675 23857
rect 27617 23848 27629 23851
rect 26108 23820 27629 23848
rect 26108 23808 26114 23820
rect 27617 23817 27629 23820
rect 27663 23817 27675 23851
rect 27617 23811 27675 23817
rect 29822 23780 29828 23792
rect 22112 23752 23428 23780
rect 29783 23752 29828 23780
rect 17773 23715 17831 23721
rect 17773 23681 17785 23715
rect 17819 23681 17831 23715
rect 18966 23712 18972 23724
rect 17773 23675 17831 23681
rect 18156 23684 18972 23712
rect 17092 23616 17172 23644
rect 17865 23647 17923 23653
rect 17092 23604 17098 23616
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 18046 23644 18052 23656
rect 17911 23616 18052 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18046 23604 18052 23616
rect 18104 23604 18110 23656
rect 7377 23579 7435 23585
rect 7377 23545 7389 23579
rect 7423 23576 7435 23579
rect 7742 23576 7748 23588
rect 7423 23548 7748 23576
rect 7423 23545 7435 23548
rect 7377 23539 7435 23545
rect 7742 23536 7748 23548
rect 7800 23576 7806 23588
rect 18156 23576 18184 23684
rect 18966 23672 18972 23684
rect 19024 23672 19030 23724
rect 19069 23715 19127 23721
rect 19069 23681 19081 23715
rect 19115 23712 19127 23715
rect 20162 23712 20168 23724
rect 19115 23684 20168 23712
rect 19115 23681 19127 23684
rect 19069 23675 19127 23681
rect 20162 23672 20168 23684
rect 20220 23672 20226 23724
rect 20346 23712 20352 23724
rect 20307 23684 20352 23712
rect 20346 23672 20352 23684
rect 20404 23672 20410 23724
rect 22112 23721 22140 23752
rect 23400 23724 23428 23752
rect 29822 23740 29828 23752
rect 29880 23740 29886 23792
rect 22097 23715 22155 23721
rect 22097 23681 22109 23715
rect 22143 23681 22155 23715
rect 22097 23675 22155 23681
rect 22922 23672 22928 23724
rect 22980 23712 22986 23724
rect 23109 23715 23167 23721
rect 23109 23712 23121 23715
rect 22980 23684 23121 23712
rect 22980 23672 22986 23684
rect 23109 23681 23121 23684
rect 23155 23681 23167 23715
rect 23382 23712 23388 23724
rect 23343 23684 23388 23712
rect 23109 23675 23167 23681
rect 23382 23672 23388 23684
rect 23440 23672 23446 23724
rect 25869 23715 25927 23721
rect 25869 23712 25881 23715
rect 23492 23684 25881 23712
rect 19150 23644 19156 23656
rect 7800 23548 18184 23576
rect 18248 23616 19156 23644
rect 7800 23536 7806 23548
rect 4617 23511 4675 23517
rect 4617 23477 4629 23511
rect 4663 23508 4675 23511
rect 4706 23508 4712 23520
rect 4663 23480 4712 23508
rect 4663 23477 4675 23480
rect 4617 23471 4675 23477
rect 4706 23468 4712 23480
rect 4764 23468 4770 23520
rect 12345 23511 12403 23517
rect 12345 23477 12357 23511
rect 12391 23508 12403 23511
rect 12894 23508 12900 23520
rect 12391 23480 12900 23508
rect 12391 23477 12403 23480
rect 12345 23471 12403 23477
rect 12894 23468 12900 23480
rect 12952 23468 12958 23520
rect 15286 23508 15292 23520
rect 15247 23480 15292 23508
rect 15286 23468 15292 23480
rect 15344 23468 15350 23520
rect 16022 23468 16028 23520
rect 16080 23508 16086 23520
rect 16669 23511 16727 23517
rect 16669 23508 16681 23511
rect 16080 23480 16681 23508
rect 16080 23468 16086 23480
rect 16669 23477 16681 23480
rect 16715 23477 16727 23511
rect 17126 23508 17132 23520
rect 17039 23480 17132 23508
rect 16669 23471 16727 23477
rect 17126 23468 17132 23480
rect 17184 23508 17190 23520
rect 18049 23511 18107 23517
rect 18049 23508 18061 23511
rect 17184 23480 18061 23508
rect 17184 23468 17190 23480
rect 18049 23477 18061 23480
rect 18095 23508 18107 23511
rect 18248 23508 18276 23616
rect 19150 23604 19156 23616
rect 19208 23604 19214 23656
rect 19242 23604 19248 23656
rect 19300 23644 19306 23656
rect 20073 23647 20131 23653
rect 20073 23644 20085 23647
rect 19300 23616 20085 23644
rect 19300 23604 19306 23616
rect 20073 23613 20085 23616
rect 20119 23613 20131 23647
rect 20180 23644 20208 23672
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 20180 23616 21833 23644
rect 20073 23607 20131 23613
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 21821 23607 21879 23613
rect 22462 23604 22468 23656
rect 22520 23644 22526 23656
rect 23201 23647 23259 23653
rect 23201 23644 23213 23647
rect 22520 23616 23213 23644
rect 22520 23604 22526 23616
rect 23201 23613 23213 23616
rect 23247 23613 23259 23647
rect 23492 23644 23520 23684
rect 25869 23681 25881 23684
rect 25915 23712 25927 23715
rect 26234 23712 26240 23724
rect 25915 23684 26240 23712
rect 25915 23681 25927 23684
rect 25869 23675 25927 23681
rect 26234 23672 26240 23684
rect 26292 23672 26298 23724
rect 30009 23715 30067 23721
rect 30009 23681 30021 23715
rect 30055 23712 30067 23715
rect 30650 23712 30656 23724
rect 30055 23684 30656 23712
rect 30055 23681 30067 23684
rect 30009 23675 30067 23681
rect 30650 23672 30656 23684
rect 30708 23672 30714 23724
rect 34330 23712 34336 23724
rect 34291 23684 34336 23712
rect 34330 23672 34336 23684
rect 34388 23672 34394 23724
rect 23201 23607 23259 23613
rect 23308 23616 23520 23644
rect 24581 23647 24639 23653
rect 18506 23536 18512 23588
rect 18564 23576 18570 23588
rect 18877 23579 18935 23585
rect 18877 23576 18889 23579
rect 18564 23548 18889 23576
rect 18564 23536 18570 23548
rect 18877 23545 18889 23548
rect 18923 23545 18935 23579
rect 18877 23539 18935 23545
rect 18966 23536 18972 23588
rect 19024 23576 19030 23588
rect 23308 23576 23336 23616
rect 24581 23613 24593 23647
rect 24627 23613 24639 23647
rect 24854 23644 24860 23656
rect 24815 23616 24860 23644
rect 24581 23607 24639 23613
rect 19024 23548 23336 23576
rect 23569 23579 23627 23585
rect 19024 23536 19030 23548
rect 23569 23545 23581 23579
rect 23615 23576 23627 23579
rect 24596 23576 24624 23607
rect 24854 23604 24860 23616
rect 24912 23604 24918 23656
rect 28166 23644 28172 23656
rect 28127 23616 28172 23644
rect 28166 23604 28172 23616
rect 28224 23604 28230 23656
rect 23615 23548 24624 23576
rect 23615 23545 23627 23548
rect 23569 23539 23627 23545
rect 18095 23480 18276 23508
rect 18095 23477 18107 23480
rect 18049 23471 18107 23477
rect 19150 23468 19156 23520
rect 19208 23508 19214 23520
rect 23106 23508 23112 23520
rect 19208 23480 23112 23508
rect 19208 23468 19214 23480
rect 23106 23468 23112 23480
rect 23164 23468 23170 23520
rect 27062 23508 27068 23520
rect 27023 23480 27068 23508
rect 27062 23468 27068 23480
rect 27120 23468 27126 23520
rect 30466 23508 30472 23520
rect 30427 23480 30472 23508
rect 30466 23468 30472 23480
rect 30524 23468 30530 23520
rect 32674 23508 32680 23520
rect 32635 23480 32680 23508
rect 32674 23468 32680 23480
rect 32732 23468 32738 23520
rect 34514 23508 34520 23520
rect 34475 23480 34520 23508
rect 34514 23468 34520 23480
rect 34572 23468 34578 23520
rect 34790 23468 34796 23520
rect 34848 23508 34854 23520
rect 34977 23511 35035 23517
rect 34977 23508 34989 23511
rect 34848 23480 34989 23508
rect 34848 23468 34854 23480
rect 34977 23477 34989 23480
rect 35023 23477 35035 23511
rect 34977 23471 35035 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 4433 23307 4491 23313
rect 4433 23273 4445 23307
rect 4479 23304 4491 23307
rect 4798 23304 4804 23316
rect 4479 23276 4804 23304
rect 4479 23273 4491 23276
rect 4433 23267 4491 23273
rect 4798 23264 4804 23276
rect 4856 23264 4862 23316
rect 6638 23304 6644 23316
rect 6599 23276 6644 23304
rect 6638 23264 6644 23276
rect 6696 23264 6702 23316
rect 12526 23304 12532 23316
rect 12487 23276 12532 23304
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 13262 23304 13268 23316
rect 13223 23276 13268 23304
rect 13262 23264 13268 23276
rect 13320 23264 13326 23316
rect 17773 23307 17831 23313
rect 17773 23273 17785 23307
rect 17819 23304 17831 23307
rect 18138 23304 18144 23316
rect 17819 23276 18144 23304
rect 17819 23273 17831 23276
rect 17773 23267 17831 23273
rect 18138 23264 18144 23276
rect 18196 23304 18202 23316
rect 18509 23307 18567 23313
rect 18509 23304 18521 23307
rect 18196 23276 18521 23304
rect 18196 23264 18202 23276
rect 18509 23273 18521 23276
rect 18555 23304 18567 23307
rect 19242 23304 19248 23316
rect 18555 23276 19248 23304
rect 18555 23273 18567 23276
rect 18509 23267 18567 23273
rect 19242 23264 19248 23276
rect 19300 23264 19306 23316
rect 20346 23304 20352 23316
rect 20307 23276 20352 23304
rect 20346 23264 20352 23276
rect 20404 23264 20410 23316
rect 36078 23264 36084 23316
rect 36136 23304 36142 23316
rect 36173 23307 36231 23313
rect 36173 23304 36185 23307
rect 36136 23276 36185 23304
rect 36136 23264 36142 23276
rect 36173 23273 36185 23276
rect 36219 23273 36231 23307
rect 36173 23267 36231 23273
rect 3973 23239 4031 23245
rect 3973 23205 3985 23239
rect 4019 23205 4031 23239
rect 13280 23236 13308 23264
rect 19978 23236 19984 23248
rect 13280 23208 19984 23236
rect 3973 23199 4031 23205
rect 1394 23100 1400 23112
rect 1355 23072 1400 23100
rect 1394 23060 1400 23072
rect 1452 23060 1458 23112
rect 2593 23103 2651 23109
rect 2593 23069 2605 23103
rect 2639 23100 2651 23103
rect 2774 23100 2780 23112
rect 2639 23072 2780 23100
rect 2639 23069 2651 23072
rect 2593 23063 2651 23069
rect 2774 23060 2780 23072
rect 2832 23060 2838 23112
rect 3237 23103 3295 23109
rect 3237 23069 3249 23103
rect 3283 23100 3295 23103
rect 3988 23100 4016 23199
rect 19978 23196 19984 23208
rect 20036 23196 20042 23248
rect 4341 23171 4399 23177
rect 4341 23137 4353 23171
rect 4387 23168 4399 23171
rect 4614 23168 4620 23180
rect 4387 23140 4620 23168
rect 4387 23137 4399 23140
rect 4341 23131 4399 23137
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 10597 23171 10655 23177
rect 10597 23168 10609 23171
rect 9272 23140 10609 23168
rect 9272 23128 9278 23140
rect 10597 23137 10609 23140
rect 10643 23137 10655 23171
rect 10597 23131 10655 23137
rect 15286 23128 15292 23180
rect 15344 23168 15350 23180
rect 16853 23171 16911 23177
rect 16853 23168 16865 23171
rect 15344 23140 16865 23168
rect 15344 23128 15350 23140
rect 16853 23137 16865 23140
rect 16899 23137 16911 23171
rect 17678 23168 17684 23180
rect 17591 23140 17684 23168
rect 16853 23131 16911 23137
rect 17678 23128 17684 23140
rect 17736 23168 17742 23180
rect 18325 23171 18383 23177
rect 18325 23168 18337 23171
rect 17736 23140 18337 23168
rect 17736 23128 17742 23140
rect 18325 23137 18337 23140
rect 18371 23137 18383 23171
rect 18325 23131 18383 23137
rect 20257 23171 20315 23177
rect 20257 23137 20269 23171
rect 20303 23168 20315 23171
rect 24486 23168 24492 23180
rect 20303 23140 24492 23168
rect 20303 23137 20315 23140
rect 20257 23131 20315 23137
rect 24486 23128 24492 23140
rect 24544 23128 24550 23180
rect 24854 23128 24860 23180
rect 24912 23168 24918 23180
rect 27433 23171 27491 23177
rect 27433 23168 27445 23171
rect 24912 23140 27445 23168
rect 24912 23128 24918 23140
rect 27433 23137 27445 23140
rect 27479 23137 27491 23171
rect 27433 23131 27491 23137
rect 27617 23171 27675 23177
rect 27617 23137 27629 23171
rect 27663 23168 27675 23171
rect 29730 23168 29736 23180
rect 27663 23140 29736 23168
rect 27663 23137 27675 23140
rect 27617 23131 27675 23137
rect 29730 23128 29736 23140
rect 29788 23128 29794 23180
rect 30653 23171 30711 23177
rect 30653 23137 30665 23171
rect 30699 23168 30711 23171
rect 30926 23168 30932 23180
rect 30699 23140 30932 23168
rect 30699 23137 30711 23140
rect 30653 23131 30711 23137
rect 30926 23128 30932 23140
rect 30984 23128 30990 23180
rect 4154 23100 4160 23112
rect 3283 23072 4016 23100
rect 4115 23072 4160 23100
rect 3283 23069 3295 23072
rect 3237 23063 3295 23069
rect 4154 23060 4160 23072
rect 4212 23060 4218 23112
rect 4982 23060 4988 23112
rect 5040 23100 5046 23112
rect 7653 23103 7711 23109
rect 7653 23100 7665 23103
rect 5040 23072 7665 23100
rect 5040 23060 5046 23072
rect 7653 23069 7665 23072
rect 7699 23069 7711 23103
rect 10870 23100 10876 23112
rect 10831 23072 10876 23100
rect 7653 23063 7711 23069
rect 10870 23060 10876 23072
rect 10928 23060 10934 23112
rect 11330 23100 11336 23112
rect 11291 23072 11336 23100
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 12713 23103 12771 23109
rect 12713 23069 12725 23103
rect 12759 23100 12771 23103
rect 12894 23100 12900 23112
rect 12759 23072 12900 23100
rect 12759 23069 12771 23072
rect 12713 23063 12771 23069
rect 12894 23060 12900 23072
rect 12952 23060 12958 23112
rect 13449 23103 13507 23109
rect 13449 23069 13461 23103
rect 13495 23100 13507 23103
rect 13998 23100 14004 23112
rect 13495 23072 14004 23100
rect 13495 23069 13507 23072
rect 13449 23063 13507 23069
rect 13998 23060 14004 23072
rect 14056 23060 14062 23112
rect 17497 23103 17555 23109
rect 17497 23069 17509 23103
rect 17543 23069 17555 23103
rect 17497 23063 17555 23069
rect 17773 23103 17831 23109
rect 17773 23069 17785 23103
rect 17819 23100 17831 23103
rect 18230 23100 18236 23112
rect 17819 23072 18236 23100
rect 17819 23069 17831 23072
rect 17773 23063 17831 23069
rect 4433 23035 4491 23041
rect 4433 23001 4445 23035
rect 4479 23032 4491 23035
rect 4706 23032 4712 23044
rect 4479 23004 4712 23032
rect 4479 23001 4491 23004
rect 4433 22995 4491 23001
rect 4706 22992 4712 23004
rect 4764 22992 4770 23044
rect 7834 23032 7840 23044
rect 7795 23004 7840 23032
rect 7834 22992 7840 23004
rect 7892 22992 7898 23044
rect 15013 23035 15071 23041
rect 15013 23001 15025 23035
rect 15059 23032 15071 23035
rect 15286 23032 15292 23044
rect 15059 23004 15292 23032
rect 15059 23001 15071 23004
rect 15013 22995 15071 23001
rect 15286 22992 15292 23004
rect 15344 22992 15350 23044
rect 16666 23032 16672 23044
rect 16627 23004 16672 23032
rect 16666 22992 16672 23004
rect 16724 22992 16730 23044
rect 17512 23032 17540 23063
rect 18230 23060 18236 23072
rect 18288 23060 18294 23112
rect 18506 23100 18512 23112
rect 18467 23072 18512 23100
rect 18506 23060 18512 23072
rect 18564 23060 18570 23112
rect 20162 23060 20168 23112
rect 20220 23100 20226 23112
rect 20349 23103 20407 23109
rect 20349 23100 20361 23103
rect 20220 23072 20361 23100
rect 20220 23060 20226 23072
rect 20349 23069 20361 23072
rect 20395 23069 20407 23103
rect 29914 23100 29920 23112
rect 29875 23072 29920 23100
rect 20349 23063 20407 23069
rect 29914 23060 29920 23072
rect 29972 23060 29978 23112
rect 30834 23100 30840 23112
rect 30795 23072 30840 23100
rect 30834 23060 30840 23072
rect 30892 23060 30898 23112
rect 31021 23103 31079 23109
rect 31021 23069 31033 23103
rect 31067 23100 31079 23103
rect 31665 23103 31723 23109
rect 31665 23100 31677 23103
rect 31067 23072 31677 23100
rect 31067 23069 31079 23072
rect 31021 23063 31079 23069
rect 31665 23069 31677 23072
rect 31711 23069 31723 23103
rect 31665 23063 31723 23069
rect 33870 23060 33876 23112
rect 33928 23100 33934 23112
rect 33965 23103 34023 23109
rect 33965 23100 33977 23103
rect 33928 23072 33977 23100
rect 33928 23060 33934 23072
rect 33965 23069 33977 23072
rect 34011 23069 34023 23103
rect 34790 23100 34796 23112
rect 34751 23072 34796 23100
rect 33965 23063 34023 23069
rect 34790 23060 34796 23072
rect 34848 23060 34854 23112
rect 18524 23032 18552 23060
rect 17512 23004 18552 23032
rect 18966 22992 18972 23044
rect 19024 23032 19030 23044
rect 20073 23035 20131 23041
rect 20073 23032 20085 23035
rect 19024 23004 20085 23032
rect 19024 22992 19030 23004
rect 20073 23001 20085 23004
rect 20119 23001 20131 23035
rect 20073 22995 20131 23001
rect 25777 23035 25835 23041
rect 25777 23001 25789 23035
rect 25823 23032 25835 23035
rect 25958 23032 25964 23044
rect 25823 23004 25964 23032
rect 25823 23001 25835 23004
rect 25777 22995 25835 23001
rect 25958 22992 25964 23004
rect 26016 22992 26022 23044
rect 35038 23035 35096 23041
rect 35038 23032 35050 23035
rect 34164 23004 35050 23032
rect 1578 22964 1584 22976
rect 1539 22936 1584 22964
rect 1578 22924 1584 22936
rect 1636 22924 1642 22976
rect 2958 22924 2964 22976
rect 3016 22964 3022 22976
rect 3053 22967 3111 22973
rect 3053 22964 3065 22967
rect 3016 22936 3065 22964
rect 3016 22924 3022 22936
rect 3053 22933 3065 22936
rect 3099 22933 3111 22967
rect 3053 22927 3111 22933
rect 16850 22924 16856 22976
rect 16908 22964 16914 22976
rect 17313 22967 17371 22973
rect 17313 22964 17325 22967
rect 16908 22936 17325 22964
rect 16908 22924 16914 22936
rect 17313 22933 17325 22936
rect 17359 22933 17371 22967
rect 17313 22927 17371 22933
rect 18693 22967 18751 22973
rect 18693 22933 18705 22967
rect 18739 22964 18751 22967
rect 19426 22964 19432 22976
rect 18739 22936 19432 22964
rect 18739 22933 18751 22936
rect 18693 22927 18751 22933
rect 19426 22924 19432 22936
rect 19484 22924 19490 22976
rect 20533 22967 20591 22973
rect 20533 22933 20545 22967
rect 20579 22964 20591 22967
rect 20806 22964 20812 22976
rect 20579 22936 20812 22964
rect 20579 22933 20591 22936
rect 20533 22927 20591 22933
rect 20806 22924 20812 22936
rect 20864 22924 20870 22976
rect 22922 22964 22928 22976
rect 22883 22936 22928 22964
rect 22922 22924 22928 22936
rect 22980 22924 22986 22976
rect 25222 22964 25228 22976
rect 25183 22936 25228 22964
rect 25222 22924 25228 22936
rect 25280 22924 25286 22976
rect 30098 22964 30104 22976
rect 30059 22936 30104 22964
rect 30098 22924 30104 22936
rect 30156 22924 30162 22976
rect 31478 22964 31484 22976
rect 31439 22936 31484 22964
rect 31478 22924 31484 22936
rect 31536 22924 31542 22976
rect 34164 22973 34192 23004
rect 35038 23001 35050 23004
rect 35084 23001 35096 23035
rect 35038 22995 35096 23001
rect 34149 22967 34207 22973
rect 34149 22933 34161 22967
rect 34195 22933 34207 22967
rect 34149 22927 34207 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 4154 22720 4160 22772
rect 4212 22760 4218 22772
rect 6365 22763 6423 22769
rect 6365 22760 6377 22763
rect 4212 22732 6377 22760
rect 4212 22720 4218 22732
rect 6365 22729 6377 22732
rect 6411 22729 6423 22763
rect 6365 22723 6423 22729
rect 7834 22720 7840 22772
rect 7892 22760 7898 22772
rect 8202 22760 8208 22772
rect 7892 22732 8208 22760
rect 7892 22720 7898 22732
rect 8202 22720 8208 22732
rect 8260 22760 8266 22772
rect 25222 22760 25228 22772
rect 8260 22732 25228 22760
rect 8260 22720 8266 22732
rect 25222 22720 25228 22732
rect 25280 22720 25286 22772
rect 29914 22760 29920 22772
rect 29875 22732 29920 22760
rect 29914 22720 29920 22732
rect 29972 22720 29978 22772
rect 30558 22720 30564 22772
rect 30616 22760 30622 22772
rect 30653 22763 30711 22769
rect 30653 22760 30665 22763
rect 30616 22732 30665 22760
rect 30616 22720 30622 22732
rect 30653 22729 30665 22732
rect 30699 22729 30711 22763
rect 30653 22723 30711 22729
rect 31113 22763 31171 22769
rect 31113 22729 31125 22763
rect 31159 22760 31171 22763
rect 33686 22760 33692 22772
rect 31159 22732 33692 22760
rect 31159 22729 31171 22732
rect 31113 22723 31171 22729
rect 33686 22720 33692 22732
rect 33744 22720 33750 22772
rect 33870 22760 33876 22772
rect 33831 22732 33876 22760
rect 33870 22720 33876 22732
rect 33928 22720 33934 22772
rect 1394 22692 1400 22704
rect 1355 22664 1400 22692
rect 1394 22652 1400 22664
rect 1452 22652 1458 22704
rect 2958 22692 2964 22704
rect 2919 22664 2964 22692
rect 2958 22652 2964 22664
rect 3016 22652 3022 22704
rect 7650 22692 7656 22704
rect 7563 22664 7656 22692
rect 7650 22652 7656 22664
rect 7708 22692 7714 22704
rect 18141 22695 18199 22701
rect 7708 22664 13124 22692
rect 7708 22652 7714 22664
rect 2774 22624 2780 22636
rect 2735 22596 2780 22624
rect 2774 22584 2780 22596
rect 2832 22584 2838 22636
rect 5258 22624 5264 22636
rect 5219 22596 5264 22624
rect 5258 22584 5264 22596
rect 5316 22584 5322 22636
rect 6549 22627 6607 22633
rect 6549 22593 6561 22627
rect 6595 22624 6607 22627
rect 6638 22624 6644 22636
rect 6595 22596 6644 22624
rect 6595 22593 6607 22596
rect 6549 22587 6607 22593
rect 6638 22584 6644 22596
rect 6696 22584 6702 22636
rect 9398 22584 9404 22636
rect 9456 22624 9462 22636
rect 10137 22627 10195 22633
rect 10137 22624 10149 22627
rect 9456 22596 10149 22624
rect 9456 22584 9462 22596
rect 10137 22593 10149 22596
rect 10183 22593 10195 22627
rect 10137 22587 10195 22593
rect 11517 22627 11575 22633
rect 11517 22593 11529 22627
rect 11563 22624 11575 22627
rect 12342 22624 12348 22636
rect 11563 22596 12348 22624
rect 11563 22593 11575 22596
rect 11517 22587 11575 22593
rect 12342 22584 12348 22596
rect 12400 22584 12406 22636
rect 3234 22556 3240 22568
rect 3195 22528 3240 22556
rect 3234 22516 3240 22528
rect 3292 22556 3298 22568
rect 9858 22556 9864 22568
rect 3292 22528 6914 22556
rect 9819 22528 9864 22556
rect 3292 22516 3298 22528
rect 6886 22488 6914 22528
rect 9858 22516 9864 22528
rect 9916 22516 9922 22568
rect 12526 22556 12532 22568
rect 11440 22528 12532 22556
rect 11440 22488 11468 22528
rect 12526 22516 12532 22528
rect 12584 22516 12590 22568
rect 6886 22460 11468 22488
rect 11514 22448 11520 22500
rect 11572 22488 11578 22500
rect 12161 22491 12219 22497
rect 12161 22488 12173 22491
rect 11572 22460 12173 22488
rect 11572 22448 11578 22460
rect 12161 22457 12173 22460
rect 12207 22457 12219 22491
rect 12161 22451 12219 22457
rect 5074 22420 5080 22432
rect 5035 22392 5080 22420
rect 5074 22380 5080 22392
rect 5132 22380 5138 22432
rect 5810 22420 5816 22432
rect 5771 22392 5816 22420
rect 5810 22380 5816 22392
rect 5868 22380 5874 22432
rect 7098 22420 7104 22432
rect 7059 22392 7104 22420
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 11698 22420 11704 22432
rect 11659 22392 11704 22420
rect 11698 22380 11704 22392
rect 11756 22380 11762 22432
rect 13096 22429 13124 22664
rect 18141 22661 18153 22695
rect 18187 22692 18199 22695
rect 18230 22692 18236 22704
rect 18187 22664 18236 22692
rect 18187 22661 18199 22664
rect 18141 22655 18199 22661
rect 18230 22652 18236 22664
rect 18288 22692 18294 22704
rect 19061 22695 19119 22701
rect 19061 22692 19073 22695
rect 18288 22664 19073 22692
rect 18288 22652 18294 22664
rect 19061 22661 19073 22664
rect 19107 22661 19119 22695
rect 23382 22692 23388 22704
rect 19061 22655 19119 22661
rect 23124 22664 23388 22692
rect 16022 22624 16028 22636
rect 15983 22596 16028 22624
rect 16022 22584 16028 22596
rect 16080 22584 16086 22636
rect 16850 22624 16856 22636
rect 16811 22596 16856 22624
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 17865 22627 17923 22633
rect 17865 22593 17877 22627
rect 17911 22624 17923 22627
rect 18506 22624 18512 22636
rect 17911 22596 18512 22624
rect 17911 22593 17923 22596
rect 17865 22587 17923 22593
rect 18506 22584 18512 22596
rect 18564 22624 18570 22636
rect 18785 22627 18843 22633
rect 18785 22624 18797 22627
rect 18564 22596 18797 22624
rect 18564 22584 18570 22596
rect 18785 22593 18797 22596
rect 18831 22593 18843 22627
rect 18785 22587 18843 22593
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 19521 22627 19579 22633
rect 19521 22624 19533 22627
rect 19484 22596 19533 22624
rect 19484 22584 19490 22596
rect 19521 22593 19533 22596
rect 19567 22593 19579 22627
rect 20806 22624 20812 22636
rect 20767 22596 20812 22624
rect 19521 22587 19579 22593
rect 20806 22584 20812 22596
rect 20864 22584 20870 22636
rect 22462 22584 22468 22636
rect 22520 22624 22526 22636
rect 22833 22627 22891 22633
rect 22833 22624 22845 22627
rect 22520 22596 22845 22624
rect 22520 22584 22526 22596
rect 22833 22593 22845 22596
rect 22879 22624 22891 22627
rect 22922 22624 22928 22636
rect 22879 22596 22928 22624
rect 22879 22593 22891 22596
rect 22833 22587 22891 22593
rect 22922 22584 22928 22596
rect 22980 22584 22986 22636
rect 23124 22633 23152 22664
rect 23382 22652 23388 22664
rect 23440 22652 23446 22704
rect 30926 22692 30932 22704
rect 29564 22664 30932 22692
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22593 23167 22627
rect 24765 22627 24823 22633
rect 24765 22624 24777 22627
rect 23109 22587 23167 22593
rect 23308 22596 24777 22624
rect 18046 22556 18052 22568
rect 17959 22528 18052 22556
rect 18046 22516 18052 22528
rect 18104 22556 18110 22568
rect 18230 22556 18236 22568
rect 18104 22528 18236 22556
rect 18104 22516 18110 22528
rect 18230 22516 18236 22528
rect 18288 22556 18294 22568
rect 18966 22556 18972 22568
rect 18288 22528 18972 22556
rect 18288 22516 18294 22528
rect 18966 22516 18972 22528
rect 19024 22516 19030 22568
rect 23017 22559 23075 22565
rect 23017 22525 23029 22559
rect 23063 22556 23075 22559
rect 23063 22528 23097 22556
rect 23063 22525 23075 22528
rect 23017 22519 23075 22525
rect 16666 22488 16672 22500
rect 16627 22460 16672 22488
rect 16666 22448 16672 22460
rect 16724 22448 16730 22500
rect 22373 22491 22431 22497
rect 18156 22460 18828 22488
rect 18156 22432 18184 22460
rect 13081 22423 13139 22429
rect 13081 22389 13093 22423
rect 13127 22420 13139 22423
rect 13998 22420 14004 22432
rect 13127 22392 14004 22420
rect 13127 22389 13139 22392
rect 13081 22383 13139 22389
rect 13998 22380 14004 22392
rect 14056 22380 14062 22432
rect 14918 22380 14924 22432
rect 14976 22420 14982 22432
rect 15013 22423 15071 22429
rect 15013 22420 15025 22423
rect 14976 22392 15025 22420
rect 14976 22380 14982 22392
rect 15013 22389 15025 22392
rect 15059 22389 15071 22423
rect 15013 22383 15071 22389
rect 15194 22380 15200 22432
rect 15252 22420 15258 22432
rect 15841 22423 15899 22429
rect 15841 22420 15853 22423
rect 15252 22392 15853 22420
rect 15252 22380 15258 22392
rect 15841 22389 15853 22392
rect 15887 22389 15899 22423
rect 17678 22420 17684 22432
rect 17639 22392 17684 22420
rect 15841 22383 15899 22389
rect 17678 22380 17684 22392
rect 17736 22380 17742 22432
rect 18138 22420 18144 22432
rect 18099 22392 18144 22420
rect 18138 22380 18144 22392
rect 18196 22380 18202 22432
rect 18598 22420 18604 22432
rect 18559 22392 18604 22420
rect 18598 22380 18604 22392
rect 18656 22380 18662 22432
rect 18800 22429 18828 22460
rect 22373 22457 22385 22491
rect 22419 22488 22431 22491
rect 23032 22488 23060 22519
rect 23308 22497 23336 22596
rect 24765 22593 24777 22596
rect 24811 22593 24823 22627
rect 27430 22624 27436 22636
rect 27391 22596 27436 22624
rect 24765 22587 24823 22593
rect 27430 22584 27436 22596
rect 27488 22584 27494 22636
rect 29564 22633 29592 22664
rect 30926 22652 30932 22664
rect 30984 22652 30990 22704
rect 34514 22652 34520 22704
rect 34572 22692 34578 22704
rect 35130 22695 35188 22701
rect 35130 22692 35142 22695
rect 34572 22664 35142 22692
rect 34572 22652 34578 22664
rect 35130 22661 35142 22664
rect 35176 22661 35188 22695
rect 35130 22655 35188 22661
rect 29549 22627 29607 22633
rect 29549 22593 29561 22627
rect 29595 22593 29607 22627
rect 29730 22624 29736 22636
rect 29691 22596 29736 22624
rect 29549 22587 29607 22593
rect 29730 22584 29736 22596
rect 29788 22584 29794 22636
rect 30006 22584 30012 22636
rect 30064 22624 30070 22636
rect 30282 22624 30288 22636
rect 30064 22596 30288 22624
rect 30064 22584 30070 22596
rect 30282 22584 30288 22596
rect 30340 22624 30346 22636
rect 30745 22627 30803 22633
rect 30745 22624 30757 22627
rect 30340 22596 30757 22624
rect 30340 22584 30346 22596
rect 30745 22593 30757 22596
rect 30791 22593 30803 22627
rect 30745 22587 30803 22593
rect 32950 22584 32956 22636
rect 33008 22624 33014 22636
rect 33689 22627 33747 22633
rect 33689 22624 33701 22627
rect 33008 22596 33701 22624
rect 33008 22584 33014 22596
rect 33689 22593 33701 22596
rect 33735 22593 33747 22627
rect 34606 22624 34612 22636
rect 33689 22587 33747 22593
rect 33796 22596 34612 22624
rect 30466 22556 30472 22568
rect 30427 22528 30472 22556
rect 30466 22516 30472 22528
rect 30524 22516 30530 22568
rect 33045 22559 33103 22565
rect 33045 22525 33057 22559
rect 33091 22556 33103 22559
rect 33505 22559 33563 22565
rect 33505 22556 33517 22559
rect 33091 22528 33517 22556
rect 33091 22525 33103 22528
rect 33045 22519 33103 22525
rect 33505 22525 33517 22528
rect 33551 22556 33563 22559
rect 33796 22556 33824 22596
rect 34606 22584 34612 22596
rect 34664 22584 34670 22636
rect 34790 22556 34796 22568
rect 33551 22528 33824 22556
rect 34532 22528 34796 22556
rect 33551 22525 33563 22528
rect 33505 22519 33563 22525
rect 23293 22491 23351 22497
rect 22419 22460 23244 22488
rect 22419 22457 22431 22460
rect 22373 22451 22431 22457
rect 18785 22423 18843 22429
rect 18785 22389 18797 22423
rect 18831 22389 18843 22423
rect 18785 22383 18843 22389
rect 19426 22380 19432 22432
rect 19484 22420 19490 22432
rect 19705 22423 19763 22429
rect 19705 22420 19717 22423
rect 19484 22392 19717 22420
rect 19484 22380 19490 22392
rect 19705 22389 19717 22392
rect 19751 22389 19763 22423
rect 19705 22383 19763 22389
rect 20346 22380 20352 22432
rect 20404 22420 20410 22432
rect 20625 22423 20683 22429
rect 20625 22420 20637 22423
rect 20404 22392 20637 22420
rect 20404 22380 20410 22392
rect 20625 22389 20637 22392
rect 20671 22389 20683 22423
rect 23106 22420 23112 22432
rect 23067 22392 23112 22420
rect 20625 22383 20683 22389
rect 23106 22380 23112 22392
rect 23164 22380 23170 22432
rect 23216 22420 23244 22460
rect 23293 22457 23305 22491
rect 23339 22457 23351 22491
rect 23293 22451 23351 22457
rect 27617 22491 27675 22497
rect 27617 22457 27629 22491
rect 27663 22488 27675 22491
rect 30742 22488 30748 22500
rect 27663 22460 30748 22488
rect 27663 22457 27675 22460
rect 27617 22451 27675 22457
rect 30742 22448 30748 22460
rect 30800 22488 30806 22500
rect 33778 22488 33784 22500
rect 30800 22460 33784 22488
rect 30800 22448 30806 22460
rect 33778 22448 33784 22460
rect 33836 22448 33842 22500
rect 34532 22432 34560 22528
rect 34790 22516 34796 22528
rect 34848 22556 34854 22568
rect 34885 22559 34943 22565
rect 34885 22556 34897 22559
rect 34848 22528 34897 22556
rect 34848 22516 34854 22528
rect 34885 22525 34897 22528
rect 34931 22525 34943 22559
rect 34885 22519 34943 22525
rect 23474 22420 23480 22432
rect 23216 22392 23480 22420
rect 23474 22380 23480 22392
rect 23532 22380 23538 22432
rect 24949 22423 25007 22429
rect 24949 22389 24961 22423
rect 24995 22420 25007 22423
rect 27522 22420 27528 22432
rect 24995 22392 27528 22420
rect 24995 22389 25007 22392
rect 24949 22383 25007 22389
rect 27522 22380 27528 22392
rect 27580 22380 27586 22432
rect 28166 22380 28172 22432
rect 28224 22420 28230 22432
rect 28997 22423 29055 22429
rect 28997 22420 29009 22423
rect 28224 22392 29009 22420
rect 28224 22380 28230 22392
rect 28997 22389 29009 22392
rect 29043 22420 29055 22423
rect 30006 22420 30012 22432
rect 29043 22392 30012 22420
rect 29043 22389 29055 22392
rect 28997 22383 29055 22389
rect 30006 22380 30012 22392
rect 30064 22380 30070 22432
rect 34425 22423 34483 22429
rect 34425 22389 34437 22423
rect 34471 22420 34483 22423
rect 34514 22420 34520 22432
rect 34471 22392 34520 22420
rect 34471 22389 34483 22392
rect 34425 22383 34483 22389
rect 34514 22380 34520 22392
rect 34572 22380 34578 22432
rect 36262 22420 36268 22432
rect 36223 22392 36268 22420
rect 36262 22380 36268 22392
rect 36320 22380 36326 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 4249 22219 4307 22225
rect 4249 22185 4261 22219
rect 4295 22185 4307 22219
rect 4249 22179 4307 22185
rect 4433 22219 4491 22225
rect 4433 22185 4445 22219
rect 4479 22216 4491 22219
rect 5258 22216 5264 22228
rect 4479 22188 5264 22216
rect 4479 22185 4491 22188
rect 4433 22179 4491 22185
rect 4264 22148 4292 22179
rect 5258 22176 5264 22188
rect 5316 22176 5322 22228
rect 6638 22176 6644 22228
rect 6696 22216 6702 22228
rect 7374 22216 7380 22228
rect 6696 22188 7380 22216
rect 6696 22176 6702 22188
rect 7374 22176 7380 22188
rect 7432 22176 7438 22228
rect 9398 22176 9404 22228
rect 9456 22216 9462 22228
rect 10137 22219 10195 22225
rect 10137 22216 10149 22219
rect 9456 22188 10149 22216
rect 9456 22176 9462 22188
rect 10137 22185 10149 22188
rect 10183 22185 10195 22219
rect 10137 22179 10195 22185
rect 29549 22219 29607 22225
rect 29549 22185 29561 22219
rect 29595 22216 29607 22219
rect 29730 22216 29736 22228
rect 29595 22188 29736 22216
rect 29595 22185 29607 22188
rect 29549 22179 29607 22185
rect 29730 22176 29736 22188
rect 29788 22176 29794 22228
rect 4798 22148 4804 22160
rect 4264 22120 4804 22148
rect 4798 22108 4804 22120
rect 4856 22108 4862 22160
rect 11072 22120 11468 22148
rect 4157 22083 4215 22089
rect 4157 22049 4169 22083
rect 4203 22080 4215 22083
rect 4614 22080 4620 22092
rect 4203 22052 4620 22080
rect 4203 22049 4215 22052
rect 4157 22043 4215 22049
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 4816 22080 4844 22108
rect 5905 22083 5963 22089
rect 5905 22080 5917 22083
rect 4816 22052 5917 22080
rect 5905 22049 5917 22052
rect 5951 22049 5963 22083
rect 5905 22043 5963 22049
rect 8386 22040 8392 22092
rect 8444 22080 8450 22092
rect 9033 22083 9091 22089
rect 9033 22080 9045 22083
rect 8444 22052 9045 22080
rect 8444 22040 8450 22052
rect 9033 22049 9045 22052
rect 9079 22080 9091 22083
rect 10321 22083 10379 22089
rect 10321 22080 10333 22083
rect 9079 22052 10333 22080
rect 9079 22049 9091 22052
rect 9033 22043 9091 22049
rect 10321 22049 10333 22052
rect 10367 22080 10379 22083
rect 11072 22080 11100 22120
rect 11440 22092 11468 22120
rect 12526 22108 12532 22160
rect 12584 22148 12590 22160
rect 15286 22148 15292 22160
rect 12584 22120 15292 22148
rect 12584 22108 12590 22120
rect 15286 22108 15292 22120
rect 15344 22148 15350 22160
rect 15344 22120 15424 22148
rect 15344 22108 15350 22120
rect 10367 22052 11100 22080
rect 11149 22083 11207 22089
rect 10367 22049 10379 22052
rect 10321 22043 10379 22049
rect 11149 22049 11161 22083
rect 11195 22080 11207 22083
rect 11330 22080 11336 22092
rect 11195 22052 11336 22080
rect 11195 22049 11207 22052
rect 11149 22043 11207 22049
rect 11330 22040 11336 22052
rect 11388 22040 11394 22092
rect 11422 22040 11428 22092
rect 11480 22040 11486 22092
rect 12618 22080 12624 22092
rect 12579 22052 12624 22080
rect 12618 22040 12624 22052
rect 12676 22040 12682 22092
rect 14918 22080 14924 22092
rect 14879 22052 14924 22080
rect 14918 22040 14924 22052
rect 14976 22040 14982 22092
rect 15105 22083 15163 22089
rect 15105 22049 15117 22083
rect 15151 22080 15163 22083
rect 15194 22080 15200 22092
rect 15151 22052 15200 22080
rect 15151 22049 15163 22052
rect 15105 22043 15163 22049
rect 15194 22040 15200 22052
rect 15252 22040 15258 22092
rect 15396 22089 15424 22120
rect 15381 22083 15439 22089
rect 15381 22049 15393 22083
rect 15427 22080 15439 22083
rect 15427 22052 15461 22080
rect 15427 22049 15439 22052
rect 15381 22043 15439 22049
rect 18046 22040 18052 22092
rect 18104 22080 18110 22092
rect 18414 22080 18420 22092
rect 18104 22052 18420 22080
rect 18104 22040 18110 22052
rect 18414 22040 18420 22052
rect 18472 22040 18478 22092
rect 20346 22080 20352 22092
rect 20307 22052 20352 22080
rect 20346 22040 20352 22052
rect 20404 22040 20410 22092
rect 20438 22040 20444 22092
rect 20496 22080 20502 22092
rect 20717 22083 20775 22089
rect 20717 22080 20729 22083
rect 20496 22052 20729 22080
rect 20496 22040 20502 22052
rect 20717 22049 20729 22052
rect 20763 22049 20775 22083
rect 27614 22080 27620 22092
rect 27575 22052 27620 22080
rect 20717 22043 20775 22049
rect 27614 22040 27620 22052
rect 27672 22040 27678 22092
rect 30193 22083 30251 22089
rect 30193 22049 30205 22083
rect 30239 22080 30251 22083
rect 31018 22080 31024 22092
rect 30239 22052 31024 22080
rect 30239 22049 30251 22052
rect 30193 22043 30251 22049
rect 31018 22040 31024 22052
rect 31076 22040 31082 22092
rect 33045 22083 33103 22089
rect 33045 22080 33057 22083
rect 32140 22052 33057 22080
rect 32140 22024 32168 22052
rect 33045 22049 33057 22052
rect 33091 22080 33103 22083
rect 34514 22080 34520 22092
rect 33091 22052 34520 22080
rect 33091 22049 33103 22052
rect 33045 22043 33103 22049
rect 34514 22040 34520 22052
rect 34572 22080 34578 22092
rect 34572 22052 35848 22080
rect 34572 22040 34578 22052
rect 35820 22024 35848 22052
rect 2682 22012 2688 22024
rect 2643 21984 2688 22012
rect 2682 21972 2688 21984
rect 2740 21972 2746 22024
rect 4246 22012 4252 22024
rect 4207 21984 4252 22012
rect 4246 21972 4252 21984
rect 4304 21972 4310 22024
rect 4982 22012 4988 22024
rect 4943 21984 4988 22012
rect 4982 21972 4988 21984
rect 5040 21972 5046 22024
rect 5629 22015 5687 22021
rect 5629 21981 5641 22015
rect 5675 22012 5687 22015
rect 5810 22012 5816 22024
rect 5675 21984 5816 22012
rect 5675 21981 5687 21984
rect 5629 21975 5687 21981
rect 5810 21972 5816 21984
rect 5868 21972 5874 22024
rect 6917 22015 6975 22021
rect 6917 21981 6929 22015
rect 6963 22012 6975 22015
rect 7098 22012 7104 22024
rect 6963 21984 7104 22012
rect 6963 21981 6975 21984
rect 6917 21975 6975 21981
rect 7098 21972 7104 21984
rect 7156 21972 7162 22024
rect 7650 22012 7656 22024
rect 7611 21984 7656 22012
rect 7650 21972 7656 21984
rect 7708 21972 7714 22024
rect 9493 22015 9551 22021
rect 9493 21981 9505 22015
rect 9539 21981 9551 22015
rect 9493 21975 9551 21981
rect 3973 21947 4031 21953
rect 3973 21913 3985 21947
rect 4019 21944 4031 21947
rect 4706 21944 4712 21956
rect 4019 21916 4712 21944
rect 4019 21913 4031 21916
rect 3973 21907 4031 21913
rect 4706 21904 4712 21916
rect 4764 21904 4770 21956
rect 5828 21944 5856 21972
rect 9508 21944 9536 21975
rect 9582 21972 9588 22024
rect 9640 22012 9646 22024
rect 10413 22015 10471 22021
rect 10413 22012 10425 22015
rect 9640 21984 10425 22012
rect 9640 21972 9646 21984
rect 10413 21981 10425 21984
rect 10459 21981 10471 22015
rect 19705 22015 19763 22021
rect 10413 21975 10471 21981
rect 12912 21984 13124 22012
rect 10137 21947 10195 21953
rect 5828 21916 7880 21944
rect 9508 21916 9904 21944
rect 7852 21888 7880 21916
rect 9876 21888 9904 21916
rect 10137 21913 10149 21947
rect 10183 21944 10195 21947
rect 11330 21944 11336 21956
rect 10183 21916 11192 21944
rect 11291 21916 11336 21944
rect 10183 21913 10195 21916
rect 10137 21907 10195 21913
rect 4614 21836 4620 21888
rect 4672 21876 4678 21888
rect 5169 21879 5227 21885
rect 5169 21876 5181 21879
rect 4672 21848 5181 21876
rect 4672 21836 4678 21848
rect 5169 21845 5181 21848
rect 5215 21845 5227 21879
rect 5169 21839 5227 21845
rect 7101 21879 7159 21885
rect 7101 21845 7113 21879
rect 7147 21876 7159 21879
rect 7374 21876 7380 21888
rect 7147 21848 7380 21876
rect 7147 21845 7159 21848
rect 7101 21839 7159 21845
rect 7374 21836 7380 21848
rect 7432 21836 7438 21888
rect 7834 21876 7840 21888
rect 7747 21848 7840 21876
rect 7834 21836 7840 21848
rect 7892 21836 7898 21888
rect 9677 21879 9735 21885
rect 9677 21845 9689 21879
rect 9723 21876 9735 21879
rect 9766 21876 9772 21888
rect 9723 21848 9772 21876
rect 9723 21845 9735 21848
rect 9677 21839 9735 21845
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 9858 21836 9864 21888
rect 9916 21836 9922 21888
rect 10594 21876 10600 21888
rect 10555 21848 10600 21876
rect 10594 21836 10600 21848
rect 10652 21836 10658 21888
rect 11164 21876 11192 21916
rect 11330 21904 11336 21916
rect 11388 21904 11394 21956
rect 11422 21904 11428 21956
rect 11480 21944 11486 21956
rect 12912 21944 12940 21984
rect 11480 21916 12940 21944
rect 13096 21944 13124 21984
rect 17236 21984 18368 22012
rect 17236 21944 17264 21984
rect 13096 21916 17264 21944
rect 17589 21947 17647 21953
rect 11480 21904 11486 21916
rect 17589 21913 17601 21947
rect 17635 21944 17647 21947
rect 18046 21944 18052 21956
rect 17635 21916 18052 21944
rect 17635 21913 17647 21916
rect 17589 21907 17647 21913
rect 18046 21904 18052 21916
rect 18104 21944 18110 21956
rect 18141 21947 18199 21953
rect 18141 21944 18153 21947
rect 18104 21916 18153 21944
rect 18104 21904 18110 21916
rect 18141 21913 18153 21916
rect 18187 21913 18199 21947
rect 18141 21907 18199 21913
rect 13538 21876 13544 21888
rect 11164 21848 13544 21876
rect 13538 21836 13544 21848
rect 13596 21836 13602 21888
rect 13814 21836 13820 21888
rect 13872 21876 13878 21888
rect 15102 21876 15108 21888
rect 13872 21848 15108 21876
rect 13872 21836 13878 21848
rect 15102 21836 15108 21848
rect 15160 21836 15166 21888
rect 18230 21876 18236 21888
rect 18191 21848 18236 21876
rect 18230 21836 18236 21848
rect 18288 21836 18294 21888
rect 18340 21876 18368 21984
rect 19705 21981 19717 22015
rect 19751 22012 19763 22015
rect 20165 22015 20223 22021
rect 20165 22012 20177 22015
rect 19751 21984 20177 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 20165 21981 20177 21984
rect 20211 21981 20223 22015
rect 23566 22012 23572 22024
rect 23527 21984 23572 22012
rect 20165 21975 20223 21981
rect 23566 21972 23572 21984
rect 23624 21972 23630 22024
rect 27801 22015 27859 22021
rect 27801 21981 27813 22015
rect 27847 22012 27859 22015
rect 30926 22012 30932 22024
rect 27847 21984 30932 22012
rect 27847 21981 27859 21984
rect 27801 21975 27859 21981
rect 30926 21972 30932 21984
rect 30984 21972 30990 22024
rect 31113 22015 31171 22021
rect 31113 21981 31125 22015
rect 31159 22012 31171 22015
rect 32122 22012 32128 22024
rect 31159 21984 32128 22012
rect 31159 21981 31171 21984
rect 31113 21975 31171 21981
rect 32122 21972 32128 21984
rect 32180 21972 32186 22024
rect 33686 21972 33692 22024
rect 33744 22012 33750 22024
rect 33781 22015 33839 22021
rect 33781 22012 33793 22015
rect 33744 21984 33793 22012
rect 33744 21972 33750 21984
rect 33781 21981 33793 21984
rect 33827 21981 33839 22015
rect 33781 21975 33839 21981
rect 34149 22015 34207 22021
rect 34149 21981 34161 22015
rect 34195 22012 34207 22015
rect 35253 22015 35311 22021
rect 35253 22012 35265 22015
rect 34195 21984 35265 22012
rect 34195 21981 34207 21984
rect 34149 21975 34207 21981
rect 35253 21981 35265 21984
rect 35299 21981 35311 22015
rect 35253 21975 35311 21981
rect 35802 21972 35808 22024
rect 35860 22012 35866 22024
rect 36081 22015 36139 22021
rect 36081 22012 36093 22015
rect 35860 21984 36093 22012
rect 35860 21972 35866 21984
rect 36081 21981 36093 21984
rect 36127 21981 36139 22015
rect 36081 21975 36139 21981
rect 24946 21944 24952 21956
rect 22066 21916 24952 21944
rect 22066 21876 22094 21916
rect 24946 21904 24952 21916
rect 25004 21904 25010 21956
rect 25958 21944 25964 21956
rect 25919 21916 25964 21944
rect 25958 21904 25964 21916
rect 26016 21904 26022 21956
rect 31380 21947 31438 21953
rect 31380 21913 31392 21947
rect 31426 21944 31438 21947
rect 31478 21944 31484 21956
rect 31426 21916 31484 21944
rect 31426 21913 31438 21916
rect 31380 21907 31438 21913
rect 31478 21904 31484 21916
rect 31536 21904 31542 21956
rect 33962 21944 33968 21956
rect 33923 21916 33968 21944
rect 33962 21904 33968 21916
rect 34020 21904 34026 21956
rect 36326 21947 36384 21953
rect 36326 21944 36338 21947
rect 35452 21916 36338 21944
rect 22462 21876 22468 21888
rect 18340 21848 22094 21876
rect 22423 21848 22468 21876
rect 22462 21836 22468 21848
rect 22520 21836 22526 21888
rect 28997 21879 29055 21885
rect 28997 21845 29009 21879
rect 29043 21876 29055 21879
rect 29638 21876 29644 21888
rect 29043 21848 29644 21876
rect 29043 21845 29055 21848
rect 28997 21839 29055 21845
rect 29638 21836 29644 21848
rect 29696 21876 29702 21888
rect 29917 21879 29975 21885
rect 29917 21876 29929 21879
rect 29696 21848 29929 21876
rect 29696 21836 29702 21848
rect 29917 21845 29929 21848
rect 29963 21845 29975 21879
rect 29917 21839 29975 21845
rect 30009 21879 30067 21885
rect 30009 21845 30021 21879
rect 30055 21876 30067 21879
rect 31754 21876 31760 21888
rect 30055 21848 31760 21876
rect 30055 21845 30067 21848
rect 30009 21839 30067 21845
rect 31754 21836 31760 21848
rect 31812 21836 31818 21888
rect 31938 21836 31944 21888
rect 31996 21876 32002 21888
rect 32306 21876 32312 21888
rect 31996 21848 32312 21876
rect 31996 21836 32002 21848
rect 32306 21836 32312 21848
rect 32364 21876 32370 21888
rect 35452 21885 35480 21916
rect 36326 21913 36338 21916
rect 36372 21913 36384 21947
rect 36326 21907 36384 21913
rect 32493 21879 32551 21885
rect 32493 21876 32505 21879
rect 32364 21848 32505 21876
rect 32364 21836 32370 21848
rect 32493 21845 32505 21848
rect 32539 21845 32551 21879
rect 32493 21839 32551 21845
rect 35437 21879 35495 21885
rect 35437 21845 35449 21879
rect 35483 21845 35495 21879
rect 35437 21839 35495 21845
rect 36630 21836 36636 21888
rect 36688 21876 36694 21888
rect 37461 21879 37519 21885
rect 37461 21876 37473 21879
rect 36688 21848 37473 21876
rect 36688 21836 36694 21848
rect 37461 21845 37473 21848
rect 37507 21845 37519 21879
rect 37461 21839 37519 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 4154 21632 4160 21684
rect 4212 21672 4218 21684
rect 6825 21675 6883 21681
rect 4212 21644 6684 21672
rect 4212 21632 4218 21644
rect 2869 21607 2927 21613
rect 2869 21573 2881 21607
rect 2915 21604 2927 21607
rect 5074 21604 5080 21616
rect 2915 21576 5080 21604
rect 2915 21573 2927 21576
rect 2869 21567 2927 21573
rect 5074 21564 5080 21576
rect 5132 21564 5138 21616
rect 5166 21564 5172 21616
rect 5224 21604 5230 21616
rect 5224 21576 6592 21604
rect 5224 21564 5230 21576
rect 1394 21536 1400 21548
rect 1355 21508 1400 21536
rect 1394 21496 1400 21508
rect 1452 21536 1458 21548
rect 2041 21539 2099 21545
rect 2041 21536 2053 21539
rect 1452 21508 2053 21536
rect 1452 21496 1458 21508
rect 2041 21505 2053 21508
rect 2087 21505 2099 21539
rect 2682 21536 2688 21548
rect 2643 21508 2688 21536
rect 2041 21499 2099 21505
rect 2682 21496 2688 21508
rect 2740 21496 2746 21548
rect 4522 21536 4528 21548
rect 4483 21508 4528 21536
rect 4522 21496 4528 21508
rect 4580 21496 4586 21548
rect 5442 21536 5448 21548
rect 5403 21508 5448 21536
rect 5442 21496 5448 21508
rect 5500 21496 5506 21548
rect 6564 21545 6592 21576
rect 6656 21545 6684 21644
rect 6825 21641 6837 21675
rect 6871 21641 6883 21675
rect 6825 21635 6883 21641
rect 6365 21539 6423 21545
rect 6365 21505 6377 21539
rect 6411 21505 6423 21539
rect 6365 21499 6423 21505
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21505 6699 21539
rect 6840 21536 6868 21635
rect 9766 21632 9772 21684
rect 9824 21672 9830 21684
rect 9950 21672 9956 21684
rect 9824 21644 9956 21672
rect 9824 21632 9830 21644
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 10226 21632 10232 21684
rect 10284 21672 10290 21684
rect 10686 21672 10692 21684
rect 10284 21644 10692 21672
rect 10284 21632 10290 21644
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 13538 21632 13544 21684
rect 13596 21672 13602 21684
rect 22462 21672 22468 21684
rect 13596 21644 22468 21672
rect 13596 21632 13602 21644
rect 22462 21632 22468 21644
rect 22520 21632 22526 21684
rect 30926 21632 30932 21684
rect 30984 21672 30990 21684
rect 31938 21672 31944 21684
rect 30984 21644 31944 21672
rect 30984 21632 30990 21644
rect 31938 21632 31944 21644
rect 31996 21632 32002 21684
rect 32122 21672 32128 21684
rect 32083 21644 32128 21672
rect 32122 21632 32128 21644
rect 32180 21632 32186 21684
rect 35802 21632 35808 21684
rect 35860 21672 35866 21684
rect 35897 21675 35955 21681
rect 35897 21672 35909 21675
rect 35860 21644 35909 21672
rect 35860 21632 35866 21644
rect 35897 21641 35909 21644
rect 35943 21641 35955 21675
rect 38010 21672 38016 21684
rect 37971 21644 38016 21672
rect 35897 21635 35955 21641
rect 38010 21632 38016 21644
rect 38068 21632 38074 21684
rect 11698 21604 11704 21616
rect 11659 21576 11704 21604
rect 11698 21564 11704 21576
rect 11756 21564 11762 21616
rect 12434 21564 12440 21616
rect 12492 21604 12498 21616
rect 18230 21604 18236 21616
rect 12492 21576 18236 21604
rect 12492 21564 12498 21576
rect 18230 21564 18236 21576
rect 18288 21564 18294 21616
rect 19426 21564 19432 21616
rect 19484 21604 19490 21616
rect 19613 21607 19671 21613
rect 19613 21604 19625 21607
rect 19484 21576 19625 21604
rect 19484 21564 19490 21576
rect 19613 21573 19625 21576
rect 19659 21573 19671 21607
rect 19613 21567 19671 21573
rect 23566 21564 23572 21616
rect 23624 21604 23630 21616
rect 30000 21607 30058 21613
rect 23624 21576 25268 21604
rect 23624 21564 23630 21576
rect 7285 21539 7343 21545
rect 7285 21536 7297 21539
rect 6840 21508 7297 21536
rect 6641 21499 6699 21505
rect 7285 21505 7297 21508
rect 7331 21505 7343 21539
rect 7285 21499 7343 21505
rect 4982 21428 4988 21480
rect 5040 21468 5046 21480
rect 5350 21468 5356 21480
rect 5040 21440 5356 21468
rect 5040 21428 5046 21440
rect 5350 21428 5356 21440
rect 5408 21428 5414 21480
rect 6380 21400 6408 21499
rect 9582 21496 9588 21548
rect 9640 21536 9646 21548
rect 9677 21539 9735 21545
rect 9677 21536 9689 21539
rect 9640 21508 9689 21536
rect 9640 21496 9646 21508
rect 9677 21505 9689 21508
rect 9723 21505 9735 21539
rect 10870 21536 10876 21548
rect 10831 21508 10876 21536
rect 9677 21499 9735 21505
rect 10870 21496 10876 21508
rect 10928 21496 10934 21548
rect 11514 21536 11520 21548
rect 11475 21508 11520 21536
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 13814 21536 13820 21548
rect 13775 21508 13820 21536
rect 13814 21496 13820 21508
rect 13872 21536 13878 21548
rect 13998 21536 14004 21548
rect 13872 21508 14004 21536
rect 13872 21496 13878 21508
rect 13998 21496 14004 21508
rect 14056 21536 14062 21548
rect 14553 21539 14611 21545
rect 14553 21536 14565 21539
rect 14056 21508 14565 21536
rect 14056 21496 14062 21508
rect 14553 21505 14565 21508
rect 14599 21505 14611 21539
rect 14553 21499 14611 21505
rect 17129 21539 17187 21545
rect 17129 21505 17141 21539
rect 17175 21536 17187 21539
rect 17678 21536 17684 21548
rect 17175 21508 17684 21536
rect 17175 21505 17187 21508
rect 17129 21499 17187 21505
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 25240 21545 25268 21576
rect 30000 21573 30012 21607
rect 30046 21604 30058 21607
rect 30098 21604 30104 21616
rect 30046 21576 30104 21604
rect 30046 21573 30058 21576
rect 30000 21567 30058 21573
rect 30098 21564 30104 21576
rect 30156 21564 30162 21616
rect 25225 21539 25283 21545
rect 25225 21505 25237 21539
rect 25271 21505 25283 21539
rect 25958 21536 25964 21548
rect 25919 21508 25964 21536
rect 25225 21499 25283 21505
rect 25958 21496 25964 21508
rect 26016 21496 26022 21548
rect 7374 21428 7380 21480
rect 7432 21468 7438 21480
rect 8941 21471 8999 21477
rect 8941 21468 8953 21471
rect 7432 21440 8953 21468
rect 7432 21428 7438 21440
rect 8941 21437 8953 21440
rect 8987 21468 8999 21471
rect 9401 21471 9459 21477
rect 9401 21468 9413 21471
rect 8987 21440 9413 21468
rect 8987 21437 8999 21440
rect 8941 21431 8999 21437
rect 9401 21437 9413 21440
rect 9447 21468 9459 21471
rect 9950 21468 9956 21480
rect 9447 21440 9956 21468
rect 9447 21437 9459 21440
rect 9401 21431 9459 21437
rect 9950 21428 9956 21440
rect 10008 21428 10014 21480
rect 12526 21468 12532 21480
rect 12487 21440 12532 21468
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 17402 21468 17408 21480
rect 17363 21440 17408 21468
rect 17402 21428 17408 21440
rect 17460 21428 17466 21480
rect 19429 21471 19487 21477
rect 19429 21437 19441 21471
rect 19475 21468 19487 21471
rect 19702 21468 19708 21480
rect 19475 21440 19708 21468
rect 19475 21437 19487 21440
rect 19429 21431 19487 21437
rect 19702 21428 19708 21440
rect 19760 21428 19766 21480
rect 19889 21471 19947 21477
rect 19889 21437 19901 21471
rect 19935 21468 19947 21471
rect 20438 21468 20444 21480
rect 19935 21440 20444 21468
rect 19935 21437 19947 21440
rect 19889 21431 19947 21437
rect 12434 21400 12440 21412
rect 6380 21372 12440 21400
rect 12434 21360 12440 21372
rect 12492 21360 12498 21412
rect 12618 21360 12624 21412
rect 12676 21400 12682 21412
rect 19904 21400 19932 21431
rect 20438 21428 20444 21440
rect 20496 21428 20502 21480
rect 23658 21468 23664 21480
rect 23619 21440 23664 21468
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 25038 21468 25044 21480
rect 24999 21440 25044 21468
rect 25038 21428 25044 21440
rect 25096 21428 25102 21480
rect 29733 21471 29791 21477
rect 29733 21437 29745 21471
rect 29779 21437 29791 21471
rect 29733 21431 29791 21437
rect 12676 21372 19932 21400
rect 12676 21360 12682 21372
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 2498 21332 2504 21344
rect 1627 21304 2504 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 2498 21292 2504 21304
rect 2556 21292 2562 21344
rect 5258 21332 5264 21344
rect 5219 21304 5264 21332
rect 5258 21292 5264 21304
rect 5316 21292 5322 21344
rect 5350 21292 5356 21344
rect 5408 21332 5414 21344
rect 6365 21335 6423 21341
rect 6365 21332 6377 21335
rect 5408 21304 6377 21332
rect 5408 21292 5414 21304
rect 6365 21301 6377 21304
rect 6411 21301 6423 21335
rect 6365 21295 6423 21301
rect 7469 21335 7527 21341
rect 7469 21301 7481 21335
rect 7515 21332 7527 21335
rect 7650 21332 7656 21344
rect 7515 21304 7656 21332
rect 7515 21301 7527 21304
rect 7469 21295 7527 21301
rect 7650 21292 7656 21304
rect 7708 21292 7714 21344
rect 7926 21332 7932 21344
rect 7887 21304 7932 21332
rect 7926 21292 7932 21304
rect 7984 21292 7990 21344
rect 13906 21292 13912 21344
rect 13964 21332 13970 21344
rect 14001 21335 14059 21341
rect 14001 21332 14013 21335
rect 13964 21304 14013 21332
rect 13964 21292 13970 21304
rect 14001 21301 14013 21304
rect 14047 21332 14059 21335
rect 22738 21332 22744 21344
rect 14047 21304 22744 21332
rect 14047 21301 14059 21304
rect 14001 21295 14059 21301
rect 22738 21292 22744 21304
rect 22796 21292 22802 21344
rect 26237 21335 26295 21341
rect 26237 21301 26249 21335
rect 26283 21332 26295 21335
rect 26326 21332 26332 21344
rect 26283 21304 26332 21332
rect 26283 21301 26295 21304
rect 26237 21295 26295 21301
rect 26326 21292 26332 21304
rect 26384 21292 26390 21344
rect 29748 21332 29776 21431
rect 32140 21400 32168 21632
rect 37826 21536 37832 21548
rect 37787 21508 37832 21536
rect 37826 21496 37832 21508
rect 37884 21496 37890 21548
rect 30668 21372 32168 21400
rect 30668 21332 30696 21372
rect 29748 21304 30696 21332
rect 31113 21335 31171 21341
rect 31113 21301 31125 21335
rect 31159 21332 31171 21335
rect 31754 21332 31760 21344
rect 31159 21304 31760 21332
rect 31159 21301 31171 21304
rect 31113 21295 31171 21301
rect 31754 21292 31760 21304
rect 31812 21292 31818 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 4617 21131 4675 21137
rect 4617 21097 4629 21131
rect 4663 21128 4675 21131
rect 4798 21128 4804 21140
rect 4663 21100 4804 21128
rect 4663 21097 4675 21100
rect 4617 21091 4675 21097
rect 4798 21088 4804 21100
rect 4856 21128 4862 21140
rect 5350 21128 5356 21140
rect 4856 21100 5356 21128
rect 4856 21088 4862 21100
rect 5350 21088 5356 21100
rect 5408 21088 5414 21140
rect 7834 21088 7840 21140
rect 7892 21128 7898 21140
rect 8297 21131 8355 21137
rect 8297 21128 8309 21131
rect 7892 21100 8309 21128
rect 7892 21088 7898 21100
rect 8297 21097 8309 21100
rect 8343 21097 8355 21131
rect 8297 21091 8355 21097
rect 11241 21131 11299 21137
rect 11241 21097 11253 21131
rect 11287 21128 11299 21131
rect 11882 21128 11888 21140
rect 11287 21100 11888 21128
rect 11287 21097 11299 21100
rect 11241 21091 11299 21097
rect 5166 21060 5172 21072
rect 4540 21032 5172 21060
rect 4540 21001 4568 21032
rect 5166 21020 5172 21032
rect 5224 21020 5230 21072
rect 4525 20995 4583 21001
rect 4525 20961 4537 20995
rect 4571 20961 4583 20995
rect 5258 20992 5264 21004
rect 5219 20964 5264 20992
rect 4525 20955 4583 20961
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5534 20992 5540 21004
rect 5495 20964 5540 20992
rect 5534 20952 5540 20964
rect 5592 20952 5598 21004
rect 8312 20992 8340 21091
rect 11882 21088 11888 21100
rect 11940 21088 11946 21140
rect 12342 21128 12348 21140
rect 12303 21100 12348 21128
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 19702 21128 19708 21140
rect 19663 21100 19708 21128
rect 19702 21088 19708 21100
rect 19760 21088 19766 21140
rect 24394 21128 24400 21140
rect 24355 21100 24400 21128
rect 24394 21088 24400 21100
rect 24452 21088 24458 21140
rect 25038 21088 25044 21140
rect 25096 21128 25102 21140
rect 25317 21131 25375 21137
rect 25317 21128 25329 21131
rect 25096 21100 25329 21128
rect 25096 21088 25102 21100
rect 25317 21097 25329 21100
rect 25363 21097 25375 21131
rect 25317 21091 25375 21097
rect 26326 21088 26332 21140
rect 26384 21128 26390 21140
rect 29546 21128 29552 21140
rect 26384 21100 29552 21128
rect 26384 21088 26390 21100
rect 29546 21088 29552 21100
rect 29604 21128 29610 21140
rect 29914 21128 29920 21140
rect 29604 21100 29920 21128
rect 29604 21088 29610 21100
rect 29914 21088 29920 21100
rect 29972 21088 29978 21140
rect 30469 21131 30527 21137
rect 30469 21097 30481 21131
rect 30515 21128 30527 21131
rect 30834 21128 30840 21140
rect 30515 21100 30840 21128
rect 30515 21097 30527 21100
rect 30469 21091 30527 21097
rect 30834 21088 30840 21100
rect 30892 21088 30898 21140
rect 9950 21020 9956 21072
rect 10008 21060 10014 21072
rect 24302 21060 24308 21072
rect 10008 21032 24308 21060
rect 10008 21020 10014 21032
rect 24302 21020 24308 21032
rect 24360 21020 24366 21072
rect 9309 20995 9367 21001
rect 9309 20992 9321 20995
rect 8312 20964 9321 20992
rect 9309 20961 9321 20964
rect 9355 20961 9367 20995
rect 9309 20955 9367 20961
rect 9398 20952 9404 21004
rect 9456 20992 9462 21004
rect 9585 20995 9643 21001
rect 9585 20992 9597 20995
rect 9456 20964 9597 20992
rect 9456 20952 9462 20964
rect 9585 20961 9597 20964
rect 9631 20961 9643 20995
rect 9585 20955 9643 20961
rect 10686 20952 10692 21004
rect 10744 20992 10750 21004
rect 11057 20995 11115 21001
rect 11057 20992 11069 20995
rect 10744 20964 11069 20992
rect 10744 20952 10750 20964
rect 11057 20961 11069 20964
rect 11103 20992 11115 20995
rect 11977 20995 12035 21001
rect 11977 20992 11989 20995
rect 11103 20964 11989 20992
rect 11103 20961 11115 20964
rect 11057 20955 11115 20961
rect 11977 20961 11989 20964
rect 12023 20961 12035 20995
rect 11977 20955 12035 20961
rect 18141 20995 18199 21001
rect 18141 20961 18153 20995
rect 18187 20992 18199 20995
rect 18598 20992 18604 21004
rect 18187 20964 18604 20992
rect 18187 20961 18199 20964
rect 18141 20955 18199 20961
rect 18598 20952 18604 20964
rect 18656 20952 18662 21004
rect 24486 20992 24492 21004
rect 24447 20964 24492 20992
rect 24486 20952 24492 20964
rect 24544 20952 24550 21004
rect 28445 20995 28503 21001
rect 28445 20961 28457 20995
rect 28491 20992 28503 20995
rect 29638 20992 29644 21004
rect 28491 20964 29644 20992
rect 28491 20961 28503 20964
rect 28445 20955 28503 20961
rect 29638 20952 29644 20964
rect 29696 20952 29702 21004
rect 31018 20992 31024 21004
rect 30979 20964 31024 20992
rect 31018 20952 31024 20964
rect 31076 20952 31082 21004
rect 4154 20884 4160 20936
rect 4212 20924 4218 20936
rect 4341 20927 4399 20933
rect 4341 20924 4353 20927
rect 4212 20896 4353 20924
rect 4212 20884 4218 20896
rect 4341 20893 4353 20896
rect 4387 20893 4399 20927
rect 4614 20924 4620 20936
rect 4575 20896 4620 20924
rect 4341 20887 4399 20893
rect 4356 20856 4384 20887
rect 4614 20884 4620 20896
rect 4672 20884 4678 20936
rect 5074 20924 5080 20936
rect 5035 20896 5080 20924
rect 5074 20884 5080 20896
rect 5132 20884 5138 20936
rect 11241 20927 11299 20933
rect 11241 20893 11253 20927
rect 11287 20924 11299 20927
rect 12161 20927 12219 20933
rect 12161 20924 12173 20927
rect 11287 20896 12173 20924
rect 11287 20893 11299 20896
rect 11241 20887 11299 20893
rect 12161 20893 12173 20896
rect 12207 20924 12219 20927
rect 12710 20924 12716 20936
rect 12207 20896 12716 20924
rect 12207 20893 12219 20896
rect 12161 20887 12219 20893
rect 12710 20884 12716 20896
rect 12768 20884 12774 20936
rect 12894 20884 12900 20936
rect 12952 20924 12958 20936
rect 13262 20924 13268 20936
rect 12952 20896 13268 20924
rect 12952 20884 12958 20896
rect 13262 20884 13268 20896
rect 13320 20884 13326 20936
rect 16298 20924 16304 20936
rect 16259 20896 16304 20924
rect 16298 20884 16304 20896
rect 16356 20884 16362 20936
rect 16942 20884 16948 20936
rect 17000 20924 17006 20936
rect 17865 20927 17923 20933
rect 17865 20924 17877 20927
rect 17000 20896 17877 20924
rect 17000 20884 17006 20896
rect 17865 20893 17877 20896
rect 17911 20893 17923 20927
rect 17865 20887 17923 20893
rect 22462 20884 22468 20936
rect 22520 20924 22526 20936
rect 22649 20927 22707 20933
rect 22649 20924 22661 20927
rect 22520 20896 22661 20924
rect 22520 20884 22526 20896
rect 22649 20893 22661 20896
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 22925 20927 22983 20933
rect 22925 20893 22937 20927
rect 22971 20924 22983 20927
rect 23934 20924 23940 20936
rect 22971 20896 23940 20924
rect 22971 20893 22983 20896
rect 22925 20887 22983 20893
rect 23934 20884 23940 20896
rect 23992 20924 23998 20936
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 23992 20896 24409 20924
rect 23992 20884 23998 20896
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 24578 20884 24584 20936
rect 24636 20924 24642 20936
rect 24673 20927 24731 20933
rect 24673 20924 24685 20927
rect 24636 20896 24685 20924
rect 24636 20884 24642 20896
rect 24673 20893 24685 20896
rect 24719 20893 24731 20927
rect 25501 20927 25559 20933
rect 25501 20924 25513 20927
rect 24673 20887 24731 20893
rect 24872 20896 25513 20924
rect 5258 20856 5264 20868
rect 4356 20828 5264 20856
rect 5258 20816 5264 20828
rect 5316 20816 5322 20868
rect 9766 20816 9772 20868
rect 9824 20856 9830 20868
rect 10965 20859 11023 20865
rect 10965 20856 10977 20859
rect 9824 20828 10977 20856
rect 9824 20816 9830 20828
rect 10965 20825 10977 20828
rect 11011 20856 11023 20859
rect 11885 20859 11943 20865
rect 11885 20856 11897 20859
rect 11011 20828 11897 20856
rect 11011 20825 11023 20828
rect 10965 20819 11023 20825
rect 11885 20825 11897 20828
rect 11931 20825 11943 20859
rect 11885 20819 11943 20825
rect 4154 20788 4160 20800
rect 4115 20760 4160 20788
rect 4154 20748 4160 20760
rect 4212 20748 4218 20800
rect 11425 20791 11483 20797
rect 11425 20757 11437 20791
rect 11471 20788 11483 20791
rect 11790 20788 11796 20800
rect 11471 20760 11796 20788
rect 11471 20757 11483 20760
rect 11425 20751 11483 20757
rect 11790 20748 11796 20760
rect 11848 20748 11854 20800
rect 13078 20788 13084 20800
rect 13039 20760 13084 20788
rect 13078 20748 13084 20760
rect 13136 20748 13142 20800
rect 24872 20797 24900 20896
rect 25501 20893 25513 20896
rect 25547 20893 25559 20927
rect 25501 20887 25559 20893
rect 28905 20927 28963 20933
rect 28905 20893 28917 20927
rect 28951 20924 28963 20927
rect 31754 20924 31760 20936
rect 28951 20896 31760 20924
rect 28951 20893 28963 20896
rect 28905 20887 28963 20893
rect 31754 20884 31760 20896
rect 31812 20924 31818 20936
rect 32582 20924 32588 20936
rect 31812 20896 32588 20924
rect 31812 20884 31818 20896
rect 32582 20884 32588 20896
rect 32640 20884 32646 20936
rect 27522 20816 27528 20868
rect 27580 20856 27586 20868
rect 28721 20859 28779 20865
rect 28721 20856 28733 20859
rect 27580 20828 28733 20856
rect 27580 20816 27586 20828
rect 28721 20825 28733 20828
rect 28767 20825 28779 20859
rect 30926 20856 30932 20868
rect 30887 20828 30932 20856
rect 28721 20819 28779 20825
rect 30926 20816 30932 20828
rect 30984 20816 30990 20868
rect 24857 20791 24915 20797
rect 24857 20757 24869 20791
rect 24903 20757 24915 20791
rect 24857 20751 24915 20757
rect 25314 20748 25320 20800
rect 25372 20788 25378 20800
rect 25958 20788 25964 20800
rect 25372 20760 25964 20788
rect 25372 20748 25378 20760
rect 25958 20748 25964 20760
rect 26016 20748 26022 20800
rect 29914 20748 29920 20800
rect 29972 20788 29978 20800
rect 30837 20791 30895 20797
rect 30837 20788 30849 20791
rect 29972 20760 30849 20788
rect 29972 20748 29978 20760
rect 30837 20757 30849 20760
rect 30883 20757 30895 20791
rect 30837 20751 30895 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 5442 20584 5448 20596
rect 5403 20556 5448 20584
rect 5442 20544 5448 20556
rect 5500 20544 5506 20596
rect 11330 20544 11336 20596
rect 11388 20584 11394 20596
rect 11609 20587 11667 20593
rect 11609 20584 11621 20587
rect 11388 20556 11621 20584
rect 11388 20544 11394 20556
rect 11609 20553 11621 20556
rect 11655 20553 11667 20587
rect 12710 20584 12716 20596
rect 12671 20556 12716 20584
rect 11609 20547 11667 20553
rect 12710 20544 12716 20556
rect 12768 20544 12774 20596
rect 14001 20587 14059 20593
rect 14001 20553 14013 20587
rect 14047 20584 14059 20587
rect 24673 20587 24731 20593
rect 14047 20556 22094 20584
rect 14047 20553 14059 20556
rect 14001 20547 14059 20553
rect 4062 20476 4068 20528
rect 4120 20516 4126 20528
rect 5534 20516 5540 20528
rect 4120 20488 5540 20516
rect 4120 20476 4126 20488
rect 5534 20476 5540 20488
rect 5592 20476 5598 20528
rect 7650 20516 7656 20528
rect 7611 20488 7656 20516
rect 7650 20476 7656 20488
rect 7708 20476 7714 20528
rect 1394 20448 1400 20460
rect 1355 20420 1400 20448
rect 1394 20408 1400 20420
rect 1452 20448 1458 20460
rect 2041 20451 2099 20457
rect 2041 20448 2053 20451
rect 1452 20420 2053 20448
rect 1452 20408 1458 20420
rect 2041 20417 2053 20420
rect 2087 20417 2099 20451
rect 2041 20411 2099 20417
rect 3329 20451 3387 20457
rect 3329 20417 3341 20451
rect 3375 20448 3387 20451
rect 4154 20448 4160 20460
rect 3375 20420 4160 20448
rect 3375 20417 3387 20420
rect 3329 20411 3387 20417
rect 4154 20408 4160 20420
rect 4212 20408 4218 20460
rect 4614 20408 4620 20460
rect 4672 20448 4678 20460
rect 4985 20451 5043 20457
rect 4985 20448 4997 20451
rect 4672 20420 4997 20448
rect 4672 20408 4678 20420
rect 4985 20417 4997 20420
rect 5031 20417 5043 20451
rect 5166 20448 5172 20460
rect 5127 20420 5172 20448
rect 4985 20411 5043 20417
rect 5166 20408 5172 20420
rect 5224 20408 5230 20460
rect 5258 20408 5264 20460
rect 5316 20448 5322 20460
rect 11790 20448 11796 20460
rect 5316 20420 5361 20448
rect 11751 20420 11796 20448
rect 5316 20408 5322 20420
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20448 12955 20451
rect 13078 20448 13084 20460
rect 12943 20420 13084 20448
rect 12943 20417 12955 20420
rect 12897 20411 12955 20417
rect 13078 20408 13084 20420
rect 13136 20448 13142 20460
rect 14016 20448 14044 20547
rect 16853 20519 16911 20525
rect 16853 20485 16865 20519
rect 16899 20516 16911 20519
rect 17402 20516 17408 20528
rect 16899 20488 17408 20516
rect 16899 20485 16911 20488
rect 16853 20479 16911 20485
rect 17402 20476 17408 20488
rect 17460 20476 17466 20528
rect 13136 20420 14044 20448
rect 13136 20408 13142 20420
rect 16298 20408 16304 20460
rect 16356 20448 16362 20460
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 16356 20420 16681 20448
rect 16356 20408 16362 20420
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 7469 20383 7527 20389
rect 7469 20349 7481 20383
rect 7515 20380 7527 20383
rect 7926 20380 7932 20392
rect 7515 20352 7932 20380
rect 7515 20349 7527 20352
rect 7469 20343 7527 20349
rect 7926 20340 7932 20352
rect 7984 20340 7990 20392
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20349 8079 20383
rect 8021 20343 8079 20349
rect 5534 20272 5540 20324
rect 5592 20312 5598 20324
rect 8036 20312 8064 20343
rect 14918 20340 14924 20392
rect 14976 20380 14982 20392
rect 17129 20383 17187 20389
rect 17129 20380 17141 20383
rect 14976 20352 17141 20380
rect 14976 20340 14982 20352
rect 17129 20349 17141 20352
rect 17175 20349 17187 20383
rect 22066 20380 22094 20556
rect 24673 20553 24685 20587
rect 24719 20553 24731 20587
rect 24673 20547 24731 20553
rect 26053 20587 26111 20593
rect 26053 20553 26065 20587
rect 26099 20584 26111 20587
rect 27522 20584 27528 20596
rect 26099 20556 27528 20584
rect 26099 20553 26111 20556
rect 26053 20547 26111 20553
rect 23934 20476 23940 20528
rect 23992 20516 23998 20528
rect 24213 20519 24271 20525
rect 24213 20516 24225 20519
rect 23992 20488 24225 20516
rect 23992 20476 23998 20488
rect 24213 20485 24225 20488
rect 24259 20485 24271 20519
rect 24213 20479 24271 20485
rect 24489 20451 24547 20457
rect 24489 20417 24501 20451
rect 24535 20448 24547 20451
rect 24578 20448 24584 20460
rect 24535 20420 24584 20448
rect 24535 20417 24547 20420
rect 24489 20411 24547 20417
rect 24578 20408 24584 20420
rect 24636 20408 24642 20460
rect 24688 20448 24716 20547
rect 27522 20544 27528 20556
rect 27580 20544 27586 20596
rect 25869 20451 25927 20457
rect 25869 20448 25881 20451
rect 24688 20420 25881 20448
rect 25869 20417 25881 20420
rect 25915 20417 25927 20451
rect 25869 20411 25927 20417
rect 23290 20380 23296 20392
rect 22066 20352 23296 20380
rect 17129 20343 17187 20349
rect 23290 20340 23296 20352
rect 23348 20340 23354 20392
rect 24302 20380 24308 20392
rect 23676 20352 24308 20380
rect 5592 20284 8064 20312
rect 5592 20272 5598 20284
rect 1581 20247 1639 20253
rect 1581 20213 1593 20247
rect 1627 20244 1639 20247
rect 2314 20244 2320 20256
rect 1627 20216 2320 20244
rect 1627 20213 1639 20216
rect 1581 20207 1639 20213
rect 2314 20204 2320 20216
rect 2372 20204 2378 20256
rect 2590 20204 2596 20256
rect 2648 20244 2654 20256
rect 3145 20247 3203 20253
rect 3145 20244 3157 20247
rect 2648 20216 3157 20244
rect 2648 20204 2654 20216
rect 3145 20213 3157 20216
rect 3191 20213 3203 20247
rect 3145 20207 3203 20213
rect 5261 20247 5319 20253
rect 5261 20213 5273 20247
rect 5307 20244 5319 20247
rect 5350 20244 5356 20256
rect 5307 20216 5356 20244
rect 5307 20213 5319 20216
rect 5261 20207 5319 20213
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 8036 20244 8064 20284
rect 9674 20272 9680 20324
rect 9732 20312 9738 20324
rect 19610 20312 19616 20324
rect 9732 20284 19616 20312
rect 9732 20272 9738 20284
rect 19610 20272 19616 20284
rect 19668 20312 19674 20324
rect 20073 20315 20131 20321
rect 20073 20312 20085 20315
rect 19668 20284 20085 20312
rect 19668 20272 19674 20284
rect 20073 20281 20085 20284
rect 20119 20281 20131 20315
rect 20073 20275 20131 20281
rect 12618 20244 12624 20256
rect 8036 20216 12624 20244
rect 12618 20204 12624 20216
rect 12676 20204 12682 20256
rect 13262 20204 13268 20256
rect 13320 20244 13326 20256
rect 13357 20247 13415 20253
rect 13357 20244 13369 20247
rect 13320 20216 13369 20244
rect 13320 20204 13326 20216
rect 13357 20213 13369 20216
rect 13403 20213 13415 20247
rect 13357 20207 13415 20213
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 19521 20247 19579 20253
rect 19521 20244 19533 20247
rect 19392 20216 19533 20244
rect 19392 20204 19398 20216
rect 19521 20213 19533 20216
rect 19567 20244 19579 20247
rect 19978 20244 19984 20256
rect 19567 20216 19984 20244
rect 19567 20213 19579 20216
rect 19521 20207 19579 20213
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 23474 20244 23480 20256
rect 22152 20216 23480 20244
rect 22152 20204 22158 20216
rect 23474 20204 23480 20216
rect 23532 20244 23538 20256
rect 23676 20253 23704 20352
rect 24302 20340 24308 20352
rect 24360 20340 24366 20392
rect 23661 20247 23719 20253
rect 23661 20244 23673 20247
rect 23532 20216 23673 20244
rect 23532 20204 23538 20216
rect 23661 20213 23673 20216
rect 23707 20213 23719 20247
rect 24394 20244 24400 20256
rect 24355 20216 24400 20244
rect 23661 20207 23719 20213
rect 24394 20204 24400 20216
rect 24452 20204 24458 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 5074 20000 5080 20052
rect 5132 20040 5138 20052
rect 5169 20043 5227 20049
rect 5169 20040 5181 20043
rect 5132 20012 5181 20040
rect 5132 20000 5138 20012
rect 5169 20009 5181 20012
rect 5215 20009 5227 20043
rect 5169 20003 5227 20009
rect 7834 20000 7840 20052
rect 7892 20040 7898 20052
rect 8021 20043 8079 20049
rect 8021 20040 8033 20043
rect 7892 20012 8033 20040
rect 7892 20000 7898 20012
rect 8021 20009 8033 20012
rect 8067 20009 8079 20043
rect 8021 20003 8079 20009
rect 22925 20043 22983 20049
rect 22925 20009 22937 20043
rect 22971 20040 22983 20043
rect 24394 20040 24400 20052
rect 22971 20012 24400 20040
rect 22971 20009 22983 20012
rect 22925 20003 22983 20009
rect 24394 20000 24400 20012
rect 24452 20000 24458 20052
rect 35986 20040 35992 20052
rect 35947 20012 35992 20040
rect 35986 20000 35992 20012
rect 36044 20000 36050 20052
rect 36998 20000 37004 20052
rect 37056 20040 37062 20052
rect 37093 20043 37151 20049
rect 37093 20040 37105 20043
rect 37056 20012 37105 20040
rect 37056 20000 37062 20012
rect 37093 20009 37105 20012
rect 37139 20009 37151 20043
rect 37093 20003 37151 20009
rect 7561 19907 7619 19913
rect 7561 19873 7573 19907
rect 7607 19904 7619 19907
rect 7852 19904 7880 20000
rect 12069 19975 12127 19981
rect 12069 19941 12081 19975
rect 12115 19972 12127 19975
rect 13906 19972 13912 19984
rect 12115 19944 13912 19972
rect 12115 19941 12127 19944
rect 12069 19935 12127 19941
rect 12544 19913 12572 19944
rect 13906 19932 13912 19944
rect 13964 19932 13970 19984
rect 20898 19932 20904 19984
rect 20956 19972 20962 19984
rect 27430 19972 27436 19984
rect 20956 19944 27436 19972
rect 20956 19932 20962 19944
rect 27430 19932 27436 19944
rect 27488 19932 27494 19984
rect 7607 19876 7880 19904
rect 12529 19907 12587 19913
rect 7607 19873 7619 19876
rect 7561 19867 7619 19873
rect 12529 19873 12541 19907
rect 12575 19873 12587 19907
rect 12529 19867 12587 19873
rect 12618 19864 12624 19916
rect 12676 19904 12682 19916
rect 14918 19904 14924 19916
rect 12676 19876 14924 19904
rect 12676 19864 12682 19876
rect 14918 19864 14924 19876
rect 14976 19864 14982 19916
rect 16942 19904 16948 19916
rect 16903 19876 16948 19904
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 17954 19904 17960 19916
rect 17915 19876 17960 19904
rect 17954 19864 17960 19876
rect 18012 19864 18018 19916
rect 24302 19864 24308 19916
rect 24360 19904 24366 19916
rect 24489 19907 24547 19913
rect 24489 19904 24501 19907
rect 24360 19876 24501 19904
rect 24360 19864 24366 19876
rect 24489 19873 24501 19876
rect 24535 19904 24547 19907
rect 25317 19907 25375 19913
rect 25317 19904 25329 19907
rect 24535 19876 25329 19904
rect 24535 19873 24547 19876
rect 24489 19867 24547 19873
rect 25317 19873 25329 19876
rect 25363 19873 25375 19907
rect 25317 19867 25375 19873
rect 36449 19907 36507 19913
rect 36449 19873 36461 19907
rect 36495 19904 36507 19907
rect 36814 19904 36820 19916
rect 36495 19876 36820 19904
rect 36495 19873 36507 19876
rect 36449 19867 36507 19873
rect 36814 19864 36820 19876
rect 36872 19904 36878 19916
rect 37553 19907 37611 19913
rect 37553 19904 37565 19907
rect 36872 19876 37565 19904
rect 36872 19864 36878 19876
rect 37553 19873 37565 19876
rect 37599 19873 37611 19907
rect 37553 19867 37611 19873
rect 37645 19907 37703 19913
rect 37645 19873 37657 19907
rect 37691 19873 37703 19907
rect 37645 19867 37703 19873
rect 2406 19836 2412 19848
rect 2367 19808 2412 19836
rect 2406 19796 2412 19808
rect 2464 19796 2470 19848
rect 7282 19836 7288 19848
rect 7243 19808 7288 19836
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 12805 19839 12863 19845
rect 12805 19805 12817 19839
rect 12851 19805 12863 19839
rect 14458 19836 14464 19848
rect 14419 19808 14464 19836
rect 12805 19799 12863 19805
rect 11882 19728 11888 19780
rect 11940 19768 11946 19780
rect 12342 19768 12348 19780
rect 11940 19740 12348 19768
rect 11940 19728 11946 19740
rect 12342 19728 12348 19740
rect 12400 19768 12406 19780
rect 12820 19768 12848 19799
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 16758 19836 16764 19848
rect 16719 19808 16764 19836
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 19610 19836 19616 19848
rect 19571 19808 19616 19836
rect 19610 19796 19616 19808
rect 19668 19796 19674 19848
rect 22281 19839 22339 19845
rect 22281 19805 22293 19839
rect 22327 19836 22339 19839
rect 22370 19836 22376 19848
rect 22327 19808 22376 19836
rect 22327 19805 22339 19808
rect 22281 19799 22339 19805
rect 22370 19796 22376 19808
rect 22428 19836 22434 19848
rect 22738 19836 22744 19848
rect 22428 19808 22744 19836
rect 22428 19796 22434 19808
rect 22738 19796 22744 19808
rect 22796 19796 22802 19848
rect 23290 19796 23296 19848
rect 23348 19836 23354 19848
rect 23385 19839 23443 19845
rect 23385 19836 23397 19839
rect 23348 19808 23397 19836
rect 23348 19796 23354 19808
rect 23385 19805 23397 19808
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 23934 19796 23940 19848
rect 23992 19836 23998 19848
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 23992 19808 24409 19836
rect 23992 19796 23998 19808
rect 24397 19805 24409 19808
rect 24443 19805 24455 19839
rect 24397 19799 24455 19805
rect 24578 19796 24584 19848
rect 24636 19836 24642 19848
rect 24673 19839 24731 19845
rect 24673 19836 24685 19839
rect 24636 19808 24685 19836
rect 24636 19796 24642 19808
rect 24673 19805 24685 19808
rect 24719 19805 24731 19839
rect 26053 19839 26111 19845
rect 26053 19836 26065 19839
rect 24673 19799 24731 19805
rect 24872 19808 26065 19836
rect 14642 19768 14648 19780
rect 12400 19740 12848 19768
rect 14603 19740 14648 19768
rect 12400 19728 12406 19740
rect 14642 19728 14648 19740
rect 14700 19728 14706 19780
rect 20898 19700 20904 19712
rect 20859 19672 20904 19700
rect 20898 19660 20904 19672
rect 20956 19660 20962 19712
rect 23569 19703 23627 19709
rect 23569 19669 23581 19703
rect 23615 19700 23627 19703
rect 24578 19700 24584 19712
rect 23615 19672 24584 19700
rect 23615 19669 23627 19672
rect 23569 19663 23627 19669
rect 24578 19660 24584 19672
rect 24636 19660 24642 19712
rect 24872 19709 24900 19808
rect 26053 19805 26065 19808
rect 26099 19805 26111 19839
rect 26053 19799 26111 19805
rect 26329 19839 26387 19845
rect 26329 19805 26341 19839
rect 26375 19836 26387 19839
rect 28902 19836 28908 19848
rect 26375 19808 28908 19836
rect 26375 19805 26387 19808
rect 26329 19799 26387 19805
rect 28902 19796 28908 19808
rect 28960 19796 28966 19848
rect 37660 19836 37688 19867
rect 36556 19808 37688 19836
rect 35986 19728 35992 19780
rect 36044 19768 36050 19780
rect 36556 19777 36584 19808
rect 36541 19771 36599 19777
rect 36541 19768 36553 19771
rect 36044 19740 36553 19768
rect 36044 19728 36050 19740
rect 36541 19737 36553 19740
rect 36587 19737 36599 19771
rect 36541 19731 36599 19737
rect 24857 19703 24915 19709
rect 24857 19669 24869 19703
rect 24903 19669 24915 19703
rect 36446 19700 36452 19712
rect 36407 19672 36452 19700
rect 24857 19663 24915 19669
rect 36446 19660 36452 19672
rect 36504 19700 36510 19712
rect 37461 19703 37519 19709
rect 37461 19700 37473 19703
rect 36504 19672 37473 19700
rect 36504 19660 36510 19672
rect 37461 19669 37473 19672
rect 37507 19669 37519 19703
rect 37461 19663 37519 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 5353 19499 5411 19505
rect 5353 19496 5365 19499
rect 5224 19468 5365 19496
rect 5224 19456 5230 19468
rect 5353 19465 5365 19468
rect 5399 19465 5411 19499
rect 8386 19496 8392 19508
rect 8347 19468 8392 19496
rect 5353 19459 5411 19465
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 19797 19499 19855 19505
rect 19797 19496 19809 19499
rect 12176 19468 19809 19496
rect 2590 19428 2596 19440
rect 2551 19400 2596 19428
rect 2590 19388 2596 19400
rect 2648 19388 2654 19440
rect 6730 19428 6736 19440
rect 5552 19400 6736 19428
rect 5552 19372 5580 19400
rect 6730 19388 6736 19400
rect 6788 19428 6794 19440
rect 6788 19400 8248 19428
rect 6788 19388 6794 19400
rect 2406 19360 2412 19372
rect 2367 19332 2412 19360
rect 2406 19320 2412 19332
rect 2464 19320 2470 19372
rect 5534 19360 5540 19372
rect 5495 19332 5540 19360
rect 5534 19320 5540 19332
rect 5592 19320 5598 19372
rect 8220 19369 8248 19400
rect 6825 19363 6883 19369
rect 6825 19329 6837 19363
rect 6871 19360 6883 19363
rect 8205 19363 8263 19369
rect 6871 19332 7420 19360
rect 6871 19329 6883 19332
rect 6825 19323 6883 19329
rect 7392 19304 7420 19332
rect 8205 19329 8217 19363
rect 8251 19329 8263 19363
rect 8205 19323 8263 19329
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 12176 19369 12204 19468
rect 19797 19465 19809 19468
rect 19843 19496 19855 19499
rect 22005 19499 22063 19505
rect 19843 19468 21956 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 18785 19431 18843 19437
rect 18785 19397 18797 19431
rect 18831 19428 18843 19431
rect 18874 19428 18880 19440
rect 18831 19400 18880 19428
rect 18831 19397 18843 19400
rect 18785 19391 18843 19397
rect 18874 19388 18880 19400
rect 18932 19388 18938 19440
rect 20717 19431 20775 19437
rect 20717 19428 20729 19431
rect 18984 19400 20729 19428
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 9916 19332 12173 19360
rect 9916 19320 9922 19332
rect 12161 19329 12173 19332
rect 12207 19329 12219 19363
rect 12802 19360 12808 19372
rect 12763 19332 12808 19360
rect 12161 19323 12219 19329
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 14458 19360 14464 19372
rect 14419 19332 14464 19360
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 16758 19320 16764 19372
rect 16816 19360 16822 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16816 19332 16865 19360
rect 16816 19320 16822 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 2866 19292 2872 19304
rect 2827 19264 2872 19292
rect 2866 19252 2872 19264
rect 2924 19252 2930 19304
rect 7374 19252 7380 19304
rect 7432 19292 7438 19304
rect 7469 19295 7527 19301
rect 7469 19292 7481 19295
rect 7432 19264 7481 19292
rect 7432 19252 7438 19264
rect 7469 19261 7481 19264
rect 7515 19261 7527 19295
rect 7469 19255 7527 19261
rect 10870 19184 10876 19236
rect 10928 19224 10934 19236
rect 18984 19233 19012 19400
rect 20717 19397 20729 19400
rect 20763 19397 20775 19431
rect 20717 19391 20775 19397
rect 19886 19360 19892 19372
rect 19847 19332 19892 19360
rect 19886 19320 19892 19332
rect 19944 19320 19950 19372
rect 20732 19360 20760 19391
rect 21821 19363 21879 19369
rect 21821 19360 21833 19363
rect 20732 19332 21833 19360
rect 21821 19329 21833 19332
rect 21867 19329 21879 19363
rect 21928 19360 21956 19468
rect 22005 19465 22017 19499
rect 22051 19496 22063 19499
rect 24581 19499 24639 19505
rect 22051 19468 24348 19496
rect 22051 19465 22063 19468
rect 22005 19459 22063 19465
rect 23290 19428 23296 19440
rect 23251 19400 23296 19428
rect 23290 19388 23296 19400
rect 23348 19388 23354 19440
rect 24320 19372 24348 19468
rect 24581 19465 24593 19499
rect 24627 19496 24639 19499
rect 26418 19496 26424 19508
rect 24627 19468 26424 19496
rect 24627 19465 24639 19468
rect 24581 19459 24639 19465
rect 26418 19456 26424 19468
rect 26476 19456 26482 19508
rect 29914 19496 29920 19508
rect 28000 19468 29920 19496
rect 28000 19440 28028 19468
rect 29914 19456 29920 19468
rect 29972 19456 29978 19508
rect 27062 19388 27068 19440
rect 27120 19428 27126 19440
rect 27249 19431 27307 19437
rect 27249 19428 27261 19431
rect 27120 19400 27261 19428
rect 27120 19388 27126 19400
rect 27249 19397 27261 19400
rect 27295 19428 27307 19431
rect 27982 19428 27988 19440
rect 27295 19400 27988 19428
rect 27295 19397 27307 19400
rect 27249 19391 27307 19397
rect 27982 19388 27988 19400
rect 28040 19388 28046 19440
rect 28902 19428 28908 19440
rect 28863 19400 28908 19428
rect 28902 19388 28908 19400
rect 28960 19388 28966 19440
rect 22462 19360 22468 19372
rect 21928 19332 22468 19360
rect 21821 19323 21879 19329
rect 22462 19320 22468 19332
rect 22520 19320 22526 19372
rect 22646 19320 22652 19372
rect 22704 19360 22710 19372
rect 23382 19360 23388 19372
rect 22704 19332 23388 19360
rect 22704 19320 22710 19332
rect 23382 19320 23388 19332
rect 23440 19360 23446 19372
rect 24118 19360 24124 19372
rect 23440 19332 24124 19360
rect 23440 19320 23446 19332
rect 24118 19320 24124 19332
rect 24176 19320 24182 19372
rect 24302 19360 24308 19372
rect 24215 19332 24308 19360
rect 24302 19320 24308 19332
rect 24360 19320 24366 19372
rect 24397 19363 24455 19369
rect 24397 19329 24409 19363
rect 24443 19360 24455 19363
rect 24578 19360 24584 19372
rect 24443 19332 24584 19360
rect 24443 19329 24455 19332
rect 24397 19323 24455 19329
rect 24578 19320 24584 19332
rect 24636 19320 24642 19372
rect 32306 19360 32312 19372
rect 32267 19332 32312 19360
rect 32306 19320 32312 19332
rect 32364 19320 32370 19372
rect 32490 19360 32496 19372
rect 32451 19332 32496 19360
rect 32490 19320 32496 19332
rect 32548 19320 32554 19372
rect 35434 19320 35440 19372
rect 35492 19360 35498 19372
rect 35601 19363 35659 19369
rect 35601 19360 35613 19363
rect 35492 19332 35613 19360
rect 35492 19320 35498 19332
rect 35601 19329 35613 19332
rect 35647 19329 35659 19363
rect 35601 19323 35659 19329
rect 29089 19295 29147 19301
rect 29089 19261 29101 19295
rect 29135 19292 29147 19295
rect 29822 19292 29828 19304
rect 29135 19264 29828 19292
rect 29135 19261 29147 19264
rect 29089 19255 29147 19261
rect 29822 19252 29828 19264
rect 29880 19252 29886 19304
rect 31662 19292 31668 19304
rect 31128 19264 31668 19292
rect 18969 19227 19027 19233
rect 18969 19224 18981 19227
rect 10928 19196 18981 19224
rect 10928 19184 10934 19196
rect 18969 19193 18981 19196
rect 19015 19193 19027 19227
rect 18969 19187 19027 19193
rect 20622 19184 20628 19236
rect 20680 19224 20686 19236
rect 31128 19224 31156 19264
rect 31662 19252 31668 19264
rect 31720 19252 31726 19304
rect 33045 19295 33103 19301
rect 33045 19261 33057 19295
rect 33091 19292 33103 19295
rect 34514 19292 34520 19304
rect 33091 19264 34520 19292
rect 33091 19261 33103 19264
rect 33045 19255 33103 19261
rect 20680 19196 31156 19224
rect 20680 19184 20686 19196
rect 31202 19184 31208 19236
rect 31260 19224 31266 19236
rect 33060 19224 33088 19255
rect 34514 19252 34520 19264
rect 34572 19292 34578 19304
rect 34793 19295 34851 19301
rect 34793 19292 34805 19295
rect 34572 19264 34805 19292
rect 34572 19252 34578 19264
rect 34793 19261 34805 19264
rect 34839 19292 34851 19295
rect 35345 19295 35403 19301
rect 35345 19292 35357 19295
rect 34839 19264 35357 19292
rect 34839 19261 34851 19264
rect 34793 19255 34851 19261
rect 35345 19261 35357 19264
rect 35391 19261 35403 19295
rect 35345 19255 35403 19261
rect 31260 19196 33088 19224
rect 31260 19184 31266 19196
rect 7006 19156 7012 19168
rect 6967 19128 7012 19156
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 12345 19159 12403 19165
rect 12345 19125 12357 19159
rect 12391 19156 12403 19159
rect 12526 19156 12532 19168
rect 12391 19128 12532 19156
rect 12391 19125 12403 19128
rect 12345 19119 12403 19125
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 12989 19159 13047 19165
rect 12989 19125 13001 19159
rect 13035 19156 13047 19159
rect 13170 19156 13176 19168
rect 13035 19128 13176 19156
rect 13035 19125 13047 19128
rect 12989 19119 13047 19125
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 13446 19156 13452 19168
rect 13407 19128 13452 19156
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 18138 19156 18144 19168
rect 18099 19128 18144 19156
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 20809 19159 20867 19165
rect 20809 19125 20821 19159
rect 20855 19156 20867 19159
rect 22094 19156 22100 19168
rect 20855 19128 22100 19156
rect 20855 19125 20867 19128
rect 20809 19119 20867 19125
rect 22094 19116 22100 19128
rect 22152 19116 22158 19168
rect 22646 19156 22652 19168
rect 22607 19128 22652 19156
rect 22646 19116 22652 19128
rect 22704 19116 22710 19168
rect 24394 19156 24400 19168
rect 24355 19128 24400 19156
rect 24394 19116 24400 19128
rect 24452 19116 24458 19168
rect 32401 19159 32459 19165
rect 32401 19125 32413 19159
rect 32447 19156 32459 19159
rect 32950 19156 32956 19168
rect 32447 19128 32956 19156
rect 32447 19125 32459 19128
rect 32401 19119 32459 19125
rect 32950 19116 32956 19128
rect 33008 19116 33014 19168
rect 34790 19116 34796 19168
rect 34848 19156 34854 19168
rect 35986 19156 35992 19168
rect 34848 19128 35992 19156
rect 34848 19116 34854 19128
rect 35986 19116 35992 19128
rect 36044 19116 36050 19168
rect 36078 19116 36084 19168
rect 36136 19156 36142 19168
rect 36446 19156 36452 19168
rect 36136 19128 36452 19156
rect 36136 19116 36142 19128
rect 36446 19116 36452 19128
rect 36504 19156 36510 19168
rect 36725 19159 36783 19165
rect 36725 19156 36737 19159
rect 36504 19128 36737 19156
rect 36504 19116 36510 19128
rect 36725 19125 36737 19128
rect 36771 19125 36783 19159
rect 36725 19119 36783 19125
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 5997 18955 6055 18961
rect 5997 18921 6009 18955
rect 6043 18952 6055 18955
rect 7282 18952 7288 18964
rect 6043 18924 7288 18952
rect 6043 18921 6055 18924
rect 5997 18915 6055 18921
rect 7282 18912 7288 18924
rect 7340 18952 7346 18964
rect 7653 18955 7711 18961
rect 7653 18952 7665 18955
rect 7340 18924 7665 18952
rect 7340 18912 7346 18924
rect 7653 18921 7665 18924
rect 7699 18921 7711 18955
rect 7653 18915 7711 18921
rect 12342 18912 12348 18964
rect 12400 18952 12406 18964
rect 12621 18955 12679 18961
rect 12621 18952 12633 18955
rect 12400 18924 12633 18952
rect 12400 18912 12406 18924
rect 12621 18921 12633 18924
rect 12667 18921 12679 18955
rect 12621 18915 12679 18921
rect 14277 18955 14335 18961
rect 14277 18921 14289 18955
rect 14323 18952 14335 18955
rect 14642 18952 14648 18964
rect 14323 18924 14648 18952
rect 14323 18921 14335 18924
rect 14277 18915 14335 18921
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 18509 18955 18567 18961
rect 18509 18921 18521 18955
rect 18555 18952 18567 18955
rect 20070 18952 20076 18964
rect 18555 18924 20076 18952
rect 18555 18921 18567 18924
rect 18509 18915 18567 18921
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 23290 18912 23296 18964
rect 23348 18952 23354 18964
rect 23569 18955 23627 18961
rect 23569 18952 23581 18955
rect 23348 18924 23581 18952
rect 23348 18912 23354 18924
rect 23569 18921 23581 18924
rect 23615 18921 23627 18955
rect 24394 18952 24400 18964
rect 24355 18924 24400 18952
rect 23569 18915 23627 18921
rect 24394 18912 24400 18924
rect 24452 18912 24458 18964
rect 29641 18955 29699 18961
rect 29641 18921 29653 18955
rect 29687 18952 29699 18955
rect 29730 18952 29736 18964
rect 29687 18924 29736 18952
rect 29687 18921 29699 18924
rect 29641 18915 29699 18921
rect 29730 18912 29736 18924
rect 29788 18952 29794 18964
rect 30466 18952 30472 18964
rect 29788 18924 30472 18952
rect 29788 18912 29794 18924
rect 30466 18912 30472 18924
rect 30524 18912 30530 18964
rect 34790 18952 34796 18964
rect 30576 18924 34796 18952
rect 8113 18887 8171 18893
rect 8113 18853 8125 18887
rect 8159 18884 8171 18887
rect 8159 18856 21680 18884
rect 8159 18853 8171 18856
rect 8113 18847 8171 18853
rect 5166 18776 5172 18828
rect 5224 18816 5230 18828
rect 5813 18819 5871 18825
rect 5813 18816 5825 18819
rect 5224 18788 5825 18816
rect 5224 18776 5230 18788
rect 5813 18785 5825 18788
rect 5859 18785 5871 18819
rect 5813 18779 5871 18785
rect 6641 18819 6699 18825
rect 6641 18785 6653 18819
rect 6687 18816 6699 18819
rect 7193 18819 7251 18825
rect 7193 18816 7205 18819
rect 6687 18788 7205 18816
rect 6687 18785 6699 18788
rect 6641 18779 6699 18785
rect 7193 18785 7205 18788
rect 7239 18816 7251 18819
rect 7374 18816 7380 18828
rect 7239 18788 7380 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 7374 18776 7380 18788
rect 7432 18816 7438 18828
rect 7742 18816 7748 18828
rect 7432 18788 7748 18816
rect 7432 18776 7438 18788
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 12768 18788 12940 18816
rect 12768 18776 12774 18788
rect 1394 18748 1400 18760
rect 1355 18720 1400 18748
rect 1394 18708 1400 18720
rect 1452 18748 1458 18760
rect 2041 18751 2099 18757
rect 2041 18748 2053 18751
rect 1452 18720 2053 18748
rect 1452 18708 1458 18720
rect 2041 18717 2053 18720
rect 2087 18717 2099 18751
rect 5074 18748 5080 18760
rect 5035 18720 5080 18748
rect 2041 18711 2099 18717
rect 5074 18708 5080 18720
rect 5132 18708 5138 18760
rect 5718 18748 5724 18760
rect 5679 18720 5724 18748
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 7006 18708 7012 18760
rect 7064 18748 7070 18760
rect 7929 18751 7987 18757
rect 7929 18748 7941 18751
rect 7064 18720 7941 18748
rect 7064 18708 7070 18720
rect 7929 18717 7941 18720
rect 7975 18717 7987 18751
rect 7929 18711 7987 18717
rect 9122 18708 9128 18760
rect 9180 18748 9186 18760
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9180 18720 9597 18748
rect 9180 18708 9186 18720
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 10870 18708 10876 18760
rect 10928 18748 10934 18760
rect 12912 18757 12940 18788
rect 18138 18776 18144 18828
rect 18196 18816 18202 18828
rect 19886 18816 19892 18828
rect 18196 18788 19892 18816
rect 18196 18776 18202 18788
rect 11977 18751 12035 18757
rect 11977 18748 11989 18751
rect 10928 18720 11989 18748
rect 10928 18708 10934 18720
rect 11977 18717 11989 18720
rect 12023 18717 12035 18751
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 11977 18711 12035 18717
rect 12452 18720 12817 18748
rect 4614 18640 4620 18692
rect 4672 18680 4678 18692
rect 5997 18683 6055 18689
rect 5997 18680 6009 18683
rect 4672 18652 6009 18680
rect 4672 18640 4678 18652
rect 5828 18624 5856 18652
rect 5997 18649 6009 18652
rect 6043 18649 6055 18683
rect 5997 18643 6055 18649
rect 7466 18640 7472 18692
rect 7524 18680 7530 18692
rect 7653 18683 7711 18689
rect 7653 18680 7665 18683
rect 7524 18652 7665 18680
rect 7524 18640 7530 18652
rect 7653 18649 7665 18652
rect 7699 18680 7711 18683
rect 8202 18680 8208 18692
rect 7699 18652 8208 18680
rect 7699 18649 7711 18652
rect 7653 18643 7711 18649
rect 8202 18640 8208 18652
rect 8260 18680 8266 18692
rect 8941 18683 8999 18689
rect 8941 18680 8953 18683
rect 8260 18652 8953 18680
rect 8260 18640 8266 18652
rect 8941 18649 8953 18652
rect 8987 18649 8999 18683
rect 8941 18643 8999 18649
rect 12452 18624 12480 18720
rect 12805 18717 12817 18720
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 12897 18751 12955 18757
rect 12897 18717 12909 18751
rect 12943 18717 12955 18751
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 12897 18711 12955 18717
rect 13096 18720 14105 18748
rect 12526 18640 12532 18692
rect 12584 18680 12590 18692
rect 12621 18683 12679 18689
rect 12621 18680 12633 18683
rect 12584 18652 12633 18680
rect 12584 18640 12590 18652
rect 12621 18649 12633 18652
rect 12667 18649 12679 18683
rect 12621 18643 12679 18649
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18612 1639 18615
rect 2590 18612 2596 18624
rect 1627 18584 2596 18612
rect 1627 18581 1639 18584
rect 1581 18575 1639 18581
rect 2590 18572 2596 18584
rect 2648 18572 2654 18624
rect 5537 18615 5595 18621
rect 5537 18581 5549 18615
rect 5583 18612 5595 18615
rect 5626 18612 5632 18624
rect 5583 18584 5632 18612
rect 5583 18581 5595 18584
rect 5537 18575 5595 18581
rect 5626 18572 5632 18584
rect 5684 18572 5690 18624
rect 5810 18572 5816 18624
rect 5868 18572 5874 18624
rect 12161 18615 12219 18621
rect 12161 18581 12173 18615
rect 12207 18612 12219 18615
rect 12434 18612 12440 18624
rect 12207 18584 12440 18612
rect 12207 18581 12219 18584
rect 12161 18575 12219 18581
rect 12434 18572 12440 18584
rect 12492 18572 12498 18624
rect 13096 18621 13124 18720
rect 14093 18717 14105 18720
rect 14139 18717 14151 18751
rect 17586 18748 17592 18760
rect 17547 18720 17592 18748
rect 14093 18711 14151 18717
rect 17586 18708 17592 18720
rect 17644 18708 17650 18760
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18748 18383 18751
rect 18414 18748 18420 18760
rect 18371 18720 18420 18748
rect 18371 18717 18383 18720
rect 18325 18711 18383 18717
rect 18414 18708 18420 18720
rect 18472 18748 18478 18760
rect 18874 18748 18880 18760
rect 18472 18720 18880 18748
rect 18472 18708 18478 18720
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19720 18757 19748 18788
rect 19886 18776 19892 18788
rect 19944 18776 19950 18828
rect 19337 18751 19395 18757
rect 19337 18748 19349 18751
rect 19024 18720 19349 18748
rect 19024 18708 19030 18720
rect 19337 18717 19349 18720
rect 19383 18717 19395 18751
rect 19337 18711 19395 18717
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 19981 18751 20039 18757
rect 19981 18717 19993 18751
rect 20027 18717 20039 18751
rect 20714 18748 20720 18760
rect 20675 18720 20720 18748
rect 19981 18711 20039 18717
rect 19996 18680 20024 18711
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 21652 18757 21680 18856
rect 23109 18819 23167 18825
rect 23109 18785 23121 18819
rect 23155 18816 23167 18819
rect 23308 18816 23336 18912
rect 27614 18844 27620 18896
rect 27672 18884 27678 18896
rect 30576 18884 30604 18924
rect 34790 18912 34796 18924
rect 34848 18912 34854 18964
rect 34977 18955 35035 18961
rect 34977 18921 34989 18955
rect 35023 18952 35035 18955
rect 35434 18952 35440 18964
rect 35023 18924 35440 18952
rect 35023 18921 35035 18924
rect 34977 18915 35035 18921
rect 35434 18912 35440 18924
rect 35492 18912 35498 18964
rect 36814 18952 36820 18964
rect 36775 18924 36820 18952
rect 36814 18912 36820 18924
rect 36872 18912 36878 18964
rect 27672 18856 30604 18884
rect 33965 18887 34023 18893
rect 27672 18844 27678 18856
rect 33965 18853 33977 18887
rect 34011 18884 34023 18887
rect 34514 18884 34520 18896
rect 34011 18856 34520 18884
rect 34011 18853 34023 18856
rect 33965 18847 34023 18853
rect 34514 18844 34520 18856
rect 34572 18884 34578 18896
rect 34572 18856 35480 18884
rect 34572 18844 34578 18856
rect 23155 18788 23336 18816
rect 23155 18785 23167 18788
rect 23109 18779 23167 18785
rect 24302 18776 24308 18828
rect 24360 18816 24366 18828
rect 24489 18819 24547 18825
rect 24489 18816 24501 18819
rect 24360 18788 24501 18816
rect 24360 18776 24366 18788
rect 24489 18785 24501 18788
rect 24535 18785 24547 18819
rect 24489 18779 24547 18785
rect 28537 18819 28595 18825
rect 28537 18785 28549 18819
rect 28583 18816 28595 18819
rect 29546 18816 29552 18828
rect 28583 18788 29552 18816
rect 28583 18785 28595 18788
rect 28537 18779 28595 18785
rect 29546 18776 29552 18788
rect 29604 18776 29610 18828
rect 35452 18825 35480 18856
rect 35437 18819 35495 18825
rect 35437 18785 35449 18819
rect 35483 18785 35495 18819
rect 35437 18779 35495 18785
rect 36446 18776 36452 18828
rect 36504 18816 36510 18828
rect 37829 18819 37887 18825
rect 37829 18816 37841 18819
rect 36504 18788 37841 18816
rect 36504 18776 36510 18788
rect 37829 18785 37841 18788
rect 37875 18785 37887 18819
rect 37829 18779 37887 18785
rect 21637 18751 21695 18757
rect 21637 18717 21649 18751
rect 21683 18717 21695 18751
rect 21637 18711 21695 18717
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 22833 18751 22891 18757
rect 22833 18748 22845 18751
rect 22796 18720 22845 18748
rect 22796 18708 22802 18720
rect 22833 18717 22845 18720
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 24118 18708 24124 18760
rect 24176 18748 24182 18760
rect 24397 18751 24455 18757
rect 24397 18748 24409 18751
rect 24176 18720 24409 18748
rect 24176 18708 24182 18720
rect 24397 18717 24409 18720
rect 24443 18717 24455 18751
rect 24397 18711 24455 18717
rect 24578 18708 24584 18760
rect 24636 18748 24642 18760
rect 24673 18751 24731 18757
rect 24673 18748 24685 18751
rect 24636 18720 24685 18748
rect 24636 18708 24642 18720
rect 24673 18717 24685 18720
rect 24719 18717 24731 18751
rect 25777 18751 25835 18757
rect 25777 18748 25789 18751
rect 24673 18711 24731 18717
rect 24872 18720 25789 18748
rect 19352 18652 20024 18680
rect 19352 18624 19380 18652
rect 13081 18615 13139 18621
rect 13081 18581 13093 18615
rect 13127 18581 13139 18615
rect 13081 18575 13139 18581
rect 19334 18572 19340 18624
rect 19392 18572 19398 18624
rect 20622 18612 20628 18624
rect 20583 18584 20628 18612
rect 20622 18572 20628 18584
rect 20680 18572 20686 18624
rect 21818 18612 21824 18624
rect 21779 18584 21824 18612
rect 21818 18572 21824 18584
rect 21876 18572 21882 18624
rect 24872 18621 24900 18720
rect 25777 18717 25789 18720
rect 25823 18717 25835 18751
rect 26418 18748 26424 18760
rect 26379 18720 26424 18748
rect 25777 18711 25835 18717
rect 26418 18708 26424 18720
rect 26476 18708 26482 18760
rect 28994 18708 29000 18760
rect 29052 18748 29058 18760
rect 30745 18751 30803 18757
rect 29052 18720 29097 18748
rect 29052 18708 29058 18720
rect 30745 18717 30757 18751
rect 30791 18748 30803 18751
rect 32582 18748 32588 18760
rect 30791 18720 31248 18748
rect 32543 18720 32588 18748
rect 30791 18717 30803 18720
rect 30745 18711 30803 18717
rect 31220 18692 31248 18720
rect 32582 18708 32588 18720
rect 32640 18708 32646 18760
rect 32677 18751 32735 18757
rect 32677 18717 32689 18751
rect 32723 18717 32735 18751
rect 32677 18711 32735 18717
rect 28813 18683 28871 18689
rect 28813 18649 28825 18683
rect 28859 18649 28871 18683
rect 28813 18643 28871 18649
rect 24857 18615 24915 18621
rect 24857 18581 24869 18615
rect 24903 18581 24915 18615
rect 25958 18612 25964 18624
rect 25919 18584 25964 18612
rect 24857 18575 24915 18581
rect 25958 18572 25964 18584
rect 26016 18572 26022 18624
rect 26605 18615 26663 18621
rect 26605 18581 26617 18615
rect 26651 18612 26663 18615
rect 28828 18612 28856 18643
rect 30834 18640 30840 18692
rect 30892 18680 30898 18692
rect 30990 18683 31048 18689
rect 30990 18680 31002 18683
rect 30892 18652 31002 18680
rect 30892 18640 30898 18652
rect 30990 18649 31002 18652
rect 31036 18649 31048 18683
rect 30990 18643 31048 18649
rect 31202 18640 31208 18692
rect 31260 18640 31266 18692
rect 26651 18584 28856 18612
rect 26651 18581 26663 18584
rect 26605 18575 26663 18581
rect 29822 18572 29828 18624
rect 29880 18612 29886 18624
rect 32125 18615 32183 18621
rect 32125 18612 32137 18615
rect 29880 18584 32137 18612
rect 29880 18572 29886 18584
rect 32125 18581 32137 18584
rect 32171 18612 32183 18615
rect 32692 18612 32720 18711
rect 32766 18708 32772 18760
rect 32824 18748 32830 18760
rect 32861 18751 32919 18757
rect 32861 18748 32873 18751
rect 32824 18720 32873 18748
rect 32824 18708 32830 18720
rect 32861 18717 32873 18720
rect 32907 18717 32919 18751
rect 32861 18711 32919 18717
rect 32950 18708 32956 18760
rect 33008 18748 33014 18760
rect 33778 18748 33784 18760
rect 33008 18720 33053 18748
rect 33739 18720 33784 18748
rect 33008 18708 33014 18720
rect 33778 18708 33784 18720
rect 33836 18708 33842 18760
rect 34606 18708 34612 18760
rect 34664 18748 34670 18760
rect 34793 18751 34851 18757
rect 34793 18748 34805 18751
rect 34664 18720 34805 18748
rect 34664 18708 34670 18720
rect 34793 18717 34805 18720
rect 34839 18717 34851 18751
rect 34793 18711 34851 18717
rect 34977 18751 35035 18757
rect 34977 18717 34989 18751
rect 35023 18748 35035 18751
rect 35526 18748 35532 18760
rect 35023 18720 35532 18748
rect 35023 18717 35035 18720
rect 34977 18711 35035 18717
rect 35526 18708 35532 18720
rect 35584 18708 35590 18760
rect 37402 18751 37460 18757
rect 37402 18748 37414 18751
rect 35820 18720 37414 18748
rect 35820 18692 35848 18720
rect 37402 18717 37414 18720
rect 37448 18717 37460 18751
rect 37402 18711 37460 18717
rect 37918 18708 37924 18760
rect 37976 18748 37982 18760
rect 37976 18720 38021 18748
rect 37976 18708 37982 18720
rect 35342 18640 35348 18692
rect 35400 18680 35406 18692
rect 35682 18683 35740 18689
rect 35682 18680 35694 18683
rect 35400 18652 35694 18680
rect 35400 18640 35406 18652
rect 35682 18649 35694 18652
rect 35728 18649 35740 18683
rect 35682 18643 35740 18649
rect 35802 18640 35808 18692
rect 35860 18640 35866 18692
rect 36814 18640 36820 18692
rect 36872 18680 36878 18692
rect 36872 18652 37504 18680
rect 36872 18640 36878 18652
rect 32171 18584 32720 18612
rect 33137 18615 33195 18621
rect 32171 18581 32183 18584
rect 32125 18575 32183 18581
rect 33137 18581 33149 18615
rect 33183 18612 33195 18615
rect 35434 18612 35440 18624
rect 33183 18584 35440 18612
rect 33183 18581 33195 18584
rect 33137 18575 33195 18581
rect 35434 18572 35440 18584
rect 35492 18572 35498 18624
rect 36906 18572 36912 18624
rect 36964 18612 36970 18624
rect 37476 18621 37504 18652
rect 37277 18615 37335 18621
rect 37277 18612 37289 18615
rect 36964 18584 37289 18612
rect 36964 18572 36970 18584
rect 37277 18581 37289 18584
rect 37323 18581 37335 18615
rect 37277 18575 37335 18581
rect 37461 18615 37519 18621
rect 37461 18581 37473 18615
rect 37507 18581 37519 18615
rect 37461 18575 37519 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 2866 18368 2872 18420
rect 2924 18408 2930 18420
rect 25409 18411 25467 18417
rect 2924 18380 7696 18408
rect 2924 18368 2930 18380
rect 7006 18340 7012 18352
rect 5736 18312 7012 18340
rect 5736 18284 5764 18312
rect 2314 18232 2320 18284
rect 2372 18272 2378 18284
rect 3145 18275 3203 18281
rect 3145 18272 3157 18275
rect 2372 18244 3157 18272
rect 2372 18232 2378 18244
rect 3145 18241 3157 18244
rect 3191 18241 3203 18275
rect 3145 18235 3203 18241
rect 4157 18275 4215 18281
rect 4157 18241 4169 18275
rect 4203 18272 4215 18275
rect 4706 18272 4712 18284
rect 4203 18244 4712 18272
rect 4203 18241 4215 18244
rect 4157 18235 4215 18241
rect 4706 18232 4712 18244
rect 4764 18232 4770 18284
rect 5537 18275 5595 18281
rect 5537 18241 5549 18275
rect 5583 18272 5595 18275
rect 5718 18272 5724 18284
rect 5583 18244 5724 18272
rect 5583 18241 5595 18244
rect 5537 18235 5595 18241
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 5810 18232 5816 18284
rect 5868 18272 5874 18284
rect 6656 18281 6684 18312
rect 7006 18300 7012 18312
rect 7064 18340 7070 18352
rect 7064 18312 7604 18340
rect 7064 18300 7070 18312
rect 6365 18275 6423 18281
rect 6365 18272 6377 18275
rect 5868 18244 6377 18272
rect 5868 18232 5874 18244
rect 6365 18241 6377 18244
rect 6411 18241 6423 18275
rect 6365 18235 6423 18241
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18241 6699 18275
rect 6641 18235 6699 18241
rect 7285 18275 7343 18281
rect 7285 18241 7297 18275
rect 7331 18272 7343 18275
rect 7466 18272 7472 18284
rect 7331 18244 7472 18272
rect 7331 18241 7343 18244
rect 7285 18235 7343 18241
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 7576 18281 7604 18312
rect 7561 18275 7619 18281
rect 7561 18241 7573 18275
rect 7607 18241 7619 18275
rect 7668 18272 7696 18380
rect 10520 18380 14872 18408
rect 9122 18272 9128 18284
rect 7668 18244 8340 18272
rect 9083 18244 9128 18272
rect 7561 18235 7619 18241
rect 5166 18164 5172 18216
rect 5224 18204 5230 18216
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 5224 18176 5641 18204
rect 5224 18164 5230 18176
rect 5629 18173 5641 18176
rect 5675 18173 5687 18207
rect 5629 18167 5687 18173
rect 6549 18207 6607 18213
rect 6549 18173 6561 18207
rect 6595 18204 6607 18207
rect 7374 18204 7380 18216
rect 6595 18176 7380 18204
rect 6595 18173 6607 18176
rect 6549 18167 6607 18173
rect 7374 18164 7380 18176
rect 7432 18204 7438 18216
rect 8205 18207 8263 18213
rect 8205 18204 8217 18207
rect 7432 18176 8217 18204
rect 7432 18164 7438 18176
rect 8205 18173 8217 18176
rect 8251 18173 8263 18207
rect 8205 18167 8263 18173
rect 4893 18139 4951 18145
rect 4893 18105 4905 18139
rect 4939 18136 4951 18139
rect 5534 18136 5540 18148
rect 4939 18108 5540 18136
rect 4939 18105 4951 18108
rect 4893 18099 4951 18105
rect 5534 18096 5540 18108
rect 5592 18096 5598 18148
rect 8312 18136 8340 18244
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 9309 18207 9367 18213
rect 9309 18173 9321 18207
rect 9355 18204 9367 18207
rect 9582 18204 9588 18216
rect 9355 18176 9588 18204
rect 9355 18173 9367 18176
rect 9309 18167 9367 18173
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18204 9735 18207
rect 10520 18204 10548 18380
rect 13170 18340 13176 18352
rect 13131 18312 13176 18340
rect 13170 18300 13176 18312
rect 13228 18300 13234 18352
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18241 12127 18275
rect 12069 18235 12127 18241
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18272 12403 18275
rect 12710 18272 12716 18284
rect 12391 18244 12716 18272
rect 12391 18241 12403 18244
rect 12345 18235 12403 18241
rect 9723 18176 10548 18204
rect 9723 18173 9735 18176
rect 9677 18167 9735 18173
rect 9692 18136 9720 18167
rect 6472 18108 7328 18136
rect 8312 18108 9720 18136
rect 12084 18136 12112 18235
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18204 12311 18207
rect 12434 18204 12440 18216
rect 12299 18176 12440 18204
rect 12299 18173 12311 18176
rect 12253 18167 12311 18173
rect 12434 18164 12440 18176
rect 12492 18204 12498 18216
rect 12618 18204 12624 18216
rect 12492 18176 12624 18204
rect 12492 18164 12498 18176
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18204 13047 18207
rect 13446 18204 13452 18216
rect 13035 18176 13452 18204
rect 13035 18173 13047 18176
rect 12989 18167 13047 18173
rect 13446 18164 13452 18176
rect 13504 18164 13510 18216
rect 14844 18213 14872 18380
rect 25409 18377 25421 18411
rect 25455 18408 25467 18411
rect 29822 18408 29828 18420
rect 25455 18380 29684 18408
rect 29783 18380 29828 18408
rect 25455 18377 25467 18380
rect 25409 18371 25467 18377
rect 17773 18343 17831 18349
rect 17773 18309 17785 18343
rect 17819 18340 17831 18343
rect 18690 18340 18696 18352
rect 17819 18312 18696 18340
rect 17819 18309 17831 18312
rect 17773 18303 17831 18309
rect 18690 18300 18696 18312
rect 18748 18300 18754 18352
rect 21818 18300 21824 18352
rect 21876 18340 21882 18352
rect 24673 18343 24731 18349
rect 24673 18340 24685 18343
rect 21876 18312 24685 18340
rect 21876 18300 21882 18312
rect 24673 18309 24685 18312
rect 24719 18309 24731 18343
rect 24673 18303 24731 18309
rect 17586 18272 17592 18284
rect 17547 18244 17592 18272
rect 17586 18232 17592 18244
rect 17644 18232 17650 18284
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18272 21327 18275
rect 22370 18272 22376 18284
rect 21315 18244 22376 18272
rect 21315 18241 21327 18244
rect 21269 18235 21327 18241
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 24857 18275 24915 18281
rect 24857 18241 24869 18275
rect 24903 18272 24915 18275
rect 25424 18272 25452 18371
rect 25958 18300 25964 18352
rect 26016 18340 26022 18352
rect 27157 18343 27215 18349
rect 27157 18340 27169 18343
rect 26016 18312 27169 18340
rect 26016 18300 26022 18312
rect 27157 18309 27169 18312
rect 27203 18309 27215 18343
rect 27157 18303 27215 18309
rect 27798 18300 27804 18352
rect 27856 18340 27862 18352
rect 28810 18340 28816 18352
rect 27856 18312 28816 18340
rect 27856 18300 27862 18312
rect 28810 18300 28816 18312
rect 28868 18300 28874 18352
rect 29656 18340 29684 18380
rect 29822 18368 29828 18380
rect 29880 18368 29886 18420
rect 29914 18368 29920 18420
rect 29972 18408 29978 18420
rect 30285 18411 30343 18417
rect 29972 18380 30017 18408
rect 29972 18368 29978 18380
rect 30285 18377 30297 18411
rect 30331 18408 30343 18411
rect 32766 18408 32772 18420
rect 30331 18380 30788 18408
rect 32727 18380 32772 18408
rect 30331 18377 30343 18380
rect 30285 18371 30343 18377
rect 30760 18349 30788 18380
rect 32766 18368 32772 18380
rect 32824 18368 32830 18420
rect 35342 18408 35348 18420
rect 35303 18380 35348 18408
rect 35342 18368 35348 18380
rect 35400 18368 35406 18420
rect 35526 18368 35532 18420
rect 35584 18408 35590 18420
rect 35897 18411 35955 18417
rect 35897 18408 35909 18411
rect 35584 18380 35909 18408
rect 35584 18368 35590 18380
rect 35897 18377 35909 18380
rect 35943 18377 35955 18411
rect 36078 18408 36084 18420
rect 36039 18380 36084 18408
rect 35897 18371 35955 18377
rect 36078 18368 36084 18380
rect 36136 18368 36142 18420
rect 37461 18411 37519 18417
rect 37461 18377 37473 18411
rect 37507 18408 37519 18411
rect 37918 18408 37924 18420
rect 37507 18380 37924 18408
rect 37507 18377 37519 18380
rect 37461 18371 37519 18377
rect 37918 18368 37924 18380
rect 37976 18368 37982 18420
rect 30745 18343 30803 18349
rect 29656 18312 30052 18340
rect 24903 18244 25452 18272
rect 30024 18272 30052 18312
rect 30745 18309 30757 18343
rect 30791 18309 30803 18343
rect 30745 18303 30803 18309
rect 30852 18312 31754 18340
rect 30852 18272 30880 18312
rect 30024 18244 30880 18272
rect 30929 18275 30987 18281
rect 24903 18241 24915 18244
rect 24857 18235 24915 18241
rect 30929 18241 30941 18275
rect 30975 18241 30987 18275
rect 31726 18272 31754 18312
rect 32306 18300 32312 18352
rect 32364 18340 32370 18352
rect 32401 18343 32459 18349
rect 32401 18340 32413 18343
rect 32364 18312 32413 18340
rect 32364 18300 32370 18312
rect 32401 18309 32413 18312
rect 32447 18309 32459 18343
rect 32401 18303 32459 18309
rect 32490 18300 32496 18352
rect 32548 18340 32554 18352
rect 32585 18343 32643 18349
rect 32585 18340 32597 18343
rect 32548 18312 32597 18340
rect 32548 18300 32554 18312
rect 32585 18309 32597 18312
rect 32631 18309 32643 18343
rect 36906 18340 36912 18352
rect 32585 18303 32643 18309
rect 35452 18312 36912 18340
rect 31726 18244 34100 18272
rect 30929 18235 30987 18241
rect 14829 18207 14887 18213
rect 14829 18173 14841 18207
rect 14875 18204 14887 18207
rect 17954 18204 17960 18216
rect 14875 18176 17960 18204
rect 14875 18173 14887 18176
rect 14829 18167 14887 18173
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 18230 18204 18236 18216
rect 18191 18176 18236 18204
rect 18230 18164 18236 18176
rect 18288 18164 18294 18216
rect 24394 18204 24400 18216
rect 24355 18176 24400 18204
rect 24394 18164 24400 18176
rect 24452 18164 24458 18216
rect 26973 18207 27031 18213
rect 26973 18173 26985 18207
rect 27019 18204 27031 18207
rect 27614 18204 27620 18216
rect 27019 18176 27620 18204
rect 27019 18173 27031 18176
rect 26973 18167 27031 18173
rect 27614 18164 27620 18176
rect 27672 18164 27678 18216
rect 29730 18204 29736 18216
rect 29691 18176 29736 18204
rect 29730 18164 29736 18176
rect 29788 18164 29794 18216
rect 30944 18204 30972 18235
rect 31662 18204 31668 18216
rect 30944 18176 31668 18204
rect 31662 18164 31668 18176
rect 31720 18204 31726 18216
rect 33962 18204 33968 18216
rect 31720 18176 33968 18204
rect 31720 18164 31726 18176
rect 33962 18164 33968 18176
rect 34020 18164 34026 18216
rect 34072 18204 34100 18244
rect 34606 18232 34612 18284
rect 34664 18272 34670 18284
rect 35452 18281 35480 18312
rect 36906 18300 36912 18312
rect 36964 18300 36970 18352
rect 35253 18275 35311 18281
rect 35253 18272 35265 18275
rect 34664 18244 35265 18272
rect 34664 18232 34670 18244
rect 35253 18241 35265 18244
rect 35299 18241 35311 18275
rect 35253 18235 35311 18241
rect 35437 18275 35495 18281
rect 35437 18241 35449 18275
rect 35483 18241 35495 18275
rect 35437 18235 35495 18241
rect 35802 18232 35808 18284
rect 35860 18272 35866 18284
rect 36022 18275 36080 18281
rect 36022 18272 36034 18275
rect 35860 18244 36034 18272
rect 35860 18232 35866 18244
rect 36022 18241 36034 18244
rect 36068 18241 36080 18275
rect 36446 18272 36452 18284
rect 36407 18244 36452 18272
rect 36022 18235 36080 18241
rect 36446 18232 36452 18244
rect 36504 18232 36510 18284
rect 36541 18275 36599 18281
rect 36541 18241 36553 18275
rect 36587 18272 36599 18275
rect 37461 18275 37519 18281
rect 37461 18272 37473 18275
rect 36587 18244 37473 18272
rect 36587 18241 36599 18244
rect 36541 18235 36599 18241
rect 37461 18241 37473 18244
rect 37507 18272 37519 18275
rect 37826 18272 37832 18284
rect 37507 18244 37832 18272
rect 37507 18241 37519 18244
rect 37461 18235 37519 18241
rect 36262 18204 36268 18216
rect 34072 18176 36268 18204
rect 36262 18164 36268 18176
rect 36320 18164 36326 18216
rect 12084 18108 12480 18136
rect 3234 18068 3240 18080
rect 3195 18040 3240 18068
rect 3234 18028 3240 18040
rect 3292 18028 3298 18080
rect 5350 18068 5356 18080
rect 5311 18040 5356 18068
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 6472 18077 6500 18108
rect 7300 18080 7328 18108
rect 12452 18080 12480 18108
rect 32582 18096 32588 18148
rect 32640 18136 32646 18148
rect 36556 18136 36584 18235
rect 37826 18232 37832 18244
rect 37884 18232 37890 18284
rect 32640 18108 36584 18136
rect 32640 18096 32646 18108
rect 5813 18071 5871 18077
rect 5813 18037 5825 18071
rect 5859 18068 5871 18071
rect 6457 18071 6515 18077
rect 6457 18068 6469 18071
rect 5859 18040 6469 18068
rect 5859 18037 5871 18040
rect 5813 18031 5871 18037
rect 6457 18037 6469 18040
rect 6503 18037 6515 18071
rect 6457 18031 6515 18037
rect 6546 18028 6552 18080
rect 6604 18068 6610 18080
rect 6825 18071 6883 18077
rect 6825 18068 6837 18071
rect 6604 18040 6837 18068
rect 6604 18028 6610 18040
rect 6825 18037 6837 18040
rect 6871 18037 6883 18071
rect 7282 18068 7288 18080
rect 7243 18040 7288 18068
rect 6825 18031 6883 18037
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 7742 18068 7748 18080
rect 7703 18040 7748 18068
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 12342 18068 12348 18080
rect 12303 18040 12348 18068
rect 12342 18028 12348 18040
rect 12400 18028 12406 18080
rect 12434 18028 12440 18080
rect 12492 18028 12498 18080
rect 12529 18071 12587 18077
rect 12529 18037 12541 18071
rect 12575 18068 12587 18071
rect 13170 18068 13176 18080
rect 12575 18040 13176 18068
rect 12575 18037 12587 18040
rect 12529 18031 12587 18037
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 20070 18068 20076 18080
rect 20031 18040 20076 18068
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 22278 18068 22284 18080
rect 22239 18040 22284 18068
rect 22278 18028 22284 18040
rect 22336 18028 22342 18080
rect 30558 18028 30564 18080
rect 30616 18068 30622 18080
rect 31113 18071 31171 18077
rect 31113 18068 31125 18071
rect 30616 18040 31125 18068
rect 30616 18028 30622 18040
rect 31113 18037 31125 18040
rect 31159 18037 31171 18071
rect 31113 18031 31171 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1578 17824 1584 17876
rect 1636 17864 1642 17876
rect 2130 17864 2136 17876
rect 1636 17836 2136 17864
rect 1636 17824 1642 17836
rect 2130 17824 2136 17836
rect 2188 17864 2194 17876
rect 2501 17867 2559 17873
rect 2501 17864 2513 17867
rect 2188 17836 2513 17864
rect 2188 17824 2194 17836
rect 2501 17833 2513 17836
rect 2547 17833 2559 17867
rect 2501 17827 2559 17833
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 3927 17867 3985 17873
rect 3927 17864 3939 17867
rect 3108 17836 3939 17864
rect 3108 17824 3114 17836
rect 3927 17833 3939 17836
rect 3973 17833 3985 17867
rect 3927 17827 3985 17833
rect 5074 17824 5080 17876
rect 5132 17824 5138 17876
rect 7466 17824 7472 17876
rect 7524 17864 7530 17876
rect 7745 17867 7803 17873
rect 7745 17864 7757 17867
rect 7524 17836 7757 17864
rect 7524 17824 7530 17836
rect 7745 17833 7757 17836
rect 7791 17833 7803 17867
rect 8386 17864 8392 17876
rect 8347 17836 8392 17864
rect 7745 17827 7803 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 9398 17864 9404 17876
rect 9359 17836 9404 17864
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 9582 17824 9588 17876
rect 9640 17864 9646 17876
rect 10229 17867 10287 17873
rect 10229 17864 10241 17867
rect 9640 17836 10241 17864
rect 9640 17824 9646 17836
rect 10229 17833 10241 17836
rect 10275 17833 10287 17867
rect 12342 17864 12348 17876
rect 12303 17836 12348 17864
rect 10229 17827 10287 17833
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 12452 17836 12848 17864
rect 3602 17756 3608 17808
rect 3660 17796 3666 17808
rect 4062 17796 4068 17808
rect 3660 17768 4068 17796
rect 3660 17756 3666 17768
rect 4062 17756 4068 17768
rect 4120 17756 4126 17808
rect 2590 17728 2596 17740
rect 2551 17700 2596 17728
rect 2590 17688 2596 17700
rect 2648 17688 2654 17740
rect 3234 17688 3240 17740
rect 3292 17728 3298 17740
rect 5092 17737 5120 17824
rect 5166 17756 5172 17808
rect 5224 17796 5230 17808
rect 9674 17796 9680 17808
rect 5224 17768 9680 17796
rect 5224 17756 5230 17768
rect 9674 17756 9680 17768
rect 9732 17756 9738 17808
rect 9769 17799 9827 17805
rect 9769 17765 9781 17799
rect 9815 17765 9827 17799
rect 12452 17796 12480 17836
rect 9769 17759 9827 17765
rect 10796 17768 12480 17796
rect 4157 17731 4215 17737
rect 4157 17728 4169 17731
rect 3292 17700 4169 17728
rect 3292 17688 3298 17700
rect 4157 17697 4169 17700
rect 4203 17697 4215 17731
rect 4157 17691 4215 17697
rect 5077 17731 5135 17737
rect 5077 17697 5089 17731
rect 5123 17697 5135 17731
rect 5534 17728 5540 17740
rect 5495 17700 5540 17728
rect 5077 17691 5135 17697
rect 1394 17660 1400 17672
rect 1355 17632 1400 17660
rect 1394 17620 1400 17632
rect 1452 17620 1458 17672
rect 2498 17660 2504 17672
rect 2459 17632 2504 17660
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 3789 17595 3847 17601
rect 3789 17561 3801 17595
rect 3835 17561 3847 17595
rect 4172 17592 4200 17691
rect 5534 17688 5540 17700
rect 5592 17688 5598 17740
rect 8386 17688 8392 17740
rect 8444 17728 8450 17740
rect 9401 17731 9459 17737
rect 9401 17728 9413 17731
rect 8444 17700 9413 17728
rect 8444 17688 8450 17700
rect 9401 17697 9413 17700
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 9582 17620 9588 17672
rect 9640 17660 9646 17672
rect 9784 17660 9812 17759
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 9640 17632 9685 17660
rect 9784 17632 10425 17660
rect 9640 17620 9646 17632
rect 10413 17629 10425 17632
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 5074 17592 5080 17604
rect 4172 17564 5080 17592
rect 3789 17555 3847 17561
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17524 1639 17527
rect 2590 17524 2596 17536
rect 1627 17496 2596 17524
rect 1627 17493 1639 17496
rect 1581 17487 1639 17493
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 2869 17527 2927 17533
rect 2869 17493 2881 17527
rect 2915 17524 2927 17527
rect 3804 17524 3832 17555
rect 5074 17552 5080 17564
rect 5132 17552 5138 17604
rect 5261 17595 5319 17601
rect 5261 17561 5273 17595
rect 5307 17592 5319 17595
rect 5442 17592 5448 17604
rect 5307 17564 5448 17592
rect 5307 17561 5319 17564
rect 5261 17555 5319 17561
rect 5442 17552 5448 17564
rect 5500 17552 5506 17604
rect 9306 17592 9312 17604
rect 9267 17564 9312 17592
rect 9306 17552 9312 17564
rect 9364 17552 9370 17604
rect 10796 17592 10824 17768
rect 12526 17756 12532 17808
rect 12584 17796 12590 17808
rect 12820 17796 12848 17836
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 16117 17867 16175 17873
rect 16117 17864 16129 17867
rect 15252 17836 16129 17864
rect 15252 17824 15258 17836
rect 16117 17833 16129 17836
rect 16163 17833 16175 17867
rect 16117 17827 16175 17833
rect 16298 17824 16304 17876
rect 16356 17864 16362 17876
rect 16850 17864 16856 17876
rect 16356 17836 16856 17864
rect 16356 17824 16362 17836
rect 16850 17824 16856 17836
rect 16908 17864 16914 17876
rect 18233 17867 18291 17873
rect 18233 17864 18245 17867
rect 16908 17836 18245 17864
rect 16908 17824 16914 17836
rect 18233 17833 18245 17836
rect 18279 17864 18291 17867
rect 18598 17864 18604 17876
rect 18279 17836 18604 17864
rect 18279 17833 18291 17836
rect 18233 17827 18291 17833
rect 18598 17824 18604 17836
rect 18656 17864 18662 17876
rect 20254 17864 20260 17876
rect 18656 17836 20260 17864
rect 18656 17824 18662 17836
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 29641 17867 29699 17873
rect 29641 17833 29653 17867
rect 29687 17864 29699 17867
rect 29914 17864 29920 17876
rect 29687 17836 29920 17864
rect 29687 17833 29699 17836
rect 29641 17827 29699 17833
rect 29914 17824 29920 17836
rect 29972 17824 29978 17876
rect 30745 17867 30803 17873
rect 30745 17833 30757 17867
rect 30791 17864 30803 17867
rect 30834 17864 30840 17876
rect 30791 17836 30840 17864
rect 30791 17833 30803 17836
rect 30745 17827 30803 17833
rect 30834 17824 30840 17836
rect 30892 17824 30898 17876
rect 32582 17864 32588 17876
rect 32543 17836 32588 17864
rect 32582 17824 32588 17836
rect 32640 17824 32646 17876
rect 38010 17864 38016 17876
rect 37971 17836 38016 17864
rect 38010 17824 38016 17836
rect 38068 17824 38074 17876
rect 18138 17796 18144 17808
rect 12584 17768 12756 17796
rect 12820 17768 18144 17796
rect 12584 17756 12590 17768
rect 12728 17740 12756 17768
rect 18138 17756 18144 17768
rect 18196 17756 18202 17808
rect 18782 17756 18788 17808
rect 18840 17796 18846 17808
rect 27154 17796 27160 17808
rect 18840 17768 27160 17796
rect 18840 17756 18846 17768
rect 27154 17756 27160 17768
rect 27212 17756 27218 17808
rect 12437 17731 12495 17737
rect 12437 17697 12449 17731
rect 12483 17728 12495 17731
rect 12618 17728 12624 17740
rect 12483 17700 12624 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 12710 17688 12716 17740
rect 12768 17688 12774 17740
rect 18506 17728 18512 17740
rect 13004 17700 18512 17728
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17660 12311 17663
rect 12342 17660 12348 17672
rect 12299 17632 12348 17660
rect 12299 17629 12311 17632
rect 12253 17623 12311 17629
rect 12342 17620 12348 17632
rect 12400 17620 12406 17672
rect 12526 17660 12532 17672
rect 12487 17632 12532 17660
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 13004 17660 13032 17700
rect 18506 17688 18512 17700
rect 18564 17688 18570 17740
rect 20070 17728 20076 17740
rect 20031 17700 20076 17728
rect 20070 17688 20076 17700
rect 20128 17688 20134 17740
rect 21913 17731 21971 17737
rect 21913 17697 21925 17731
rect 21959 17728 21971 17731
rect 23842 17728 23848 17740
rect 21959 17700 23848 17728
rect 21959 17697 21971 17700
rect 21913 17691 21971 17697
rect 23842 17688 23848 17700
rect 23900 17688 23906 17740
rect 13170 17660 13176 17672
rect 12636 17632 13032 17660
rect 13131 17632 13176 17660
rect 12636 17592 12664 17632
rect 13170 17620 13176 17632
rect 13228 17620 13234 17672
rect 13354 17620 13360 17672
rect 13412 17660 13418 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13412 17632 14105 17660
rect 13412 17620 13418 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 16298 17660 16304 17672
rect 16259 17632 16304 17660
rect 14093 17623 14151 17629
rect 16298 17620 16304 17632
rect 16356 17620 16362 17672
rect 30558 17660 30564 17672
rect 16408 17632 19380 17660
rect 30519 17632 30564 17660
rect 9784 17564 10824 17592
rect 12406 17564 12664 17592
rect 9784 17563 9812 17564
rect 2915 17496 3832 17524
rect 4433 17527 4491 17533
rect 2915 17493 2927 17496
rect 2869 17487 2927 17493
rect 4433 17493 4445 17527
rect 4479 17524 4491 17527
rect 4982 17524 4988 17536
rect 4479 17496 4988 17524
rect 4479 17493 4491 17496
rect 4433 17487 4491 17493
rect 4982 17484 4988 17496
rect 5040 17524 5046 17536
rect 9692 17535 9812 17563
rect 9692 17524 9720 17535
rect 5040 17496 9720 17524
rect 5040 17484 5046 17496
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 12406 17524 12434 17564
rect 12894 17552 12900 17604
rect 12952 17592 12958 17604
rect 16408 17592 16436 17632
rect 12952 17564 16436 17592
rect 18141 17595 18199 17601
rect 12952 17552 12958 17564
rect 18141 17561 18153 17595
rect 18187 17592 18199 17595
rect 19242 17592 19248 17604
rect 18187 17564 19248 17592
rect 18187 17561 18199 17564
rect 18141 17555 18199 17561
rect 9916 17496 12434 17524
rect 12713 17527 12771 17533
rect 9916 17484 9922 17496
rect 12713 17493 12725 17527
rect 12759 17524 12771 17527
rect 12802 17524 12808 17536
rect 12759 17496 12808 17524
rect 12759 17493 12771 17496
rect 12713 17487 12771 17493
rect 12802 17484 12808 17496
rect 12860 17484 12866 17536
rect 13357 17527 13415 17533
rect 13357 17493 13369 17527
rect 13403 17524 13415 17527
rect 13538 17524 13544 17536
rect 13403 17496 13544 17524
rect 13403 17493 13415 17496
rect 13357 17487 13415 17493
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 17589 17527 17647 17533
rect 17589 17493 17601 17527
rect 17635 17524 17647 17527
rect 17770 17524 17776 17536
rect 17635 17496 17776 17524
rect 17635 17493 17647 17496
rect 17589 17487 17647 17493
rect 17770 17484 17776 17496
rect 17828 17524 17834 17536
rect 18156 17524 18184 17555
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 17828 17496 18184 17524
rect 19352 17524 19380 17632
rect 30558 17620 30564 17632
rect 30616 17620 30622 17672
rect 31202 17660 31208 17672
rect 31163 17632 31208 17660
rect 31202 17620 31208 17632
rect 31260 17660 31266 17672
rect 33137 17663 33195 17669
rect 33137 17660 33149 17663
rect 31260 17632 33149 17660
rect 31260 17620 31266 17632
rect 33137 17629 33149 17632
rect 33183 17660 33195 17663
rect 35253 17663 35311 17669
rect 35253 17660 35265 17663
rect 33183 17632 35265 17660
rect 33183 17629 33195 17632
rect 33137 17623 33195 17629
rect 35253 17629 35265 17632
rect 35299 17660 35311 17663
rect 35618 17660 35624 17672
rect 35299 17632 35624 17660
rect 35299 17629 35311 17632
rect 35253 17623 35311 17629
rect 35618 17620 35624 17632
rect 35676 17620 35682 17672
rect 37369 17663 37427 17669
rect 37369 17629 37381 17663
rect 37415 17660 37427 17663
rect 37734 17660 37740 17672
rect 37415 17632 37740 17660
rect 37415 17629 37427 17632
rect 37369 17623 37427 17629
rect 37734 17620 37740 17632
rect 37792 17660 37798 17672
rect 37829 17663 37887 17669
rect 37829 17660 37841 17663
rect 37792 17632 37841 17660
rect 37792 17620 37798 17632
rect 37829 17629 37841 17632
rect 37875 17629 37887 17663
rect 37829 17623 37887 17629
rect 20254 17592 20260 17604
rect 20215 17564 20260 17592
rect 20254 17552 20260 17564
rect 20312 17552 20318 17604
rect 31478 17601 31484 17604
rect 31472 17555 31484 17601
rect 31536 17592 31542 17604
rect 31536 17564 31572 17592
rect 31478 17552 31484 17555
rect 31536 17552 31542 17564
rect 22738 17524 22744 17536
rect 19352 17496 22744 17524
rect 17828 17484 17834 17496
rect 22738 17484 22744 17496
rect 22796 17484 22802 17536
rect 30558 17484 30564 17536
rect 30616 17524 30622 17536
rect 31386 17524 31392 17536
rect 30616 17496 31392 17524
rect 30616 17484 30622 17496
rect 31386 17484 31392 17496
rect 31444 17484 31450 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 3421 17323 3479 17329
rect 3421 17289 3433 17323
rect 3467 17320 3479 17323
rect 5442 17320 5448 17332
rect 3467 17292 5304 17320
rect 5403 17292 5448 17320
rect 3467 17289 3479 17292
rect 3421 17283 3479 17289
rect 1394 17252 1400 17264
rect 1355 17224 1400 17252
rect 1394 17212 1400 17224
rect 1452 17212 1458 17264
rect 2958 17252 2964 17264
rect 2871 17224 2964 17252
rect 2958 17212 2964 17224
rect 3016 17252 3022 17264
rect 3973 17255 4031 17261
rect 3973 17252 3985 17255
rect 3016 17224 3985 17252
rect 3016 17212 3022 17224
rect 3973 17221 3985 17224
rect 4019 17221 4031 17255
rect 5276 17252 5304 17292
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 9306 17280 9312 17332
rect 9364 17320 9370 17332
rect 10134 17320 10140 17332
rect 9364 17292 10140 17320
rect 9364 17280 9370 17292
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 18782 17320 18788 17332
rect 12406 17292 18184 17320
rect 18743 17292 18788 17320
rect 12406 17252 12434 17292
rect 18156 17264 18184 17292
rect 18782 17280 18788 17292
rect 18840 17280 18846 17332
rect 20714 17280 20720 17332
rect 20772 17320 20778 17332
rect 20809 17323 20867 17329
rect 20809 17320 20821 17323
rect 20772 17292 20821 17320
rect 20772 17280 20778 17292
rect 20809 17289 20821 17292
rect 20855 17320 20867 17323
rect 29546 17320 29552 17332
rect 20855 17292 26234 17320
rect 29459 17292 29552 17320
rect 20855 17289 20867 17292
rect 20809 17283 20867 17289
rect 13538 17252 13544 17264
rect 5276 17224 12434 17252
rect 13499 17224 13544 17252
rect 3973 17215 4031 17221
rect 13538 17212 13544 17224
rect 13596 17212 13602 17264
rect 18138 17252 18144 17264
rect 18051 17224 18144 17252
rect 18138 17212 18144 17224
rect 18196 17212 18202 17264
rect 22465 17255 22523 17261
rect 22465 17221 22477 17255
rect 22511 17252 22523 17255
rect 23106 17252 23112 17264
rect 22511 17224 23112 17252
rect 22511 17221 22523 17224
rect 22465 17215 22523 17221
rect 23106 17212 23112 17224
rect 23164 17252 23170 17264
rect 23382 17252 23388 17264
rect 23164 17224 23388 17252
rect 23164 17212 23170 17224
rect 23382 17212 23388 17224
rect 23440 17212 23446 17264
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2498 17184 2504 17196
rect 2179 17156 2504 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 2682 17144 2688 17196
rect 2740 17184 2746 17196
rect 3142 17184 3148 17196
rect 2740 17156 3148 17184
rect 2740 17144 2746 17156
rect 3142 17144 3148 17156
rect 3200 17184 3206 17196
rect 3237 17187 3295 17193
rect 3237 17184 3249 17187
rect 3200 17156 3249 17184
rect 3200 17144 3206 17156
rect 3237 17153 3249 17156
rect 3283 17153 3295 17187
rect 3237 17147 3295 17153
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17153 4307 17187
rect 5626 17184 5632 17196
rect 5587 17156 5632 17184
rect 4249 17147 4307 17153
rect 2225 17119 2283 17125
rect 2225 17085 2237 17119
rect 2271 17116 2283 17119
rect 2314 17116 2320 17128
rect 2271 17088 2320 17116
rect 2271 17085 2283 17088
rect 2225 17079 2283 17085
rect 2314 17076 2320 17088
rect 2372 17076 2378 17128
rect 3050 17116 3056 17128
rect 3011 17088 3056 17116
rect 3050 17076 3056 17088
rect 3108 17116 3114 17128
rect 3970 17116 3976 17128
rect 3108 17088 3976 17116
rect 3108 17076 3114 17088
rect 3970 17076 3976 17088
rect 4028 17116 4034 17128
rect 4065 17119 4123 17125
rect 4065 17116 4077 17119
rect 4028 17088 4077 17116
rect 4028 17076 4034 17088
rect 4065 17085 4077 17088
rect 4111 17085 4123 17119
rect 4065 17079 4123 17085
rect 2332 17048 2360 17076
rect 4264 17048 4292 17147
rect 5626 17144 5632 17156
rect 5684 17144 5690 17196
rect 9674 17184 9680 17196
rect 9646 17144 9680 17184
rect 9732 17144 9738 17196
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12713 17187 12771 17193
rect 12492 17156 12537 17184
rect 12492 17144 12498 17156
rect 12713 17153 12725 17187
rect 12759 17184 12771 17187
rect 12894 17184 12900 17196
rect 12759 17156 12900 17184
rect 12759 17153 12771 17156
rect 12713 17147 12771 17153
rect 12894 17144 12900 17156
rect 12952 17144 12958 17196
rect 13354 17184 13360 17196
rect 13315 17156 13360 17184
rect 13354 17144 13360 17156
rect 13412 17144 13418 17196
rect 22738 17184 22744 17196
rect 22699 17156 22744 17184
rect 22738 17144 22744 17156
rect 22796 17184 22802 17196
rect 23198 17184 23204 17196
rect 22796 17156 23204 17184
rect 22796 17144 22802 17156
rect 23198 17144 23204 17156
rect 23256 17184 23262 17196
rect 23661 17187 23719 17193
rect 23661 17184 23673 17187
rect 23256 17156 23673 17184
rect 23256 17144 23262 17156
rect 23661 17153 23673 17156
rect 23707 17153 23719 17187
rect 23661 17147 23719 17153
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 9646 17116 9674 17144
rect 12618 17116 12624 17128
rect 5592 17088 9674 17116
rect 12579 17088 12624 17116
rect 5592 17076 5598 17088
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 15102 17116 15108 17128
rect 15015 17088 15108 17116
rect 15102 17076 15108 17088
rect 15160 17116 15166 17128
rect 18230 17116 18236 17128
rect 15160 17088 18236 17116
rect 15160 17076 15166 17088
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 18506 17116 18512 17128
rect 18467 17088 18512 17116
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 22649 17119 22707 17125
rect 22649 17085 22661 17119
rect 22695 17116 22707 17119
rect 23474 17116 23480 17128
rect 22695 17088 23480 17116
rect 22695 17085 22707 17088
rect 22649 17079 22707 17085
rect 23474 17076 23480 17088
rect 23532 17116 23538 17128
rect 24302 17116 24308 17128
rect 23532 17088 24308 17116
rect 23532 17076 23538 17088
rect 24302 17076 24308 17088
rect 24360 17076 24366 17128
rect 26206 17116 26234 17292
rect 29546 17280 29552 17292
rect 29604 17320 29610 17332
rect 30377 17323 30435 17329
rect 30377 17320 30389 17323
rect 29604 17292 30389 17320
rect 29604 17280 29610 17292
rect 30377 17289 30389 17292
rect 30423 17320 30435 17323
rect 30558 17320 30564 17332
rect 30423 17292 30564 17320
rect 30423 17289 30435 17292
rect 30377 17283 30435 17289
rect 30558 17280 30564 17292
rect 30616 17280 30622 17332
rect 31389 17323 31447 17329
rect 31389 17289 31401 17323
rect 31435 17320 31447 17323
rect 31478 17320 31484 17332
rect 31435 17292 31484 17320
rect 31435 17289 31447 17292
rect 31389 17283 31447 17289
rect 31478 17280 31484 17292
rect 31536 17280 31542 17332
rect 35618 17320 35624 17332
rect 35579 17292 35624 17320
rect 35618 17280 35624 17292
rect 35676 17280 35682 17332
rect 28994 17212 29000 17264
rect 29052 17252 29058 17264
rect 30469 17255 30527 17261
rect 30469 17252 30481 17255
rect 29052 17224 30481 17252
rect 29052 17212 29058 17224
rect 30469 17221 30481 17224
rect 30515 17252 30527 17255
rect 32582 17252 32588 17264
rect 30515 17224 32588 17252
rect 30515 17221 30527 17224
rect 30469 17215 30527 17221
rect 32582 17212 32588 17224
rect 32640 17212 32646 17264
rect 27246 17184 27252 17196
rect 27207 17156 27252 17184
rect 27246 17144 27252 17156
rect 27304 17144 27310 17196
rect 30190 17144 30196 17196
rect 30248 17184 30254 17196
rect 30248 17156 30604 17184
rect 30248 17144 30254 17156
rect 30576 17125 30604 17156
rect 30650 17144 30656 17196
rect 30708 17184 30714 17196
rect 31205 17187 31263 17193
rect 31205 17184 31217 17187
rect 30708 17156 31217 17184
rect 30708 17144 30714 17156
rect 31205 17153 31217 17156
rect 31251 17153 31263 17187
rect 31205 17147 31263 17153
rect 30561 17119 30619 17125
rect 26206 17088 30512 17116
rect 22278 17048 22284 17060
rect 2332 17020 4292 17048
rect 12728 17020 22284 17048
rect 12728 16992 12756 17020
rect 22278 17008 22284 17020
rect 22336 17048 22342 17060
rect 22336 17020 23428 17048
rect 22336 17008 22342 17020
rect 2130 16980 2136 16992
rect 2091 16952 2136 16980
rect 2130 16940 2136 16952
rect 2188 16980 2194 16992
rect 2406 16980 2412 16992
rect 2188 16952 2412 16980
rect 2188 16940 2194 16952
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 2501 16983 2559 16989
rect 2501 16949 2513 16983
rect 2547 16980 2559 16983
rect 2866 16980 2872 16992
rect 2547 16952 2872 16980
rect 2547 16949 2559 16952
rect 2501 16943 2559 16949
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 3237 16983 3295 16989
rect 3237 16949 3249 16983
rect 3283 16980 3295 16983
rect 4062 16980 4068 16992
rect 3283 16952 4068 16980
rect 3283 16949 3295 16952
rect 3237 16943 3295 16949
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 4433 16983 4491 16989
rect 4433 16949 4445 16983
rect 4479 16980 4491 16983
rect 8386 16980 8392 16992
rect 4479 16952 8392 16980
rect 4479 16949 4491 16952
rect 4433 16943 4491 16949
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 9122 16980 9128 16992
rect 9083 16952 9128 16980
rect 9122 16940 9128 16952
rect 9180 16940 9186 16992
rect 12710 16980 12716 16992
rect 12623 16952 12716 16980
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 18322 16989 18328 16992
rect 18306 16983 18328 16989
rect 18306 16949 18318 16983
rect 18306 16943 18328 16949
rect 18322 16940 18328 16943
rect 18380 16940 18386 16992
rect 18414 16940 18420 16992
rect 18472 16980 18478 16992
rect 22480 16989 22508 17020
rect 23400 16992 23428 17020
rect 27154 17008 27160 17060
rect 27212 17048 27218 17060
rect 29730 17048 29736 17060
rect 27212 17020 29736 17048
rect 27212 17008 27218 17020
rect 29730 17008 29736 17020
rect 29788 17008 29794 17060
rect 22465 16983 22523 16989
rect 18472 16952 18517 16980
rect 18472 16940 18478 16952
rect 22465 16949 22477 16983
rect 22511 16949 22523 16983
rect 22922 16980 22928 16992
rect 22883 16952 22928 16980
rect 22465 16943 22523 16949
rect 22922 16940 22928 16952
rect 22980 16940 22986 16992
rect 23382 16980 23388 16992
rect 23295 16952 23388 16980
rect 23382 16940 23388 16952
rect 23440 16940 23446 16992
rect 23842 16980 23848 16992
rect 23803 16952 23848 16980
rect 23842 16940 23848 16952
rect 23900 16940 23906 16992
rect 26878 16940 26884 16992
rect 26936 16980 26942 16992
rect 27065 16983 27123 16989
rect 27065 16980 27077 16983
rect 26936 16952 27077 16980
rect 26936 16940 26942 16952
rect 27065 16949 27077 16952
rect 27111 16949 27123 16983
rect 27065 16943 27123 16949
rect 30009 16983 30067 16989
rect 30009 16949 30021 16983
rect 30055 16980 30067 16983
rect 30282 16980 30288 16992
rect 30055 16952 30288 16980
rect 30055 16949 30067 16952
rect 30009 16943 30067 16949
rect 30282 16940 30288 16952
rect 30340 16940 30346 16992
rect 30484 16980 30512 17088
rect 30561 17085 30573 17119
rect 30607 17116 30619 17119
rect 31018 17116 31024 17128
rect 30607 17088 31024 17116
rect 30607 17085 30619 17088
rect 30561 17079 30619 17085
rect 31018 17076 31024 17088
rect 31076 17076 31082 17128
rect 32674 16980 32680 16992
rect 30484 16952 32680 16980
rect 32674 16940 32680 16952
rect 32732 16940 32738 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 2958 16776 2964 16788
rect 2919 16748 2964 16776
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 3970 16785 3976 16788
rect 3954 16779 3976 16785
rect 3954 16745 3966 16779
rect 3954 16739 3976 16745
rect 3970 16736 3976 16739
rect 4028 16736 4034 16788
rect 4062 16736 4068 16788
rect 4120 16776 4126 16788
rect 12710 16776 12716 16788
rect 4120 16748 4165 16776
rect 12671 16748 12716 16776
rect 4120 16736 4126 16748
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 18325 16779 18383 16785
rect 18325 16745 18337 16779
rect 18371 16776 18383 16779
rect 18598 16776 18604 16788
rect 18371 16748 18604 16776
rect 18371 16745 18383 16748
rect 18325 16739 18383 16745
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 23382 16776 23388 16788
rect 23343 16748 23388 16776
rect 23382 16736 23388 16748
rect 23440 16736 23446 16788
rect 27614 16776 27620 16788
rect 26620 16748 27620 16776
rect 8386 16668 8392 16720
rect 8444 16708 8450 16720
rect 15930 16708 15936 16720
rect 8444 16680 15936 16708
rect 8444 16668 8450 16680
rect 15930 16668 15936 16680
rect 15988 16668 15994 16720
rect 17221 16711 17279 16717
rect 17221 16677 17233 16711
rect 17267 16708 17279 16711
rect 18414 16708 18420 16720
rect 17267 16680 18420 16708
rect 17267 16677 17279 16680
rect 17221 16671 17279 16677
rect 18414 16668 18420 16680
rect 18472 16668 18478 16720
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4614 16640 4620 16652
rect 4203 16612 4620 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 9122 16640 9128 16652
rect 9083 16612 9128 16640
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16640 9738 16652
rect 9732 16612 10548 16640
rect 9732 16600 9738 16612
rect 2498 16532 2504 16584
rect 2556 16572 2562 16584
rect 2593 16575 2651 16581
rect 2593 16572 2605 16575
rect 2556 16544 2605 16572
rect 2556 16532 2562 16544
rect 2593 16541 2605 16544
rect 2639 16541 2651 16575
rect 2593 16535 2651 16541
rect 2866 16532 2872 16584
rect 2924 16572 2930 16584
rect 3789 16575 3847 16581
rect 3789 16572 3801 16575
rect 2924 16544 3801 16572
rect 2924 16532 2930 16544
rect 3789 16541 3801 16544
rect 3835 16541 3847 16575
rect 7742 16572 7748 16584
rect 7703 16544 7748 16572
rect 3789 16535 3847 16541
rect 7742 16532 7748 16544
rect 7800 16532 7806 16584
rect 10520 16572 10548 16612
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 12713 16643 12771 16649
rect 12713 16640 12725 16643
rect 12676 16612 12725 16640
rect 12676 16600 12682 16612
rect 12713 16609 12725 16612
rect 12759 16609 12771 16643
rect 18322 16640 18328 16652
rect 18235 16612 18328 16640
rect 12713 16603 12771 16609
rect 18322 16600 18328 16612
rect 18380 16640 18386 16652
rect 18966 16640 18972 16652
rect 18380 16612 18972 16640
rect 18380 16600 18386 16612
rect 18966 16600 18972 16612
rect 19024 16600 19030 16652
rect 19889 16643 19947 16649
rect 19889 16609 19901 16643
rect 19935 16640 19947 16643
rect 19978 16640 19984 16652
rect 19935 16612 19984 16640
rect 19935 16609 19947 16612
rect 19889 16603 19947 16609
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 20165 16643 20223 16649
rect 20165 16609 20177 16643
rect 20211 16640 20223 16643
rect 20254 16640 20260 16652
rect 20211 16612 20260 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 23293 16643 23351 16649
rect 23293 16609 23305 16643
rect 23339 16640 23351 16643
rect 23474 16640 23480 16652
rect 23339 16612 23480 16640
rect 23339 16609 23351 16612
rect 23293 16603 23351 16609
rect 23474 16600 23480 16612
rect 23532 16600 23538 16652
rect 26620 16649 26648 16748
rect 27614 16736 27620 16748
rect 27672 16776 27678 16788
rect 28537 16779 28595 16785
rect 28537 16776 28549 16779
rect 27672 16748 28549 16776
rect 27672 16736 27678 16748
rect 28537 16745 28549 16748
rect 28583 16776 28595 16779
rect 31202 16776 31208 16788
rect 28583 16748 31208 16776
rect 28583 16745 28595 16748
rect 28537 16739 28595 16745
rect 31202 16736 31208 16748
rect 31260 16736 31266 16788
rect 34698 16736 34704 16788
rect 34756 16776 34762 16788
rect 35253 16779 35311 16785
rect 35253 16776 35265 16779
rect 34756 16748 35265 16776
rect 34756 16736 34762 16748
rect 35253 16745 35265 16748
rect 35299 16776 35311 16779
rect 35526 16776 35532 16788
rect 35299 16748 35532 16776
rect 35299 16745 35311 16748
rect 35253 16739 35311 16745
rect 35526 16736 35532 16748
rect 35584 16736 35590 16788
rect 30469 16711 30527 16717
rect 30469 16677 30481 16711
rect 30515 16708 30527 16711
rect 30650 16708 30656 16720
rect 30515 16680 30656 16708
rect 30515 16677 30527 16680
rect 30469 16671 30527 16677
rect 30650 16668 30656 16680
rect 30708 16668 30714 16720
rect 26605 16643 26663 16649
rect 26605 16609 26617 16643
rect 26651 16609 26663 16643
rect 26605 16603 26663 16609
rect 35618 16600 35624 16652
rect 35676 16640 35682 16652
rect 35805 16643 35863 16649
rect 35805 16640 35817 16643
rect 35676 16612 35817 16640
rect 35676 16600 35682 16612
rect 35805 16609 35817 16612
rect 35851 16609 35863 16643
rect 35805 16603 35863 16609
rect 12897 16575 12955 16581
rect 10520 16544 12756 16572
rect 2406 16464 2412 16516
rect 2464 16504 2470 16516
rect 2777 16507 2835 16513
rect 2777 16504 2789 16507
rect 2464 16476 2789 16504
rect 2464 16464 2470 16476
rect 2777 16473 2789 16476
rect 2823 16473 2835 16507
rect 2777 16467 2835 16473
rect 4525 16507 4583 16513
rect 4525 16473 4537 16507
rect 4571 16504 4583 16507
rect 8202 16504 8208 16516
rect 4571 16476 8208 16504
rect 4571 16473 4583 16476
rect 4525 16467 4583 16473
rect 8202 16464 8208 16476
rect 8260 16464 8266 16516
rect 9309 16507 9367 16513
rect 9309 16473 9321 16507
rect 9355 16504 9367 16507
rect 9398 16504 9404 16516
rect 9355 16476 9404 16504
rect 9355 16473 9367 16476
rect 9309 16467 9367 16473
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 12434 16464 12440 16516
rect 12492 16504 12498 16516
rect 12621 16507 12679 16513
rect 12621 16504 12633 16507
rect 12492 16476 12633 16504
rect 12492 16464 12498 16476
rect 12621 16473 12633 16476
rect 12667 16473 12679 16507
rect 12728 16504 12756 16544
rect 12897 16541 12909 16575
rect 12943 16572 12955 16575
rect 12986 16572 12992 16584
rect 12943 16544 12992 16572
rect 12943 16541 12955 16544
rect 12897 16535 12955 16541
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 18138 16572 18144 16584
rect 18099 16544 18144 16572
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16572 18475 16575
rect 18506 16572 18512 16584
rect 18463 16544 18512 16572
rect 18463 16541 18475 16544
rect 18417 16535 18475 16541
rect 18506 16532 18512 16544
rect 18564 16532 18570 16584
rect 23106 16572 23112 16584
rect 23067 16544 23112 16572
rect 23106 16532 23112 16544
rect 23164 16532 23170 16584
rect 23198 16532 23204 16584
rect 23256 16572 23262 16584
rect 26878 16581 26884 16584
rect 23385 16575 23443 16581
rect 23385 16572 23397 16575
rect 23256 16544 23397 16572
rect 23256 16532 23262 16544
rect 23385 16541 23397 16544
rect 23431 16541 23443 16575
rect 23385 16535 23443 16541
rect 26872 16535 26884 16581
rect 26936 16572 26942 16584
rect 30101 16575 30159 16581
rect 30101 16572 30113 16575
rect 26936 16544 26972 16572
rect 29564 16544 30113 16572
rect 26878 16532 26884 16535
rect 26936 16532 26942 16544
rect 15102 16504 15108 16516
rect 12728 16476 15108 16504
rect 12621 16467 12679 16473
rect 15102 16464 15108 16476
rect 15160 16464 15166 16516
rect 17037 16507 17095 16513
rect 17037 16504 17049 16507
rect 16408 16476 17049 16504
rect 7558 16436 7564 16448
rect 7519 16408 7564 16436
rect 7558 16396 7564 16408
rect 7616 16396 7622 16448
rect 13078 16436 13084 16448
rect 13039 16408 13084 16436
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 16206 16396 16212 16448
rect 16264 16436 16270 16448
rect 16408 16445 16436 16476
rect 17037 16473 17049 16476
rect 17083 16473 17095 16507
rect 17037 16467 17095 16473
rect 16393 16439 16451 16445
rect 16393 16436 16405 16439
rect 16264 16408 16405 16436
rect 16264 16396 16270 16408
rect 16393 16405 16405 16408
rect 16439 16405 16451 16439
rect 18598 16436 18604 16448
rect 18559 16408 18604 16436
rect 16393 16399 16451 16405
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 23569 16439 23627 16445
rect 23569 16405 23581 16439
rect 23615 16436 23627 16439
rect 24854 16436 24860 16448
rect 23615 16408 24860 16436
rect 23615 16405 23627 16408
rect 23569 16399 23627 16405
rect 24854 16396 24860 16408
rect 24912 16396 24918 16448
rect 27706 16396 27712 16448
rect 27764 16436 27770 16448
rect 27985 16439 28043 16445
rect 27985 16436 27997 16439
rect 27764 16408 27997 16436
rect 27764 16396 27770 16408
rect 27985 16405 27997 16408
rect 28031 16405 28043 16439
rect 27985 16399 28043 16405
rect 29086 16396 29092 16448
rect 29144 16436 29150 16448
rect 29564 16445 29592 16544
rect 30101 16541 30113 16544
rect 30147 16541 30159 16575
rect 30282 16572 30288 16584
rect 30243 16544 30288 16572
rect 30101 16535 30159 16541
rect 30282 16532 30288 16544
rect 30340 16532 30346 16584
rect 36072 16507 36130 16513
rect 36072 16473 36084 16507
rect 36118 16504 36130 16507
rect 36262 16504 36268 16516
rect 36118 16476 36268 16504
rect 36118 16473 36130 16476
rect 36072 16467 36130 16473
rect 36262 16464 36268 16476
rect 36320 16464 36326 16516
rect 29549 16439 29607 16445
rect 29549 16436 29561 16439
rect 29144 16408 29561 16436
rect 29144 16396 29150 16408
rect 29549 16405 29561 16408
rect 29595 16405 29607 16439
rect 37182 16436 37188 16448
rect 37143 16408 37188 16436
rect 29549 16399 29607 16405
rect 37182 16396 37188 16408
rect 37240 16396 37246 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 9398 16232 9404 16244
rect 9359 16204 9404 16232
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 27157 16235 27215 16241
rect 27157 16201 27169 16235
rect 27203 16232 27215 16235
rect 27246 16232 27252 16244
rect 27203 16204 27252 16232
rect 27203 16201 27215 16204
rect 27157 16195 27215 16201
rect 27246 16192 27252 16204
rect 27304 16192 27310 16244
rect 27706 16192 27712 16244
rect 27764 16232 27770 16244
rect 28445 16235 28503 16241
rect 28445 16232 28457 16235
rect 27764 16204 28457 16232
rect 27764 16192 27770 16204
rect 28445 16201 28457 16204
rect 28491 16201 28503 16235
rect 36262 16232 36268 16244
rect 36223 16204 36268 16232
rect 28445 16195 28503 16201
rect 36262 16192 36268 16204
rect 36320 16192 36326 16244
rect 27798 16124 27804 16176
rect 27856 16164 27862 16176
rect 28353 16167 28411 16173
rect 28353 16164 28365 16167
rect 27856 16136 28365 16164
rect 27856 16124 27862 16136
rect 28353 16133 28365 16136
rect 28399 16133 28411 16167
rect 28353 16127 28411 16133
rect 35161 16167 35219 16173
rect 35161 16133 35173 16167
rect 35207 16164 35219 16167
rect 36078 16164 36084 16176
rect 35207 16136 35848 16164
rect 35207 16133 35219 16136
rect 35161 16127 35219 16133
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16096 1458 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 1452 16068 2053 16096
rect 1452 16056 1458 16068
rect 2041 16065 2053 16068
rect 2087 16065 2099 16099
rect 3142 16096 3148 16108
rect 3103 16068 3148 16096
rect 2041 16059 2099 16065
rect 3142 16056 3148 16068
rect 3200 16056 3206 16108
rect 6546 16096 6552 16108
rect 6507 16068 6552 16096
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 9582 16096 9588 16108
rect 9543 16068 9588 16096
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 12894 16096 12900 16108
rect 12855 16068 12900 16096
rect 12894 16056 12900 16068
rect 12952 16056 12958 16108
rect 15930 16056 15936 16108
rect 15988 16096 15994 16108
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 15988 16068 16681 16096
rect 15988 16056 15994 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16942 16096 16948 16108
rect 16903 16068 16948 16096
rect 16669 16059 16727 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16096 17831 16099
rect 17862 16096 17868 16108
rect 17819 16068 17868 16096
rect 17819 16065 17831 16068
rect 17773 16059 17831 16065
rect 17862 16056 17868 16068
rect 17920 16056 17926 16108
rect 24854 16096 24860 16108
rect 24815 16068 24860 16096
rect 24854 16056 24860 16068
rect 24912 16056 24918 16108
rect 27341 16099 27399 16105
rect 27341 16065 27353 16099
rect 27387 16096 27399 16099
rect 27387 16068 28028 16096
rect 27387 16065 27399 16068
rect 27341 16059 27399 16065
rect 16853 16031 16911 16037
rect 16853 15997 16865 16031
rect 16899 16028 16911 16031
rect 18322 16028 18328 16040
rect 16899 16000 18328 16028
rect 16899 15997 16911 16000
rect 16853 15991 16911 15997
rect 18322 15988 18328 16000
rect 18380 15988 18386 16040
rect 22554 16028 22560 16040
rect 22515 16000 22560 16028
rect 22554 15988 22560 16000
rect 22612 15988 22618 16040
rect 22741 16031 22799 16037
rect 22741 15997 22753 16031
rect 22787 16028 22799 16031
rect 23198 16028 23204 16040
rect 22787 16000 23204 16028
rect 22787 15997 22799 16000
rect 22741 15991 22799 15997
rect 23198 15988 23204 16000
rect 23256 15988 23262 16040
rect 23474 16028 23480 16040
rect 23435 16000 23480 16028
rect 23474 15988 23480 16000
rect 23532 15988 23538 16040
rect 27525 16031 27583 16037
rect 27525 15997 27537 16031
rect 27571 15997 27583 16031
rect 27525 15991 27583 15997
rect 3237 15963 3295 15969
rect 3237 15929 3249 15963
rect 3283 15960 3295 15963
rect 4614 15960 4620 15972
rect 3283 15932 4620 15960
rect 3283 15929 3295 15932
rect 3237 15923 3295 15929
rect 4614 15920 4620 15932
rect 4672 15920 4678 15972
rect 17954 15960 17960 15972
rect 17915 15932 17960 15960
rect 17954 15920 17960 15932
rect 18012 15920 18018 15972
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 2498 15892 2504 15904
rect 1627 15864 2504 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 6362 15892 6368 15904
rect 6323 15864 6368 15892
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 12710 15892 12716 15904
rect 12671 15864 12716 15892
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 13262 15852 13268 15904
rect 13320 15892 13326 15904
rect 13357 15895 13415 15901
rect 13357 15892 13369 15895
rect 13320 15864 13369 15892
rect 13320 15852 13326 15864
rect 13357 15861 13369 15864
rect 13403 15892 13415 15895
rect 13814 15892 13820 15904
rect 13403 15864 13820 15892
rect 13403 15861 13415 15864
rect 13357 15855 13415 15861
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 16850 15892 16856 15904
rect 16811 15864 16856 15892
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 17129 15895 17187 15901
rect 17129 15861 17141 15895
rect 17175 15892 17187 15895
rect 17402 15892 17408 15904
rect 17175 15864 17408 15892
rect 17175 15861 17187 15864
rect 17129 15855 17187 15861
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 20806 15892 20812 15904
rect 20767 15864 20812 15892
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 25041 15895 25099 15901
rect 25041 15861 25053 15895
rect 25087 15892 25099 15895
rect 26050 15892 26056 15904
rect 25087 15864 26056 15892
rect 25087 15861 25099 15864
rect 25041 15855 25099 15861
rect 26050 15852 26056 15864
rect 26108 15852 26114 15904
rect 27540 15892 27568 15991
rect 28000 15969 28028 16068
rect 32490 16056 32496 16108
rect 32548 16096 32554 16108
rect 34885 16099 34943 16105
rect 34885 16096 34897 16099
rect 32548 16068 34897 16096
rect 32548 16056 32554 16068
rect 34885 16065 34897 16068
rect 34931 16065 34943 16099
rect 34885 16059 34943 16065
rect 28629 16031 28687 16037
rect 28629 15997 28641 16031
rect 28675 16028 28687 16031
rect 30190 16028 30196 16040
rect 28675 16000 30196 16028
rect 28675 15997 28687 16000
rect 28629 15991 28687 15997
rect 30190 15988 30196 16000
rect 30248 15988 30254 16040
rect 27985 15963 28043 15969
rect 27985 15929 27997 15963
rect 28031 15929 28043 15963
rect 34900 15960 34928 16059
rect 35526 16056 35532 16108
rect 35584 16096 35590 16108
rect 35820 16105 35848 16136
rect 35912 16136 36084 16164
rect 35912 16105 35940 16136
rect 36078 16124 36084 16136
rect 36136 16164 36142 16176
rect 36446 16164 36452 16176
rect 36136 16136 36452 16164
rect 36136 16124 36142 16136
rect 36446 16124 36452 16136
rect 36504 16124 36510 16176
rect 35621 16099 35679 16105
rect 35621 16096 35633 16099
rect 35584 16068 35633 16096
rect 35584 16056 35590 16068
rect 35621 16065 35633 16068
rect 35667 16065 35679 16099
rect 35621 16059 35679 16065
rect 35805 16099 35863 16105
rect 35805 16065 35817 16099
rect 35851 16065 35863 16099
rect 35805 16059 35863 16065
rect 35897 16099 35955 16105
rect 35897 16065 35909 16099
rect 35943 16065 35955 16099
rect 35897 16059 35955 16065
rect 35989 16099 36047 16105
rect 35989 16065 36001 16099
rect 36035 16096 36047 16099
rect 37182 16096 37188 16108
rect 36035 16068 37188 16096
rect 36035 16065 36047 16068
rect 35989 16059 36047 16065
rect 35161 16031 35219 16037
rect 35161 15997 35173 16031
rect 35207 16028 35219 16031
rect 35912 16028 35940 16059
rect 35207 16000 35940 16028
rect 35207 15997 35219 16000
rect 35161 15991 35219 15997
rect 36004 15960 36032 16059
rect 37182 16056 37188 16068
rect 37240 16056 37246 16108
rect 34900 15932 36032 15960
rect 27985 15923 28043 15929
rect 29086 15892 29092 15904
rect 27540 15864 29092 15892
rect 29086 15852 29092 15864
rect 29144 15852 29150 15904
rect 34977 15895 35035 15901
rect 34977 15861 34989 15895
rect 35023 15892 35035 15895
rect 35342 15892 35348 15904
rect 35023 15864 35348 15892
rect 35023 15861 35035 15864
rect 34977 15855 35035 15861
rect 35342 15852 35348 15864
rect 35400 15852 35406 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 16942 15688 16948 15700
rect 13188 15660 16948 15688
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 13078 15552 13084 15564
rect 5767 15524 13084 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 13078 15512 13084 15524
rect 13136 15512 13142 15564
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 5445 15487 5503 15493
rect 5445 15484 5457 15487
rect 4212 15456 5457 15484
rect 4212 15444 4218 15456
rect 5445 15453 5457 15456
rect 5491 15453 5503 15487
rect 6178 15484 6184 15496
rect 6139 15456 6184 15484
rect 5445 15447 5503 15453
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 7374 15444 7380 15496
rect 7432 15484 7438 15496
rect 7469 15487 7527 15493
rect 7469 15484 7481 15487
rect 7432 15456 7481 15484
rect 7432 15444 7438 15456
rect 7469 15453 7481 15456
rect 7515 15453 7527 15487
rect 7469 15447 7527 15453
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8720 15456 8953 15484
rect 8720 15444 8726 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 12526 15444 12532 15496
rect 12584 15484 12590 15496
rect 12621 15487 12679 15493
rect 12621 15484 12633 15487
rect 12584 15456 12633 15484
rect 12584 15444 12590 15456
rect 12621 15453 12633 15456
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 4614 15376 4620 15428
rect 4672 15416 4678 15428
rect 13188 15416 13216 15660
rect 16206 15620 16212 15632
rect 16167 15592 16212 15620
rect 16206 15580 16212 15592
rect 16264 15580 16270 15632
rect 16316 15561 16344 15660
rect 16942 15648 16948 15660
rect 17000 15648 17006 15700
rect 17313 15691 17371 15697
rect 17313 15657 17325 15691
rect 17359 15688 17371 15691
rect 18046 15688 18052 15700
rect 17359 15660 18052 15688
rect 17359 15657 17371 15660
rect 17313 15651 17371 15657
rect 18046 15648 18052 15660
rect 18104 15688 18110 15700
rect 18322 15688 18328 15700
rect 18104 15660 18328 15688
rect 18104 15648 18110 15660
rect 18322 15648 18328 15660
rect 18380 15648 18386 15700
rect 23198 15688 23204 15700
rect 23159 15660 23204 15688
rect 23198 15648 23204 15660
rect 23256 15648 23262 15700
rect 32674 15688 32680 15700
rect 32635 15660 32680 15688
rect 32674 15648 32680 15660
rect 32732 15648 32738 15700
rect 35805 15691 35863 15697
rect 35805 15657 35817 15691
rect 35851 15688 35863 15691
rect 35894 15688 35900 15700
rect 35851 15660 35900 15688
rect 35851 15657 35863 15660
rect 35805 15651 35863 15657
rect 35894 15648 35900 15660
rect 35952 15648 35958 15700
rect 36078 15688 36084 15700
rect 36039 15660 36084 15688
rect 36078 15648 36084 15660
rect 36136 15648 36142 15700
rect 24670 15620 24676 15632
rect 22204 15592 24676 15620
rect 22204 15564 22232 15592
rect 24670 15580 24676 15592
rect 24728 15580 24734 15632
rect 16301 15555 16359 15561
rect 16301 15521 16313 15555
rect 16347 15521 16359 15555
rect 16301 15515 16359 15521
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18693 15555 18751 15561
rect 18693 15552 18705 15555
rect 18012 15524 18705 15552
rect 18012 15512 18018 15524
rect 18693 15521 18705 15524
rect 18739 15552 18751 15555
rect 19245 15555 19303 15561
rect 19245 15552 19257 15555
rect 18739 15524 19257 15552
rect 18739 15521 18751 15524
rect 18693 15515 18751 15521
rect 19245 15521 19257 15524
rect 19291 15521 19303 15555
rect 20806 15552 20812 15564
rect 20767 15524 20812 15552
rect 19245 15515 19303 15521
rect 20806 15512 20812 15524
rect 20864 15512 20870 15564
rect 22186 15552 22192 15564
rect 22147 15524 22192 15552
rect 22186 15512 22192 15524
rect 22244 15512 22250 15564
rect 23842 15512 23848 15564
rect 23900 15552 23906 15564
rect 25133 15555 25191 15561
rect 25133 15552 25145 15555
rect 23900 15524 25145 15552
rect 23900 15512 23906 15524
rect 25133 15521 25145 15524
rect 25179 15521 25191 15555
rect 35802 15552 35808 15564
rect 35763 15524 35808 15552
rect 25133 15515 25191 15521
rect 35802 15512 35808 15524
rect 35860 15512 35866 15564
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 13449 15487 13507 15493
rect 13320 15456 13365 15484
rect 13320 15444 13326 15456
rect 13449 15453 13461 15487
rect 13495 15453 13507 15487
rect 15930 15484 15936 15496
rect 15891 15456 15936 15484
rect 13449 15447 13507 15453
rect 4672 15388 13216 15416
rect 4672 15376 4678 15388
rect 13354 15376 13360 15428
rect 13412 15416 13418 15428
rect 13464 15416 13492 15447
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 16080 15487 16138 15493
rect 16080 15453 16092 15487
rect 16126 15484 16138 15487
rect 17129 15487 17187 15493
rect 17129 15484 17141 15487
rect 16126 15453 16160 15484
rect 16080 15447 16160 15453
rect 16132 15416 16160 15447
rect 16592 15456 17141 15484
rect 16592 15416 16620 15456
rect 17129 15453 17141 15456
rect 17175 15453 17187 15487
rect 17129 15447 17187 15453
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 19484 15456 19533 15484
rect 19484 15444 19490 15456
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 22922 15444 22928 15496
rect 22980 15484 22986 15496
rect 23385 15487 23443 15493
rect 23385 15484 23397 15487
rect 22980 15456 23397 15484
rect 22980 15444 22986 15456
rect 23385 15453 23397 15456
rect 23431 15453 23443 15487
rect 25406 15484 25412 15496
rect 25367 15456 25412 15484
rect 23385 15447 23443 15453
rect 25406 15444 25412 15456
rect 25464 15444 25470 15496
rect 29730 15444 29736 15496
rect 29788 15484 29794 15496
rect 30009 15487 30067 15493
rect 30009 15484 30021 15487
rect 29788 15456 30021 15484
rect 29788 15444 29794 15456
rect 30009 15453 30021 15456
rect 30055 15453 30067 15487
rect 30009 15447 30067 15453
rect 32214 15444 32220 15496
rect 32272 15484 32278 15496
rect 32493 15487 32551 15493
rect 32493 15484 32505 15487
rect 32272 15456 32505 15484
rect 32272 15444 32278 15456
rect 32493 15453 32505 15456
rect 32539 15453 32551 15487
rect 32493 15447 32551 15453
rect 35434 15444 35440 15496
rect 35492 15484 35498 15496
rect 35713 15487 35771 15493
rect 35713 15484 35725 15487
rect 35492 15456 35725 15484
rect 35492 15444 35498 15456
rect 35713 15453 35725 15456
rect 35759 15453 35771 15487
rect 35713 15447 35771 15453
rect 13412 15388 13492 15416
rect 15212 15388 16620 15416
rect 16669 15419 16727 15425
rect 13412 15376 13418 15388
rect 12161 15351 12219 15357
rect 12161 15317 12173 15351
rect 12207 15348 12219 15351
rect 13372 15348 13400 15376
rect 12207 15320 13400 15348
rect 13449 15351 13507 15357
rect 12207 15317 12219 15320
rect 12161 15311 12219 15317
rect 13449 15317 13461 15351
rect 13495 15348 13507 15351
rect 15212 15348 15240 15388
rect 16669 15385 16681 15419
rect 16715 15416 16727 15419
rect 20714 15416 20720 15428
rect 16715 15388 20720 15416
rect 16715 15385 16727 15388
rect 16669 15379 16727 15385
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 20990 15416 20996 15428
rect 20951 15388 20996 15416
rect 20990 15376 20996 15388
rect 21048 15376 21054 15428
rect 30190 15416 30196 15428
rect 30151 15388 30196 15416
rect 30190 15376 30196 15388
rect 30248 15376 30254 15428
rect 13495 15320 15240 15348
rect 13495 15317 13507 15320
rect 13449 15311 13507 15317
rect 15286 15308 15292 15360
rect 15344 15348 15350 15360
rect 15381 15351 15439 15357
rect 15381 15348 15393 15351
rect 15344 15320 15393 15348
rect 15344 15308 15350 15320
rect 15381 15317 15393 15320
rect 15427 15348 15439 15351
rect 16206 15348 16212 15360
rect 15427 15320 16212 15348
rect 15427 15317 15439 15320
rect 15381 15311 15439 15317
rect 16206 15308 16212 15320
rect 16264 15308 16270 15360
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 17862 15348 17868 15360
rect 16908 15320 17868 15348
rect 16908 15308 16914 15320
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 27798 15348 27804 15360
rect 27759 15320 27804 15348
rect 27798 15308 27804 15320
rect 27856 15308 27862 15360
rect 28445 15351 28503 15357
rect 28445 15317 28457 15351
rect 28491 15348 28503 15351
rect 29086 15348 29092 15360
rect 28491 15320 29092 15348
rect 28491 15317 28503 15320
rect 28445 15311 28503 15317
rect 29086 15308 29092 15320
rect 29144 15308 29150 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 9582 15104 9588 15156
rect 9640 15144 9646 15156
rect 9677 15147 9735 15153
rect 9677 15144 9689 15147
rect 9640 15116 9689 15144
rect 9640 15104 9646 15116
rect 9677 15113 9689 15116
rect 9723 15113 9735 15147
rect 9677 15107 9735 15113
rect 19705 15147 19763 15153
rect 19705 15113 19717 15147
rect 19751 15144 19763 15147
rect 19978 15144 19984 15156
rect 19751 15116 19984 15144
rect 19751 15113 19763 15116
rect 19705 15107 19763 15113
rect 19978 15104 19984 15116
rect 20036 15104 20042 15156
rect 20533 15147 20591 15153
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 20990 15144 20996 15156
rect 20579 15116 20996 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 25406 15104 25412 15156
rect 25464 15144 25470 15156
rect 29730 15144 29736 15156
rect 25464 15116 26234 15144
rect 29691 15116 29736 15144
rect 25464 15104 25470 15116
rect 4154 15076 4160 15088
rect 4115 15048 4160 15076
rect 4154 15036 4160 15048
rect 4212 15036 4218 15088
rect 7558 15076 7564 15088
rect 7519 15048 7564 15076
rect 7558 15036 7564 15048
rect 7616 15036 7622 15088
rect 10134 15076 10140 15088
rect 10095 15048 10140 15076
rect 10134 15036 10140 15048
rect 10192 15036 10198 15088
rect 12710 15076 12716 15088
rect 12671 15048 12716 15076
rect 12710 15036 12716 15048
rect 12768 15036 12774 15088
rect 18601 15079 18659 15085
rect 18601 15045 18613 15079
rect 18647 15076 18659 15079
rect 24394 15076 24400 15088
rect 18647 15048 22094 15076
rect 24355 15048 24400 15076
rect 18647 15045 18659 15048
rect 18601 15039 18659 15045
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 15008 1458 15020
rect 2041 15011 2099 15017
rect 2041 15008 2053 15011
rect 1452 14980 2053 15008
rect 1452 14968 1458 14980
rect 2041 14977 2053 14980
rect 2087 14977 2099 15011
rect 7374 15008 7380 15020
rect 7335 14980 7380 15008
rect 2041 14971 2099 14977
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 9490 14968 9496 15020
rect 9548 15008 9554 15020
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 9548 14980 9873 15008
rect 9548 14968 9554 14980
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 12526 15008 12532 15020
rect 12487 14980 12532 15008
rect 9861 14971 9919 14977
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 19245 15011 19303 15017
rect 19245 14977 19257 15011
rect 19291 14977 19303 15011
rect 19245 14971 19303 14977
rect 19521 15011 19579 15017
rect 19521 14977 19533 15011
rect 19567 15008 19579 15011
rect 19610 15008 19616 15020
rect 19567 14980 19616 15008
rect 19567 14977 19579 14980
rect 19521 14971 19579 14977
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 3973 14943 4031 14949
rect 3973 14940 3985 14943
rect 3292 14912 3985 14940
rect 3292 14900 3298 14912
rect 3973 14909 3985 14912
rect 4019 14909 4031 14943
rect 4433 14943 4491 14949
rect 4433 14940 4445 14943
rect 3973 14903 4031 14909
rect 4080 14912 4445 14940
rect 4080 14884 4108 14912
rect 4433 14909 4445 14912
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 7837 14943 7895 14949
rect 7837 14909 7849 14943
rect 7883 14909 7895 14943
rect 10042 14940 10048 14952
rect 10003 14912 10048 14940
rect 7837 14903 7895 14909
rect 4062 14832 4068 14884
rect 4120 14832 4126 14884
rect 7852 14872 7880 14903
rect 10042 14900 10048 14912
rect 10100 14900 10106 14952
rect 12986 14940 12992 14952
rect 12947 14912 12992 14940
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14940 16175 14943
rect 16761 14943 16819 14949
rect 16761 14940 16773 14943
rect 16163 14912 16773 14940
rect 16163 14909 16175 14912
rect 16117 14903 16175 14909
rect 16761 14909 16773 14912
rect 16807 14909 16819 14943
rect 16942 14940 16948 14952
rect 16903 14912 16948 14940
rect 16761 14903 16819 14909
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 9766 14872 9772 14884
rect 7852 14844 9772 14872
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 2774 14804 2780 14816
rect 1627 14776 2780 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 2774 14764 2780 14776
rect 2832 14764 2838 14816
rect 3878 14764 3884 14816
rect 3936 14804 3942 14816
rect 7852 14804 7880 14844
rect 9766 14832 9772 14844
rect 9824 14832 9830 14884
rect 19260 14872 19288 14971
rect 19610 14968 19616 14980
rect 19668 14968 19674 15020
rect 19794 14968 19800 15020
rect 19852 15008 19858 15020
rect 20349 15011 20407 15017
rect 20349 15008 20361 15011
rect 19852 14980 20361 15008
rect 19852 14968 19858 14980
rect 20349 14977 20361 14980
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 19426 14940 19432 14952
rect 19387 14912 19432 14940
rect 19426 14900 19432 14912
rect 19484 14900 19490 14952
rect 22066 14940 22094 15048
rect 24394 15036 24400 15048
rect 24452 15036 24458 15088
rect 26050 15076 26056 15088
rect 26011 15048 26056 15076
rect 26050 15036 26056 15048
rect 26108 15036 26114 15088
rect 26206 15076 26234 15116
rect 29730 15104 29736 15116
rect 29788 15104 29794 15156
rect 27157 15079 27215 15085
rect 27157 15076 27169 15079
rect 26206 15048 27169 15076
rect 27157 15045 27169 15048
rect 27203 15045 27215 15079
rect 27157 15039 27215 15045
rect 28813 15079 28871 15085
rect 28813 15045 28825 15079
rect 28859 15076 28871 15079
rect 29270 15076 29276 15088
rect 28859 15048 29276 15076
rect 28859 15045 28871 15048
rect 28813 15039 28871 15045
rect 29270 15036 29276 15048
rect 29328 15036 29334 15088
rect 35437 15079 35495 15085
rect 35437 15045 35449 15079
rect 35483 15076 35495 15079
rect 35894 15076 35900 15088
rect 35483 15048 35900 15076
rect 35483 15045 35495 15048
rect 35437 15039 35495 15045
rect 35894 15036 35900 15048
rect 35952 15076 35958 15088
rect 36446 15076 36452 15088
rect 35952 15048 36452 15076
rect 35952 15036 35958 15048
rect 36446 15036 36452 15048
rect 36504 15036 36510 15088
rect 22554 14968 22560 15020
rect 22612 15008 22618 15020
rect 22649 15011 22707 15017
rect 22649 15008 22661 15011
rect 22612 14980 22661 15008
rect 22612 14968 22618 14980
rect 22649 14977 22661 14980
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 34790 14968 34796 15020
rect 34848 15008 34854 15020
rect 35253 15011 35311 15017
rect 35253 15008 35265 15011
rect 34848 14980 35265 15008
rect 34848 14968 34854 14980
rect 35253 14977 35265 14980
rect 35299 14977 35311 15011
rect 35526 15008 35532 15020
rect 35487 14980 35532 15008
rect 35253 14971 35311 14977
rect 35526 14968 35532 14980
rect 35584 14968 35590 15020
rect 22186 14940 22192 14952
rect 22066 14912 22192 14940
rect 22186 14900 22192 14912
rect 22244 14900 22250 14952
rect 26237 14943 26295 14949
rect 26237 14909 26249 14943
rect 26283 14909 26295 14943
rect 26237 14903 26295 14909
rect 26973 14943 27031 14949
rect 26973 14909 26985 14943
rect 27019 14940 27031 14943
rect 27890 14940 27896 14952
rect 27019 14912 27896 14940
rect 27019 14909 27031 14912
rect 26973 14903 27031 14909
rect 19518 14872 19524 14884
rect 19260 14844 19524 14872
rect 19518 14832 19524 14844
rect 19576 14872 19582 14884
rect 20530 14872 20536 14884
rect 19576 14844 20536 14872
rect 19576 14832 19582 14844
rect 20530 14832 20536 14844
rect 20588 14832 20594 14884
rect 26252 14872 26280 14903
rect 27890 14900 27896 14912
rect 27948 14900 27954 14952
rect 30374 14872 30380 14884
rect 26252 14844 30380 14872
rect 30374 14832 30380 14844
rect 30432 14832 30438 14884
rect 35253 14875 35311 14881
rect 35253 14841 35265 14875
rect 35299 14872 35311 14875
rect 35342 14872 35348 14884
rect 35299 14844 35348 14872
rect 35299 14841 35311 14844
rect 35253 14835 35311 14841
rect 35342 14832 35348 14844
rect 35400 14832 35406 14884
rect 3936 14776 7880 14804
rect 3936 14764 3942 14776
rect 9306 14764 9312 14816
rect 9364 14804 9370 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9364 14776 9873 14804
rect 9364 14764 9370 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 19334 14804 19340 14816
rect 19295 14776 19340 14804
rect 9861 14767 9919 14773
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 3234 14600 3240 14612
rect 3195 14572 3240 14600
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 9306 14560 9312 14612
rect 9364 14600 9370 14612
rect 9401 14603 9459 14609
rect 9401 14600 9413 14603
rect 9364 14572 9413 14600
rect 9364 14560 9370 14572
rect 9401 14569 9413 14572
rect 9447 14600 9459 14603
rect 10321 14603 10379 14609
rect 10321 14600 10333 14603
rect 9447 14572 10333 14600
rect 9447 14569 9459 14572
rect 9401 14563 9459 14569
rect 10321 14569 10333 14572
rect 10367 14569 10379 14603
rect 19334 14600 19340 14612
rect 19295 14572 19340 14600
rect 10321 14563 10379 14569
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 19794 14600 19800 14612
rect 19755 14572 19800 14600
rect 19794 14560 19800 14572
rect 19852 14560 19858 14612
rect 33965 14603 34023 14609
rect 33965 14569 33977 14603
rect 34011 14600 34023 14603
rect 34330 14600 34336 14612
rect 34011 14572 34336 14600
rect 34011 14569 34023 14572
rect 33965 14563 34023 14569
rect 34330 14560 34336 14572
rect 34388 14600 34394 14612
rect 34885 14603 34943 14609
rect 34388 14572 34744 14600
rect 34388 14560 34394 14572
rect 3970 14492 3976 14544
rect 4028 14532 4034 14544
rect 4028 14504 6500 14532
rect 4028 14492 4034 14504
rect 5350 14464 5356 14476
rect 5311 14436 5356 14464
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 5997 14467 6055 14473
rect 5997 14433 6009 14467
rect 6043 14464 6055 14467
rect 6178 14464 6184 14476
rect 6043 14436 6184 14464
rect 6043 14433 6055 14436
rect 5997 14427 6055 14433
rect 6178 14424 6184 14436
rect 6236 14424 6242 14476
rect 6472 14473 6500 14504
rect 18598 14492 18604 14544
rect 18656 14532 18662 14544
rect 18656 14504 33824 14532
rect 18656 14492 18662 14504
rect 6457 14467 6515 14473
rect 6457 14433 6469 14467
rect 6503 14464 6515 14467
rect 9122 14464 9128 14476
rect 6503 14436 9128 14464
rect 6503 14433 6515 14436
rect 6457 14427 6515 14433
rect 9122 14424 9128 14436
rect 9180 14424 9186 14476
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 10042 14464 10048 14476
rect 9631 14436 10048 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 10042 14424 10048 14436
rect 10100 14464 10106 14476
rect 10505 14467 10563 14473
rect 10505 14464 10517 14467
rect 10100 14436 10517 14464
rect 10100 14424 10106 14436
rect 10505 14433 10517 14436
rect 10551 14464 10563 14467
rect 10594 14464 10600 14476
rect 10551 14436 10600 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 19426 14464 19432 14476
rect 19387 14436 19432 14464
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 22097 14467 22155 14473
rect 22097 14464 22109 14467
rect 19536 14436 22109 14464
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5166 14396 5172 14408
rect 5123 14368 5172 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 3988 14328 4016 14359
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14396 9459 14399
rect 9490 14396 9496 14408
rect 9447 14368 9496 14396
rect 9447 14365 9459 14368
rect 9401 14359 9459 14365
rect 9490 14356 9496 14368
rect 9548 14396 9554 14408
rect 10321 14399 10379 14405
rect 10321 14396 10333 14399
rect 9548 14368 10333 14396
rect 9548 14356 9554 14368
rect 10321 14365 10333 14368
rect 10367 14365 10379 14399
rect 10321 14359 10379 14365
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14396 15807 14399
rect 16209 14399 16267 14405
rect 16209 14396 16221 14399
rect 15795 14368 16221 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 16209 14365 16221 14368
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14396 18107 14399
rect 19536 14396 19564 14436
rect 22097 14433 22109 14436
rect 22143 14464 22155 14467
rect 23658 14464 23664 14476
rect 22143 14436 23664 14464
rect 22143 14433 22155 14436
rect 22097 14427 22155 14433
rect 23658 14424 23664 14436
rect 23716 14424 23722 14476
rect 27154 14464 27160 14476
rect 27115 14436 27160 14464
rect 27154 14424 27160 14436
rect 27212 14424 27218 14476
rect 30190 14424 30196 14476
rect 30248 14464 30254 14476
rect 30285 14467 30343 14473
rect 30285 14464 30297 14467
rect 30248 14436 30297 14464
rect 30248 14424 30254 14436
rect 30285 14433 30297 14436
rect 30331 14433 30343 14467
rect 30285 14427 30343 14433
rect 18095 14368 19564 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 19610 14356 19616 14408
rect 19668 14396 19674 14408
rect 19978 14396 19984 14408
rect 19668 14368 19984 14396
rect 19668 14356 19674 14368
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 21177 14399 21235 14405
rect 21177 14365 21189 14399
rect 21223 14396 21235 14399
rect 21637 14399 21695 14405
rect 21637 14396 21649 14399
rect 21223 14368 21649 14396
rect 21223 14365 21235 14368
rect 21177 14359 21235 14365
rect 21637 14365 21649 14368
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 26973 14399 27031 14405
rect 26973 14365 26985 14399
rect 27019 14396 27031 14399
rect 29270 14396 29276 14408
rect 27019 14368 29276 14396
rect 27019 14365 27031 14368
rect 26973 14359 27031 14365
rect 5350 14328 5356 14340
rect 3988 14300 5356 14328
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 6181 14331 6239 14337
rect 6181 14297 6193 14331
rect 6227 14328 6239 14331
rect 6362 14328 6368 14340
rect 6227 14300 6368 14328
rect 6227 14297 6239 14300
rect 6181 14291 6239 14297
rect 6362 14288 6368 14300
rect 6420 14288 6426 14340
rect 9677 14331 9735 14337
rect 9677 14297 9689 14331
rect 9723 14328 9735 14331
rect 10226 14328 10232 14340
rect 9723 14300 10232 14328
rect 9723 14297 9735 14300
rect 9677 14291 9735 14297
rect 10226 14288 10232 14300
rect 10284 14328 10290 14340
rect 10597 14331 10655 14337
rect 10597 14328 10609 14331
rect 10284 14300 10609 14328
rect 10284 14288 10290 14300
rect 10597 14297 10609 14300
rect 10643 14297 10655 14331
rect 10597 14291 10655 14297
rect 16393 14331 16451 14337
rect 16393 14297 16405 14331
rect 16439 14328 16451 14331
rect 17310 14328 17316 14340
rect 16439 14300 17316 14328
rect 16439 14297 16451 14300
rect 16393 14291 16451 14297
rect 17310 14288 17316 14300
rect 17368 14288 17374 14340
rect 18693 14331 18751 14337
rect 18693 14297 18705 14331
rect 18739 14328 18751 14331
rect 19242 14328 19248 14340
rect 18739 14300 19248 14328
rect 18739 14297 18751 14300
rect 18693 14291 18751 14297
rect 19242 14288 19248 14300
rect 19300 14328 19306 14340
rect 19337 14331 19395 14337
rect 19337 14328 19349 14331
rect 19300 14300 19349 14328
rect 19300 14288 19306 14300
rect 19337 14297 19349 14300
rect 19383 14328 19395 14331
rect 19518 14328 19524 14340
rect 19383 14300 19524 14328
rect 19383 14297 19395 14300
rect 19337 14291 19395 14297
rect 19518 14288 19524 14300
rect 19576 14288 19582 14340
rect 21818 14328 21824 14340
rect 21779 14300 21824 14328
rect 21818 14288 21824 14300
rect 21876 14288 21882 14340
rect 26988 14328 27016 14359
rect 29270 14356 29276 14368
rect 29328 14356 29334 14408
rect 30101 14399 30159 14405
rect 30101 14365 30113 14399
rect 30147 14396 30159 14399
rect 31846 14396 31852 14408
rect 30147 14368 31852 14396
rect 30147 14365 30159 14368
rect 30101 14359 30159 14365
rect 26160 14300 27016 14328
rect 28997 14331 29055 14337
rect 26160 14272 26188 14300
rect 28997 14297 29009 14331
rect 29043 14328 29055 14331
rect 29546 14328 29552 14340
rect 29043 14300 29552 14328
rect 29043 14297 29055 14300
rect 28997 14291 29055 14297
rect 29546 14288 29552 14300
rect 29604 14328 29610 14340
rect 30116 14328 30144 14359
rect 31846 14356 31852 14368
rect 31904 14356 31910 14408
rect 32214 14356 32220 14408
rect 32272 14396 32278 14408
rect 33796 14405 33824 14504
rect 34716 14473 34744 14572
rect 34885 14569 34897 14603
rect 34931 14600 34943 14603
rect 35526 14600 35532 14612
rect 34931 14572 35532 14600
rect 34931 14569 34943 14572
rect 34885 14563 34943 14569
rect 35526 14560 35532 14572
rect 35584 14560 35590 14612
rect 34701 14467 34759 14473
rect 34701 14433 34713 14467
rect 34747 14464 34759 14467
rect 36446 14464 36452 14476
rect 34747 14436 36452 14464
rect 34747 14433 34759 14436
rect 34701 14427 34759 14433
rect 36446 14424 36452 14436
rect 36504 14424 36510 14476
rect 33137 14399 33195 14405
rect 33137 14396 33149 14399
rect 32272 14368 33149 14396
rect 32272 14356 32278 14368
rect 33137 14365 33149 14368
rect 33183 14365 33195 14399
rect 33137 14359 33195 14365
rect 33321 14399 33379 14405
rect 33321 14365 33333 14399
rect 33367 14365 33379 14399
rect 33321 14359 33379 14365
rect 33781 14399 33839 14405
rect 33781 14365 33793 14399
rect 33827 14365 33839 14399
rect 33781 14359 33839 14365
rect 33965 14399 34023 14405
rect 33965 14365 33977 14399
rect 34011 14365 34023 14399
rect 33965 14359 34023 14365
rect 29604 14300 30144 14328
rect 30193 14331 30251 14337
rect 29604 14288 29610 14300
rect 30193 14297 30205 14331
rect 30239 14328 30251 14331
rect 30374 14328 30380 14340
rect 30239 14300 30380 14328
rect 30239 14297 30251 14300
rect 30193 14291 30251 14297
rect 30374 14288 30380 14300
rect 30432 14288 30438 14340
rect 33336 14328 33364 14359
rect 33980 14328 34008 14359
rect 34974 14356 34980 14408
rect 35032 14396 35038 14408
rect 35032 14368 35077 14396
rect 35032 14356 35038 14368
rect 34992 14328 35020 14356
rect 33336 14300 35020 14328
rect 37369 14331 37427 14337
rect 37369 14297 37381 14331
rect 37415 14328 37427 14331
rect 38010 14328 38016 14340
rect 37415 14300 38016 14328
rect 37415 14297 37427 14300
rect 37369 14291 37427 14297
rect 38010 14288 38016 14300
rect 38068 14288 38074 14340
rect 9214 14260 9220 14272
rect 9175 14232 9220 14260
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 10134 14260 10140 14272
rect 10095 14232 10140 14260
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 26142 14260 26148 14272
rect 26103 14232 26148 14260
rect 26142 14220 26148 14232
rect 26200 14220 26206 14272
rect 26602 14260 26608 14272
rect 26563 14232 26608 14260
rect 26602 14220 26608 14232
rect 26660 14220 26666 14272
rect 27065 14263 27123 14269
rect 27065 14229 27077 14263
rect 27111 14260 27123 14263
rect 27890 14260 27896 14272
rect 27111 14232 27896 14260
rect 27111 14229 27123 14232
rect 27065 14223 27123 14229
rect 27890 14220 27896 14232
rect 27948 14220 27954 14272
rect 29178 14220 29184 14272
rect 29236 14260 29242 14272
rect 29733 14263 29791 14269
rect 29733 14260 29745 14263
rect 29236 14232 29745 14260
rect 29236 14220 29242 14232
rect 29733 14229 29745 14232
rect 29779 14229 29791 14263
rect 33134 14260 33140 14272
rect 33095 14232 33140 14260
rect 29733 14223 29791 14229
rect 33134 14220 33140 14232
rect 33192 14220 33198 14272
rect 34149 14263 34207 14269
rect 34149 14229 34161 14263
rect 34195 14260 34207 14263
rect 34422 14260 34428 14272
rect 34195 14232 34428 14260
rect 34195 14229 34207 14232
rect 34149 14223 34207 14229
rect 34422 14220 34428 14232
rect 34480 14220 34486 14272
rect 34698 14260 34704 14272
rect 34659 14232 34704 14260
rect 34698 14220 34704 14232
rect 34756 14220 34762 14272
rect 37918 14260 37924 14272
rect 37879 14232 37924 14260
rect 37918 14220 37924 14232
rect 37976 14220 37982 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 15749 14059 15807 14065
rect 15749 14025 15761 14059
rect 15795 14056 15807 14059
rect 16114 14056 16120 14068
rect 15795 14028 16120 14056
rect 15795 14025 15807 14028
rect 15749 14019 15807 14025
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 16853 14059 16911 14065
rect 16853 14025 16865 14059
rect 16899 14056 16911 14059
rect 16942 14056 16948 14068
rect 16899 14028 16948 14056
rect 16899 14025 16911 14028
rect 16853 14019 16911 14025
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 17310 14056 17316 14068
rect 17271 14028 17316 14056
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 19242 14056 19248 14068
rect 19203 14028 19248 14056
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 21177 14059 21235 14065
rect 21177 14025 21189 14059
rect 21223 14056 21235 14059
rect 21818 14056 21824 14068
rect 21223 14028 21824 14056
rect 21223 14025 21235 14028
rect 21177 14019 21235 14025
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 26329 14059 26387 14065
rect 26329 14025 26341 14059
rect 26375 14056 26387 14059
rect 27154 14056 27160 14068
rect 26375 14028 27160 14056
rect 26375 14025 26387 14028
rect 26329 14019 26387 14025
rect 27154 14016 27160 14028
rect 27212 14016 27218 14068
rect 30193 14059 30251 14065
rect 30193 14025 30205 14059
rect 30239 14056 30251 14059
rect 30374 14056 30380 14068
rect 30239 14028 30380 14056
rect 30239 14025 30251 14028
rect 30193 14019 30251 14025
rect 30374 14016 30380 14028
rect 30432 14016 30438 14068
rect 32214 14056 32220 14068
rect 32175 14028 32220 14056
rect 32214 14016 32220 14028
rect 32272 14016 32278 14068
rect 34974 14016 34980 14068
rect 35032 14016 35038 14068
rect 35345 14059 35403 14065
rect 35345 14025 35357 14059
rect 35391 14056 35403 14059
rect 35802 14056 35808 14068
rect 35391 14028 35808 14056
rect 35391 14025 35403 14028
rect 35345 14019 35403 14025
rect 35802 14016 35808 14028
rect 35860 14056 35866 14068
rect 37369 14059 37427 14065
rect 37369 14056 37381 14059
rect 35860 14028 37381 14056
rect 35860 14016 35866 14028
rect 37369 14025 37381 14028
rect 37415 14025 37427 14059
rect 37369 14019 37427 14025
rect 5166 13988 5172 14000
rect 5127 13960 5172 13988
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 10134 13988 10140 14000
rect 7300 13960 10140 13988
rect 5350 13880 5356 13932
rect 5408 13920 5414 13932
rect 7300 13929 7328 13960
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 12986 13988 12992 14000
rect 10244 13960 12992 13988
rect 7285 13923 7343 13929
rect 5408 13892 5453 13920
rect 5408 13880 5414 13892
rect 7285 13889 7297 13923
rect 7331 13889 7343 13923
rect 8662 13920 8668 13932
rect 8623 13892 8668 13920
rect 7285 13883 7343 13889
rect 8662 13880 8668 13892
rect 8720 13880 8726 13932
rect 3970 13852 3976 13864
rect 3931 13824 3976 13852
rect 3970 13812 3976 13824
rect 4028 13812 4034 13864
rect 7006 13852 7012 13864
rect 6967 13824 7012 13852
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 8846 13852 8852 13864
rect 8807 13824 8852 13852
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 9122 13852 9128 13864
rect 9083 13824 9128 13852
rect 9122 13812 9128 13824
rect 9180 13852 9186 13864
rect 10244 13852 10272 13960
rect 12986 13948 12992 13960
rect 13044 13948 13050 14000
rect 28537 13991 28595 13997
rect 28537 13957 28549 13991
rect 28583 13988 28595 13991
rect 29086 13988 29092 14000
rect 28583 13960 29092 13988
rect 28583 13957 28595 13960
rect 28537 13951 28595 13957
rect 10594 13880 10600 13932
rect 10652 13920 10658 13932
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 10652 13892 12081 13920
rect 10652 13880 10658 13892
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13920 16727 13923
rect 17218 13920 17224 13932
rect 16715 13892 17224 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 17494 13920 17500 13932
rect 17455 13892 17500 13920
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 20990 13920 20996 13932
rect 20951 13892 20996 13920
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 29012 13929 29040 13960
rect 29086 13948 29092 13960
rect 29144 13948 29150 14000
rect 34149 13991 34207 13997
rect 34149 13988 34161 13991
rect 30300 13960 34161 13988
rect 28997 13923 29055 13929
rect 28997 13889 29009 13923
rect 29043 13920 29055 13923
rect 29178 13920 29184 13932
rect 29043 13892 29077 13920
rect 29139 13892 29184 13920
rect 29043 13889 29055 13892
rect 28997 13883 29055 13889
rect 29178 13880 29184 13892
rect 29236 13880 29242 13932
rect 30300 13929 30328 13960
rect 30285 13923 30343 13929
rect 30285 13889 30297 13923
rect 30331 13889 30343 13923
rect 31021 13923 31079 13929
rect 31021 13920 31033 13923
rect 30285 13883 30343 13889
rect 30576 13892 31033 13920
rect 9180 13824 10272 13852
rect 12345 13855 12403 13861
rect 9180 13812 9186 13824
rect 12345 13821 12357 13855
rect 12391 13852 12403 13855
rect 12526 13852 12532 13864
rect 12391 13824 12532 13852
rect 12391 13821 12403 13824
rect 12345 13815 12403 13821
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 14642 13852 14648 13864
rect 14603 13824 14648 13852
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 14826 13852 14832 13864
rect 14787 13824 14832 13852
rect 14826 13812 14832 13824
rect 14884 13812 14890 13864
rect 29825 13855 29883 13861
rect 29825 13852 29837 13855
rect 29104 13824 29837 13852
rect 27890 13744 27896 13796
rect 27948 13784 27954 13796
rect 29104 13784 29132 13824
rect 29825 13821 29837 13824
rect 29871 13821 29883 13855
rect 29825 13815 29883 13821
rect 30009 13855 30067 13861
rect 30009 13821 30021 13855
rect 30055 13852 30067 13855
rect 30576 13852 30604 13892
rect 31021 13889 31033 13892
rect 31067 13889 31079 13923
rect 31021 13883 31079 13889
rect 30055 13824 30604 13852
rect 30745 13855 30803 13861
rect 30055 13821 30067 13824
rect 30009 13815 30067 13821
rect 30745 13821 30757 13855
rect 30791 13821 30803 13855
rect 30745 13815 30803 13821
rect 30837 13855 30895 13861
rect 30837 13821 30849 13855
rect 30883 13852 30895 13855
rect 31128 13852 31156 13960
rect 34149 13957 34161 13960
rect 34195 13957 34207 13991
rect 34992 13988 35020 14016
rect 36265 13991 36323 13997
rect 36265 13988 36277 13991
rect 34149 13951 34207 13957
rect 34440 13960 36277 13988
rect 33318 13880 33324 13932
rect 33376 13929 33382 13932
rect 33376 13920 33388 13929
rect 33376 13892 33421 13920
rect 33376 13883 33388 13892
rect 33376 13880 33382 13883
rect 31478 13852 31484 13864
rect 30883 13824 31484 13852
rect 30883 13821 30895 13824
rect 30837 13815 30895 13821
rect 27948 13756 29132 13784
rect 27948 13744 27954 13756
rect 30374 13744 30380 13796
rect 30432 13784 30438 13796
rect 30760 13784 30788 13815
rect 31478 13812 31484 13824
rect 31536 13812 31542 13864
rect 33594 13852 33600 13864
rect 33555 13824 33600 13852
rect 33594 13812 33600 13824
rect 33652 13812 33658 13864
rect 30926 13784 30932 13796
rect 30432 13756 30932 13784
rect 30432 13744 30438 13756
rect 30926 13744 30932 13756
rect 30984 13744 30990 13796
rect 34164 13784 34192 13951
rect 34330 13920 34336 13932
rect 34291 13892 34336 13920
rect 34330 13880 34336 13892
rect 34388 13880 34394 13932
rect 34440 13929 34468 13960
rect 36265 13957 36277 13960
rect 36311 13957 36323 13991
rect 36265 13951 36323 13957
rect 34425 13923 34483 13929
rect 34425 13889 34437 13923
rect 34471 13889 34483 13923
rect 34425 13883 34483 13889
rect 34977 13923 35035 13929
rect 34977 13889 34989 13923
rect 35023 13920 35035 13923
rect 35250 13920 35256 13932
rect 35023 13892 35256 13920
rect 35023 13889 35035 13892
rect 34977 13883 35035 13889
rect 35250 13880 35256 13892
rect 35308 13880 35314 13932
rect 35437 13923 35495 13929
rect 35437 13889 35449 13923
rect 35483 13920 35495 13923
rect 35526 13920 35532 13932
rect 35483 13892 35532 13920
rect 35483 13889 35495 13892
rect 35437 13883 35495 13889
rect 35526 13880 35532 13892
rect 35584 13880 35590 13932
rect 36449 13923 36507 13929
rect 36449 13889 36461 13923
rect 36495 13920 36507 13923
rect 37274 13920 37280 13932
rect 36495 13892 37280 13920
rect 36495 13889 36507 13892
rect 36449 13883 36507 13889
rect 37274 13880 37280 13892
rect 37332 13880 37338 13932
rect 34514 13812 34520 13864
rect 34572 13852 34578 13864
rect 35069 13855 35127 13861
rect 35069 13852 35081 13855
rect 34572 13824 35081 13852
rect 34572 13812 34578 13824
rect 35069 13821 35081 13824
rect 35115 13821 35127 13855
rect 35069 13815 35127 13821
rect 35161 13787 35219 13793
rect 35161 13784 35173 13787
rect 34164 13756 35173 13784
rect 35161 13753 35173 13756
rect 35207 13753 35219 13787
rect 35161 13747 35219 13753
rect 29362 13716 29368 13728
rect 29323 13688 29368 13716
rect 29362 13676 29368 13688
rect 29420 13676 29426 13728
rect 31205 13719 31263 13725
rect 31205 13685 31217 13719
rect 31251 13716 31263 13719
rect 37642 13716 37648 13728
rect 31251 13688 37648 13716
rect 31251 13685 31263 13688
rect 31205 13679 31263 13685
rect 37642 13676 37648 13688
rect 37700 13676 37706 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8904 13484 9045 13512
rect 8904 13472 8910 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 10042 13512 10048 13524
rect 9955 13484 10048 13512
rect 9033 13475 9091 13481
rect 10042 13472 10048 13484
rect 10100 13512 10106 13524
rect 10226 13512 10232 13524
rect 10100 13484 10232 13512
rect 10100 13472 10106 13484
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 10502 13472 10508 13524
rect 10560 13512 10566 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 10560 13484 11621 13512
rect 10560 13472 10566 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 11609 13475 11667 13481
rect 13265 13515 13323 13521
rect 13265 13481 13277 13515
rect 13311 13512 13323 13515
rect 14826 13512 14832 13524
rect 13311 13484 14832 13512
rect 13311 13481 13323 13484
rect 13265 13475 13323 13481
rect 14826 13472 14832 13484
rect 14884 13472 14890 13524
rect 16117 13515 16175 13521
rect 16117 13481 16129 13515
rect 16163 13512 16175 13515
rect 16758 13512 16764 13524
rect 16163 13484 16764 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 16758 13472 16764 13484
rect 16816 13472 16822 13524
rect 17218 13512 17224 13524
rect 17179 13484 17224 13512
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19705 13515 19763 13521
rect 19705 13512 19717 13515
rect 19392 13484 19717 13512
rect 19392 13472 19398 13484
rect 19705 13481 19717 13484
rect 19751 13481 19763 13515
rect 19705 13475 19763 13481
rect 20165 13515 20223 13521
rect 20165 13481 20177 13515
rect 20211 13512 20223 13515
rect 20990 13512 20996 13524
rect 20211 13484 20996 13512
rect 20211 13481 20223 13484
rect 20165 13475 20223 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 27614 13512 27620 13524
rect 26528 13484 27620 13512
rect 7006 13404 7012 13456
rect 7064 13404 7070 13456
rect 8202 13404 8208 13456
rect 8260 13444 8266 13456
rect 10873 13447 10931 13453
rect 10873 13444 10885 13447
rect 8260 13416 10885 13444
rect 8260 13404 8266 13416
rect 10873 13413 10885 13416
rect 10919 13413 10931 13447
rect 10873 13407 10931 13413
rect 15289 13447 15347 13453
rect 15289 13413 15301 13447
rect 15335 13413 15347 13447
rect 15289 13407 15347 13413
rect 16301 13447 16359 13453
rect 16301 13413 16313 13447
rect 16347 13444 16359 13447
rect 17494 13444 17500 13456
rect 16347 13416 17500 13444
rect 16347 13413 16359 13416
rect 16301 13407 16359 13413
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 5169 13379 5227 13385
rect 5169 13376 5181 13379
rect 4212 13348 5181 13376
rect 4212 13336 4218 13348
rect 5169 13345 5181 13348
rect 5215 13376 5227 13379
rect 5534 13376 5540 13388
rect 5215 13348 5540 13376
rect 5215 13345 5227 13348
rect 5169 13339 5227 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 6825 13379 6883 13385
rect 6825 13345 6837 13379
rect 6871 13376 6883 13379
rect 7024 13376 7052 13404
rect 6871 13348 7052 13376
rect 6871 13345 6883 13348
rect 6825 13339 6883 13345
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13308 1458 13320
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 1452 13280 2053 13308
rect 1452 13268 1458 13280
rect 2041 13277 2053 13280
rect 2087 13277 2099 13311
rect 2041 13271 2099 13277
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 8386 13308 8392 13320
rect 7064 13280 7109 13308
rect 8347 13280 8392 13308
rect 7064 13268 7070 13280
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 9214 13308 9220 13320
rect 9175 13280 9220 13308
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13308 10287 13311
rect 10502 13308 10508 13320
rect 10275 13280 10508 13308
rect 10275 13277 10287 13280
rect 10229 13271 10287 13277
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 10888 13308 10916 13407
rect 15304 13376 15332 13407
rect 17494 13404 17500 13416
rect 17552 13404 17558 13456
rect 16022 13376 16028 13388
rect 15304 13348 16028 13376
rect 16022 13336 16028 13348
rect 16080 13376 16086 13388
rect 16853 13379 16911 13385
rect 16853 13376 16865 13379
rect 16080 13348 16865 13376
rect 16080 13336 16086 13348
rect 16853 13345 16865 13348
rect 16899 13376 16911 13379
rect 17681 13379 17739 13385
rect 17681 13376 17693 13379
rect 16899 13348 17693 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 17681 13345 17693 13348
rect 17727 13345 17739 13379
rect 17681 13339 17739 13345
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 19484 13348 19901 13376
rect 19484 13336 19490 13348
rect 19889 13345 19901 13348
rect 19935 13376 19947 13379
rect 20530 13376 20536 13388
rect 19935 13348 20536 13376
rect 19935 13345 19947 13348
rect 19889 13339 19947 13345
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 26528 13385 26556 13484
rect 27614 13472 27620 13484
rect 27672 13512 27678 13524
rect 28353 13515 28411 13521
rect 28353 13512 28365 13515
rect 27672 13484 28365 13512
rect 27672 13472 27678 13484
rect 28353 13481 28365 13484
rect 28399 13481 28411 13515
rect 30926 13512 30932 13524
rect 30887 13484 30932 13512
rect 28353 13475 28411 13481
rect 30926 13472 30932 13484
rect 30984 13472 30990 13524
rect 33318 13472 33324 13524
rect 33376 13512 33382 13524
rect 33413 13515 33471 13521
rect 33413 13512 33425 13515
rect 33376 13484 33425 13512
rect 33376 13472 33382 13484
rect 33413 13481 33425 13484
rect 33459 13481 33471 13515
rect 36446 13512 36452 13524
rect 36407 13484 36452 13512
rect 33413 13475 33471 13481
rect 36446 13472 36452 13484
rect 36504 13472 36510 13524
rect 27890 13444 27896 13456
rect 27851 13416 27896 13444
rect 27890 13404 27896 13416
rect 27948 13404 27954 13456
rect 26513 13379 26571 13385
rect 26513 13345 26525 13379
rect 26559 13345 26571 13379
rect 32125 13379 32183 13385
rect 32125 13376 32137 13379
rect 26513 13339 26571 13345
rect 31726 13348 32137 13376
rect 11425 13311 11483 13317
rect 11425 13308 11437 13311
rect 10888 13280 11437 13308
rect 11425 13277 11437 13280
rect 11471 13277 11483 13311
rect 12526 13308 12532 13320
rect 12439 13280 12532 13308
rect 11425 13271 11483 13277
rect 11440 13240 11468 13271
rect 12526 13268 12532 13280
rect 12584 13308 12590 13320
rect 15105 13311 15163 13317
rect 15105 13308 15117 13311
rect 12584 13280 15117 13308
rect 12584 13268 12590 13280
rect 15105 13277 15117 13280
rect 15151 13308 15163 13311
rect 15194 13308 15200 13320
rect 15151 13280 15200 13308
rect 15151 13277 15163 13280
rect 15105 13271 15163 13277
rect 15194 13268 15200 13280
rect 15252 13268 15258 13320
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13308 16175 13311
rect 17037 13311 17095 13317
rect 17037 13308 17049 13311
rect 16163 13280 17049 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 17037 13277 17049 13280
rect 17083 13308 17095 13311
rect 18230 13308 18236 13320
rect 17083 13280 18236 13308
rect 17083 13277 17095 13280
rect 17037 13271 17095 13277
rect 18230 13268 18236 13280
rect 18288 13308 18294 13320
rect 19978 13308 19984 13320
rect 18288 13280 19984 13308
rect 18288 13268 18294 13280
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 22278 13268 22284 13320
rect 22336 13308 22342 13320
rect 22373 13311 22431 13317
rect 22373 13308 22385 13311
rect 22336 13280 22385 13308
rect 22336 13268 22342 13280
rect 22373 13277 22385 13280
rect 22419 13277 22431 13311
rect 22373 13271 22431 13277
rect 26053 13311 26111 13317
rect 26053 13277 26065 13311
rect 26099 13308 26111 13311
rect 26602 13308 26608 13320
rect 26099 13280 26608 13308
rect 26099 13277 26111 13280
rect 26053 13271 26111 13277
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 29549 13311 29607 13317
rect 29549 13308 29561 13311
rect 29012 13280 29561 13308
rect 11440 13212 12848 13240
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 12820 13172 12848 13212
rect 12894 13200 12900 13252
rect 12952 13240 12958 13252
rect 15841 13243 15899 13249
rect 15841 13240 15853 13243
rect 12952 13212 15853 13240
rect 12952 13200 12958 13212
rect 15841 13209 15853 13212
rect 15887 13240 15899 13243
rect 16761 13243 16819 13249
rect 16761 13240 16773 13243
rect 15887 13212 16773 13240
rect 15887 13209 15899 13212
rect 15841 13203 15899 13209
rect 16761 13209 16773 13212
rect 16807 13209 16819 13243
rect 16761 13203 16819 13209
rect 19705 13243 19763 13249
rect 19705 13209 19717 13243
rect 19751 13240 19763 13243
rect 20438 13240 20444 13252
rect 19751 13212 20444 13240
rect 19751 13209 19763 13212
rect 19705 13203 19763 13209
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 25866 13240 25872 13252
rect 25827 13212 25872 13240
rect 25866 13200 25872 13212
rect 25924 13200 25930 13252
rect 26780 13243 26838 13249
rect 26780 13209 26792 13243
rect 26826 13240 26838 13243
rect 26970 13240 26976 13252
rect 26826 13212 26976 13240
rect 26826 13209 26838 13212
rect 26780 13203 26838 13209
rect 26970 13200 26976 13212
rect 27028 13200 27034 13252
rect 29012 13184 29040 13280
rect 29549 13277 29561 13280
rect 29595 13308 29607 13311
rect 31726 13308 31754 13348
rect 32125 13345 32137 13348
rect 32171 13376 32183 13379
rect 32171 13348 33640 13376
rect 32171 13345 32183 13348
rect 32125 13339 32183 13345
rect 33612 13320 33640 13348
rect 33134 13308 33140 13320
rect 29595 13280 31754 13308
rect 33095 13280 33140 13308
rect 29595 13277 29607 13280
rect 29549 13271 29607 13277
rect 33134 13268 33140 13280
rect 33192 13268 33198 13320
rect 33594 13268 33600 13320
rect 33652 13308 33658 13320
rect 35069 13311 35127 13317
rect 35069 13308 35081 13311
rect 33652 13280 35081 13308
rect 33652 13268 33658 13280
rect 35069 13277 35081 13280
rect 35115 13308 35127 13311
rect 35115 13280 35480 13308
rect 35115 13277 35127 13280
rect 35069 13271 35127 13277
rect 35452 13252 35480 13280
rect 29822 13249 29828 13252
rect 29816 13203 29828 13249
rect 29880 13240 29886 13252
rect 29880 13212 29916 13240
rect 29822 13200 29828 13203
rect 29880 13200 29886 13212
rect 31662 13200 31668 13252
rect 31720 13240 31726 13252
rect 33413 13243 33471 13249
rect 33413 13240 33425 13243
rect 31720 13212 33425 13240
rect 31720 13200 31726 13212
rect 33413 13209 33425 13212
rect 33459 13240 33471 13243
rect 34514 13240 34520 13252
rect 33459 13212 34520 13240
rect 33459 13209 33471 13212
rect 33413 13203 33471 13209
rect 34514 13200 34520 13212
rect 34572 13200 34578 13252
rect 34790 13200 34796 13252
rect 34848 13240 34854 13252
rect 35314 13243 35372 13249
rect 35314 13240 35326 13243
rect 34848 13212 35326 13240
rect 34848 13200 34854 13212
rect 35314 13209 35326 13212
rect 35360 13209 35372 13243
rect 35314 13203 35372 13209
rect 35434 13200 35440 13252
rect 35492 13200 35498 13252
rect 16850 13172 16856 13184
rect 12820 13144 16856 13172
rect 16850 13132 16856 13144
rect 16908 13132 16914 13184
rect 25685 13175 25743 13181
rect 25685 13141 25697 13175
rect 25731 13172 25743 13175
rect 27154 13172 27160 13184
rect 25731 13144 27160 13172
rect 25731 13141 25743 13144
rect 25685 13135 25743 13141
rect 27154 13132 27160 13144
rect 27212 13132 27218 13184
rect 28994 13172 29000 13184
rect 28955 13144 29000 13172
rect 28994 13132 29000 13144
rect 29052 13132 29058 13184
rect 33229 13175 33287 13181
rect 33229 13141 33241 13175
rect 33275 13172 33287 13175
rect 34422 13172 34428 13184
rect 33275 13144 34428 13172
rect 33275 13141 33287 13144
rect 33229 13135 33287 13141
rect 34422 13132 34428 13144
rect 34480 13132 34486 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10689 12971 10747 12977
rect 10689 12968 10701 12971
rect 10560 12940 10701 12968
rect 10560 12928 10566 12940
rect 10689 12937 10701 12940
rect 10735 12968 10747 12971
rect 11422 12968 11428 12980
rect 10735 12940 11428 12968
rect 10735 12937 10747 12940
rect 10689 12931 10747 12937
rect 11422 12928 11428 12940
rect 11480 12968 11486 12980
rect 12069 12971 12127 12977
rect 12069 12968 12081 12971
rect 11480 12940 12081 12968
rect 11480 12928 11486 12940
rect 12069 12937 12081 12940
rect 12115 12937 12127 12971
rect 12069 12931 12127 12937
rect 2498 12900 2504 12912
rect 2459 12872 2504 12900
rect 2498 12860 2504 12872
rect 2556 12860 2562 12912
rect 2774 12792 2780 12844
rect 2832 12832 2838 12844
rect 5445 12835 5503 12841
rect 2832 12804 2877 12832
rect 2832 12792 2838 12804
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 7006 12832 7012 12844
rect 5491 12804 7012 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 8386 12832 8392 12844
rect 8347 12804 8392 12832
rect 8386 12792 8392 12804
rect 8444 12792 8450 12844
rect 12084 12832 12112 12931
rect 15194 12928 15200 12980
rect 15252 12968 15258 12980
rect 15473 12971 15531 12977
rect 15473 12968 15485 12971
rect 15252 12940 15485 12968
rect 15252 12928 15258 12940
rect 15473 12937 15485 12940
rect 15519 12937 15531 12971
rect 17034 12968 17040 12980
rect 16995 12940 17040 12968
rect 15473 12931 15531 12937
rect 17034 12928 17040 12940
rect 17092 12928 17098 12980
rect 19334 12968 19340 12980
rect 18248 12940 19340 12968
rect 16758 12860 16764 12912
rect 16816 12900 16822 12912
rect 18248 12900 18276 12940
rect 19334 12928 19340 12940
rect 19392 12928 19398 12980
rect 20073 12971 20131 12977
rect 20073 12937 20085 12971
rect 20119 12968 20131 12971
rect 20162 12968 20168 12980
rect 20119 12940 20168 12968
rect 20119 12937 20131 12940
rect 20073 12931 20131 12937
rect 16816 12872 18276 12900
rect 16816 12860 16822 12872
rect 12621 12835 12679 12841
rect 12621 12832 12633 12835
rect 12084 12804 12633 12832
rect 12621 12801 12633 12804
rect 12667 12801 12679 12835
rect 12894 12832 12900 12844
rect 12855 12804 12900 12832
rect 12621 12795 12679 12801
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 14642 12832 14648 12844
rect 14603 12804 14648 12832
rect 14642 12792 14648 12804
rect 14700 12792 14706 12844
rect 17126 12832 17132 12844
rect 17087 12804 17132 12832
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 18248 12841 18276 12872
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12832 19395 12835
rect 19426 12832 19432 12844
rect 19383 12804 19432 12832
rect 19383 12801 19395 12804
rect 19337 12795 19395 12801
rect 19426 12792 19432 12804
rect 19484 12832 19490 12844
rect 20088 12832 20116 12931
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 26970 12968 26976 12980
rect 26931 12940 26976 12968
rect 26970 12928 26976 12940
rect 27028 12928 27034 12980
rect 29822 12968 29828 12980
rect 29783 12940 29828 12968
rect 29822 12928 29828 12940
rect 29880 12928 29886 12980
rect 34517 12971 34575 12977
rect 34517 12937 34529 12971
rect 34563 12968 34575 12971
rect 34698 12968 34704 12980
rect 34563 12940 34704 12968
rect 34563 12937 34575 12940
rect 34517 12931 34575 12937
rect 34698 12928 34704 12940
rect 34756 12928 34762 12980
rect 20346 12832 20352 12844
rect 19484 12804 20352 12832
rect 19484 12792 19490 12804
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 22278 12832 22284 12844
rect 22239 12804 22284 12832
rect 22278 12792 22284 12804
rect 22336 12792 22342 12844
rect 27154 12832 27160 12844
rect 27115 12804 27160 12832
rect 27154 12792 27160 12804
rect 27212 12792 27218 12844
rect 29362 12792 29368 12844
rect 29420 12832 29426 12844
rect 30009 12835 30067 12841
rect 30009 12832 30021 12835
rect 29420 12804 30021 12832
rect 29420 12792 29426 12804
rect 30009 12801 30021 12804
rect 30055 12801 30067 12835
rect 34422 12832 34428 12844
rect 34383 12804 34428 12832
rect 30009 12795 30067 12801
rect 34422 12792 34428 12804
rect 34480 12792 34486 12844
rect 34698 12832 34704 12844
rect 34659 12804 34704 12832
rect 34698 12792 34704 12804
rect 34756 12792 34762 12844
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 8570 12764 8576 12776
rect 8531 12736 8576 12764
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 9766 12764 9772 12776
rect 9727 12736 9772 12764
rect 9766 12724 9772 12736
rect 9824 12724 9830 12776
rect 14921 12767 14979 12773
rect 14921 12733 14933 12767
rect 14967 12764 14979 12767
rect 17862 12764 17868 12776
rect 14967 12736 17868 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12764 18567 12767
rect 18598 12764 18604 12776
rect 18555 12736 18604 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 22462 12764 22468 12776
rect 22423 12736 22468 12764
rect 22462 12724 22468 12736
rect 22520 12724 22526 12776
rect 23474 12764 23480 12776
rect 23435 12736 23480 12764
rect 23474 12724 23480 12736
rect 23532 12724 23538 12776
rect 19521 12699 19579 12705
rect 19521 12665 19533 12699
rect 19567 12696 19579 12699
rect 20438 12696 20444 12708
rect 19567 12668 20444 12696
rect 19567 12665 19579 12668
rect 19521 12659 19579 12665
rect 20438 12656 20444 12668
rect 20496 12656 20502 12708
rect 34701 12699 34759 12705
rect 34701 12665 34713 12699
rect 34747 12696 34759 12699
rect 34790 12696 34796 12708
rect 34747 12668 34796 12696
rect 34747 12665 34759 12668
rect 34701 12659 34759 12665
rect 34790 12656 34796 12668
rect 34848 12656 34854 12708
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 2406 12628 2412 12640
rect 1636 12600 2412 12628
rect 1636 12588 1642 12600
rect 2406 12588 2412 12600
rect 2464 12628 2470 12640
rect 2501 12631 2559 12637
rect 2501 12628 2513 12631
rect 2464 12600 2513 12628
rect 2464 12588 2470 12600
rect 2501 12597 2513 12600
rect 2547 12597 2559 12631
rect 2501 12591 2559 12597
rect 2961 12631 3019 12637
rect 2961 12597 2973 12631
rect 3007 12628 3019 12631
rect 3970 12628 3976 12640
rect 3007 12600 3976 12628
rect 3007 12597 3019 12600
rect 2961 12591 3019 12597
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 4798 12628 4804 12640
rect 4759 12600 4804 12628
rect 4798 12588 4804 12600
rect 4856 12588 4862 12640
rect 35253 12631 35311 12637
rect 35253 12597 35265 12631
rect 35299 12628 35311 12631
rect 35434 12628 35440 12640
rect 35299 12600 35440 12628
rect 35299 12597 35311 12600
rect 35253 12591 35311 12597
rect 35434 12588 35440 12600
rect 35492 12588 35498 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 2590 12424 2596 12436
rect 2551 12396 2596 12424
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 10410 12384 10416 12436
rect 10468 12424 10474 12436
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 10468 12396 10701 12424
rect 10468 12384 10474 12396
rect 10689 12393 10701 12396
rect 10735 12393 10747 12427
rect 10689 12387 10747 12393
rect 14185 12427 14243 12433
rect 14185 12393 14197 12427
rect 14231 12424 14243 12427
rect 15102 12424 15108 12436
rect 14231 12396 15108 12424
rect 14231 12393 14243 12396
rect 14185 12387 14243 12393
rect 10505 12359 10563 12365
rect 10505 12356 10517 12359
rect 10060 12328 10517 12356
rect 2406 12248 2412 12300
rect 2464 12288 2470 12300
rect 2593 12291 2651 12297
rect 2593 12288 2605 12291
rect 2464 12260 2605 12288
rect 2464 12248 2470 12260
rect 2593 12257 2605 12260
rect 2639 12257 2651 12291
rect 2593 12251 2651 12257
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 5261 12291 5319 12297
rect 5261 12288 5273 12291
rect 4856 12260 5273 12288
rect 4856 12248 4862 12260
rect 5261 12257 5273 12260
rect 5307 12257 5319 12291
rect 5261 12251 5319 12257
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 5592 12260 5733 12288
rect 5592 12248 5598 12260
rect 5721 12257 5733 12260
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 10060 12297 10088 12328
rect 10505 12325 10517 12328
rect 10551 12325 10563 12359
rect 10505 12319 10563 12325
rect 9769 12291 9827 12297
rect 9769 12288 9781 12291
rect 8628 12260 9781 12288
rect 8628 12248 8634 12260
rect 9769 12257 9781 12260
rect 9815 12257 9827 12291
rect 9769 12251 9827 12257
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 10594 12248 10600 12300
rect 10652 12288 10658 12300
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 10652 12260 10793 12288
rect 10652 12248 10658 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 2498 12220 2504 12232
rect 2459 12192 2504 12220
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 10686 12220 10692 12232
rect 10647 12192 10692 12220
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 11422 12220 11428 12232
rect 11383 12192 11428 12220
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12216 12403 12223
rect 14200 12220 14228 12387
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 20165 12427 20223 12433
rect 20165 12393 20177 12427
rect 20211 12424 20223 12427
rect 20346 12424 20352 12436
rect 20211 12396 20352 12424
rect 20211 12393 20223 12396
rect 20165 12387 20223 12393
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 22462 12384 22468 12436
rect 22520 12424 22526 12436
rect 22833 12427 22891 12433
rect 22833 12424 22845 12427
rect 22520 12396 22845 12424
rect 22520 12384 22526 12396
rect 22833 12393 22845 12396
rect 22879 12393 22891 12427
rect 35434 12424 35440 12436
rect 35395 12396 35440 12424
rect 22833 12387 22891 12393
rect 35434 12384 35440 12396
rect 35492 12384 35498 12436
rect 37274 12384 37280 12436
rect 37332 12424 37338 12436
rect 37369 12427 37427 12433
rect 37369 12424 37381 12427
rect 37332 12396 37381 12424
rect 37332 12384 37338 12396
rect 37369 12393 37381 12396
rect 37415 12393 37427 12427
rect 37369 12387 37427 12393
rect 18230 12288 18236 12300
rect 18191 12260 18236 12288
rect 18230 12248 18236 12260
rect 18288 12248 18294 12300
rect 26142 12248 26148 12300
rect 26200 12288 26206 12300
rect 26513 12291 26571 12297
rect 26513 12288 26525 12291
rect 26200 12260 26525 12288
rect 26200 12248 26206 12260
rect 26513 12257 26525 12260
rect 26559 12257 26571 12291
rect 35452 12288 35480 12384
rect 35989 12291 36047 12297
rect 35989 12288 36001 12291
rect 35452 12260 36001 12288
rect 26513 12251 26571 12257
rect 35989 12257 36001 12260
rect 36035 12257 36047 12291
rect 35989 12251 36047 12257
rect 18506 12220 18512 12232
rect 12452 12216 14228 12220
rect 12391 12192 14228 12216
rect 18467 12192 18512 12220
rect 12391 12189 12480 12192
rect 12345 12188 12480 12189
rect 12345 12183 12403 12188
rect 18506 12180 18512 12192
rect 18564 12180 18570 12232
rect 19426 12220 19432 12232
rect 19387 12192 19432 12220
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 20898 12180 20904 12232
rect 20956 12220 20962 12232
rect 22281 12223 22339 12229
rect 22281 12220 22293 12223
rect 20956 12192 22293 12220
rect 20956 12180 20962 12192
rect 22281 12189 22293 12192
rect 22327 12189 22339 12223
rect 23014 12220 23020 12232
rect 22975 12192 23020 12220
rect 22281 12183 22339 12189
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 35342 12180 35348 12232
rect 35400 12220 35406 12232
rect 36245 12223 36303 12229
rect 36245 12220 36257 12223
rect 35400 12192 36257 12220
rect 35400 12180 35406 12192
rect 36245 12189 36257 12192
rect 36291 12189 36303 12223
rect 36245 12183 36303 12189
rect 5445 12155 5503 12161
rect 5445 12121 5457 12155
rect 5491 12152 5503 12155
rect 6362 12152 6368 12164
rect 5491 12124 6368 12152
rect 5491 12121 5503 12124
rect 5445 12115 5503 12121
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 10042 12112 10048 12164
rect 10100 12152 10106 12164
rect 10965 12155 11023 12161
rect 10965 12152 10977 12155
rect 10100 12124 10977 12152
rect 10100 12112 10106 12124
rect 10965 12121 10977 12124
rect 11011 12121 11023 12155
rect 10965 12115 11023 12121
rect 14642 12112 14648 12164
rect 14700 12152 14706 12164
rect 21910 12152 21916 12164
rect 14700 12124 21916 12152
rect 14700 12112 14706 12124
rect 21910 12112 21916 12124
rect 21968 12112 21974 12164
rect 22094 12152 22100 12164
rect 22055 12124 22100 12152
rect 22094 12112 22100 12124
rect 22152 12112 22158 12164
rect 25498 12112 25504 12164
rect 25556 12152 25562 12164
rect 25685 12155 25743 12161
rect 25685 12152 25697 12155
rect 25556 12124 25697 12152
rect 25556 12112 25562 12124
rect 25685 12121 25697 12124
rect 25731 12121 25743 12155
rect 25866 12152 25872 12164
rect 25827 12124 25872 12152
rect 25685 12115 25743 12121
rect 25866 12112 25872 12124
rect 25924 12152 25930 12164
rect 30374 12152 30380 12164
rect 25924 12124 30380 12152
rect 25924 12112 25930 12124
rect 30374 12112 30380 12124
rect 30432 12112 30438 12164
rect 1578 12084 1584 12096
rect 1539 12056 1584 12084
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 2869 12087 2927 12093
rect 2869 12053 2881 12087
rect 2915 12084 2927 12087
rect 2958 12084 2964 12096
rect 2915 12056 2964 12084
rect 2915 12053 2927 12056
rect 2869 12047 2927 12053
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 10686 12044 10692 12096
rect 10744 12084 10750 12096
rect 11609 12087 11667 12093
rect 11609 12084 11621 12087
rect 10744 12056 11621 12084
rect 10744 12044 10750 12056
rect 11609 12053 11621 12056
rect 11655 12053 11667 12087
rect 12526 12084 12532 12096
rect 12487 12056 12532 12084
rect 11609 12047 11667 12053
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 13354 12084 13360 12096
rect 13315 12056 13360 12084
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 19613 12087 19671 12093
rect 19613 12053 19625 12087
rect 19659 12084 19671 12087
rect 20254 12084 20260 12096
rect 19659 12056 20260 12084
rect 19659 12053 19671 12056
rect 19613 12047 19671 12053
rect 20254 12044 20260 12056
rect 20312 12044 20318 12096
rect 26053 12087 26111 12093
rect 26053 12053 26065 12087
rect 26099 12084 26111 12087
rect 26970 12084 26976 12096
rect 26099 12056 26976 12084
rect 26099 12053 26111 12056
rect 26053 12047 26111 12053
rect 26970 12044 26976 12056
rect 27028 12044 27034 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 6362 11880 6368 11892
rect 6323 11852 6368 11880
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 11422 11840 11428 11892
rect 11480 11880 11486 11892
rect 11701 11883 11759 11889
rect 11701 11880 11713 11883
rect 11480 11852 11713 11880
rect 11480 11840 11486 11852
rect 11701 11849 11713 11852
rect 11747 11849 11759 11883
rect 11701 11843 11759 11849
rect 17862 11840 17868 11892
rect 17920 11880 17926 11892
rect 19889 11883 19947 11889
rect 19889 11880 19901 11883
rect 17920 11852 19901 11880
rect 17920 11840 17926 11852
rect 19889 11849 19901 11852
rect 19935 11849 19947 11883
rect 20622 11880 20628 11892
rect 19889 11843 19947 11849
rect 20088 11852 20628 11880
rect 1394 11812 1400 11824
rect 1355 11784 1400 11812
rect 1394 11772 1400 11784
rect 1452 11772 1458 11824
rect 13998 11812 14004 11824
rect 13096 11784 14004 11812
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11744 10563 11747
rect 10686 11744 10692 11756
rect 10551 11716 10692 11744
rect 10551 11713 10563 11716
rect 10505 11707 10563 11713
rect 6564 11608 6592 11707
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 13096 11753 13124 11784
rect 13998 11772 14004 11784
rect 14056 11772 14062 11824
rect 18506 11772 18512 11824
rect 18564 11812 18570 11824
rect 18564 11784 19288 11812
rect 18564 11772 18570 11784
rect 13081 11747 13139 11753
rect 10836 11716 10881 11744
rect 10836 11704 10842 11716
rect 13081 11713 13093 11747
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 13354 11704 13360 11756
rect 13412 11744 13418 11756
rect 13633 11747 13691 11753
rect 13633 11744 13645 11747
rect 13412 11716 13645 11744
rect 13412 11704 13418 11716
rect 13633 11713 13645 11716
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 16908 11716 16957 11744
rect 16908 11704 16914 11716
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 18598 11744 18604 11756
rect 18559 11716 18604 11744
rect 16945 11707 17003 11713
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 19260 11753 19288 11784
rect 19245 11747 19303 11753
rect 19245 11713 19257 11747
rect 19291 11713 19303 11747
rect 19245 11707 19303 11713
rect 19426 11704 19432 11756
rect 19484 11744 19490 11756
rect 20088 11753 20116 11852
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 22281 11883 22339 11889
rect 22281 11849 22293 11883
rect 22327 11880 22339 11883
rect 23014 11880 23020 11892
rect 22327 11852 23020 11880
rect 22327 11849 22339 11852
rect 22281 11843 22339 11849
rect 23014 11840 23020 11852
rect 23072 11840 23078 11892
rect 25498 11880 25504 11892
rect 25459 11852 25504 11880
rect 25498 11840 25504 11852
rect 25556 11840 25562 11892
rect 29825 11883 29883 11889
rect 29825 11849 29837 11883
rect 29871 11849 29883 11883
rect 29825 11843 29883 11849
rect 30561 11883 30619 11889
rect 30561 11849 30573 11883
rect 30607 11880 30619 11883
rect 31110 11880 31116 11892
rect 30607 11852 31116 11880
rect 30607 11849 30619 11852
rect 30561 11843 30619 11849
rect 20254 11772 20260 11824
rect 20312 11812 20318 11824
rect 20349 11815 20407 11821
rect 20349 11812 20361 11815
rect 20312 11784 20361 11812
rect 20312 11772 20318 11784
rect 20349 11781 20361 11784
rect 20395 11812 20407 11815
rect 21821 11815 21879 11821
rect 21821 11812 21833 11815
rect 20395 11784 21833 11812
rect 20395 11781 20407 11784
rect 20349 11775 20407 11781
rect 21821 11781 21833 11784
rect 21867 11781 21879 11815
rect 21821 11775 21879 11781
rect 21910 11772 21916 11824
rect 21968 11812 21974 11824
rect 29086 11812 29092 11824
rect 21968 11784 29092 11812
rect 21968 11772 21974 11784
rect 29086 11772 29092 11784
rect 29144 11812 29150 11824
rect 29840 11812 29868 11843
rect 29144 11784 29868 11812
rect 29144 11772 29150 11784
rect 20073 11747 20131 11753
rect 20073 11744 20085 11747
rect 19484 11716 20085 11744
rect 19484 11704 19490 11716
rect 20073 11713 20085 11716
rect 20119 11713 20131 11747
rect 22002 11744 22008 11756
rect 20073 11707 20131 11713
rect 20180 11716 22008 11744
rect 10594 11676 10600 11688
rect 10555 11648 10600 11676
rect 10594 11636 10600 11648
rect 10652 11636 10658 11688
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 11940 11648 12817 11676
rect 11940 11636 11946 11648
rect 12805 11645 12817 11648
rect 12851 11645 12863 11679
rect 13814 11676 13820 11688
rect 13775 11648 13820 11676
rect 12805 11639 12863 11645
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 16666 11636 16672 11688
rect 16724 11676 16730 11688
rect 17126 11676 17132 11688
rect 16724 11648 17132 11676
rect 16724 11636 16730 11648
rect 17126 11636 17132 11648
rect 17184 11676 17190 11688
rect 20180 11685 20208 11716
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 17221 11679 17279 11685
rect 17221 11676 17233 11679
rect 17184 11648 17233 11676
rect 17184 11636 17190 11648
rect 17221 11645 17233 11648
rect 17267 11676 17279 11679
rect 20165 11679 20223 11685
rect 20165 11676 20177 11679
rect 17267 11648 20177 11676
rect 17267 11645 17279 11648
rect 17221 11639 17279 11645
rect 20165 11645 20177 11648
rect 20211 11645 20223 11679
rect 20165 11639 20223 11645
rect 15378 11608 15384 11620
rect 6564 11580 15384 11608
rect 15378 11568 15384 11580
rect 15436 11568 15442 11620
rect 18785 11611 18843 11617
rect 18785 11577 18797 11611
rect 18831 11608 18843 11611
rect 18831 11580 20116 11608
rect 18831 11577 18843 11580
rect 18785 11571 18843 11577
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 10594 11540 10600 11552
rect 10468 11512 10600 11540
rect 10468 11500 10474 11512
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 10962 11540 10968 11552
rect 10923 11512 10968 11540
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 15930 11540 15936 11552
rect 15891 11512 15936 11540
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 19426 11540 19432 11552
rect 19387 11512 19432 11540
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 20088 11549 20116 11580
rect 20622 11568 20628 11620
rect 20680 11608 20686 11620
rect 22112 11608 22140 11707
rect 25222 11704 25228 11756
rect 25280 11744 25286 11756
rect 25869 11747 25927 11753
rect 25869 11744 25881 11747
rect 25280 11716 25881 11744
rect 25280 11704 25286 11716
rect 25869 11713 25881 11716
rect 25915 11744 25927 11747
rect 26142 11744 26148 11756
rect 25915 11716 26148 11744
rect 25915 11713 25927 11716
rect 25869 11707 25927 11713
rect 26142 11704 26148 11716
rect 26200 11704 26206 11756
rect 26970 11744 26976 11756
rect 26931 11716 26976 11744
rect 26970 11704 26976 11716
rect 27028 11704 27034 11756
rect 30009 11747 30067 11753
rect 30009 11713 30021 11747
rect 30055 11744 30067 11747
rect 30466 11744 30472 11756
rect 30055 11716 30472 11744
rect 30055 11713 30067 11716
rect 30009 11707 30067 11713
rect 30466 11704 30472 11716
rect 30524 11744 30530 11756
rect 30576 11744 30604 11843
rect 31110 11840 31116 11852
rect 31168 11840 31174 11892
rect 30524 11716 30604 11744
rect 30524 11704 30530 11716
rect 25958 11676 25964 11688
rect 25919 11648 25964 11676
rect 25958 11636 25964 11648
rect 26016 11636 26022 11688
rect 26053 11679 26111 11685
rect 26053 11645 26065 11679
rect 26099 11645 26111 11679
rect 26053 11639 26111 11645
rect 20680 11580 22140 11608
rect 20680 11568 20686 11580
rect 25406 11568 25412 11620
rect 25464 11608 25470 11620
rect 26068 11608 26096 11639
rect 25464 11580 26096 11608
rect 25464 11568 25470 11580
rect 20073 11543 20131 11549
rect 20073 11509 20085 11543
rect 20119 11540 20131 11543
rect 20346 11540 20352 11552
rect 20119 11512 20352 11540
rect 20119 11509 20131 11512
rect 20073 11503 20131 11509
rect 20346 11500 20352 11512
rect 20404 11540 20410 11552
rect 21821 11543 21879 11549
rect 21821 11540 21833 11543
rect 20404 11512 21833 11540
rect 20404 11500 20410 11512
rect 21821 11509 21833 11512
rect 21867 11509 21879 11543
rect 27154 11540 27160 11552
rect 27115 11512 27160 11540
rect 21821 11503 21879 11509
rect 27154 11500 27160 11512
rect 27212 11500 27218 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1578 11296 1584 11348
rect 1636 11336 1642 11348
rect 2501 11339 2559 11345
rect 2501 11336 2513 11339
rect 1636 11308 2513 11336
rect 1636 11296 1642 11308
rect 2501 11305 2513 11308
rect 2547 11336 2559 11339
rect 2590 11336 2596 11348
rect 2547 11308 2596 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 10652 11308 10977 11336
rect 10652 11296 10658 11308
rect 10965 11305 10977 11308
rect 11011 11336 11023 11339
rect 11882 11336 11888 11348
rect 11011 11308 11888 11336
rect 11011 11305 11023 11308
rect 10965 11299 11023 11305
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 15378 11336 15384 11348
rect 15339 11308 15384 11336
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15565 11339 15623 11345
rect 15565 11305 15577 11339
rect 15611 11305 15623 11339
rect 16666 11336 16672 11348
rect 15565 11299 15623 11305
rect 15764 11308 16672 11336
rect 10781 11271 10839 11277
rect 10781 11237 10793 11271
rect 10827 11268 10839 11271
rect 10870 11268 10876 11280
rect 10827 11240 10876 11268
rect 10827 11237 10839 11240
rect 10781 11231 10839 11237
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 15102 11228 15108 11280
rect 15160 11268 15166 11280
rect 15580 11268 15608 11299
rect 15160 11240 15608 11268
rect 15160 11228 15166 11240
rect 2498 11160 2504 11212
rect 2556 11200 2562 11212
rect 2593 11203 2651 11209
rect 2593 11200 2605 11203
rect 2556 11172 2605 11200
rect 2556 11160 2562 11172
rect 2593 11169 2605 11172
rect 2639 11169 2651 11203
rect 2593 11163 2651 11169
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11200 11207 11203
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11195 11172 11989 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 11977 11169 11989 11172
rect 12023 11200 12035 11203
rect 12526 11200 12532 11212
rect 12023 11172 12532 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11200 13231 11203
rect 13998 11200 14004 11212
rect 13219 11172 14004 11200
rect 13219 11169 13231 11172
rect 13173 11163 13231 11169
rect 13998 11160 14004 11172
rect 14056 11200 14062 11212
rect 15764 11209 15792 11308
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 16850 11336 16856 11348
rect 16811 11308 16856 11336
rect 16850 11296 16856 11308
rect 16908 11336 16914 11348
rect 17313 11339 17371 11345
rect 17313 11336 17325 11339
rect 16908 11308 17325 11336
rect 16908 11296 16914 11308
rect 17313 11305 17325 11308
rect 17359 11336 17371 11339
rect 17586 11336 17592 11348
rect 17359 11308 17592 11336
rect 17359 11305 17371 11308
rect 17313 11299 17371 11305
rect 17586 11296 17592 11308
rect 17644 11336 17650 11348
rect 18601 11339 18659 11345
rect 18601 11336 18613 11339
rect 17644 11308 18613 11336
rect 17644 11296 17650 11308
rect 18601 11305 18613 11308
rect 18647 11305 18659 11339
rect 20346 11336 20352 11348
rect 20307 11308 20352 11336
rect 18601 11299 18659 11305
rect 20346 11296 20352 11308
rect 20404 11336 20410 11348
rect 21269 11339 21327 11345
rect 21269 11336 21281 11339
rect 20404 11308 21281 11336
rect 20404 11296 20410 11308
rect 21269 11305 21281 11308
rect 21315 11336 21327 11339
rect 22189 11339 22247 11345
rect 22189 11336 22201 11339
rect 21315 11308 22201 11336
rect 21315 11305 21327 11308
rect 21269 11299 21327 11305
rect 22189 11305 22201 11308
rect 22235 11305 22247 11339
rect 25958 11336 25964 11348
rect 22189 11299 22247 11305
rect 24964 11308 25964 11336
rect 15930 11268 15936 11280
rect 15856 11240 15936 11268
rect 15749 11203 15807 11209
rect 14056 11172 15700 11200
rect 14056 11160 14062 11172
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2777 11135 2835 11141
rect 2777 11132 2789 11135
rect 2280 11104 2789 11132
rect 2280 11092 2286 11104
rect 2777 11101 2789 11104
rect 2823 11101 2835 11135
rect 2777 11095 2835 11101
rect 10502 11092 10508 11144
rect 10560 11132 10566 11144
rect 10778 11132 10784 11144
rect 10560 11104 10784 11132
rect 10560 11092 10566 11104
rect 10778 11092 10784 11104
rect 10836 11132 10842 11144
rect 10965 11135 11023 11141
rect 10965 11132 10977 11135
rect 10836 11104 10977 11132
rect 10836 11092 10842 11104
rect 10965 11101 10977 11104
rect 11011 11132 11023 11135
rect 11882 11132 11888 11144
rect 11011 11104 11888 11132
rect 11011 11101 11023 11104
rect 10965 11095 11023 11101
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 13078 11132 13084 11144
rect 13035 11104 13084 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13872 11104 14197 11132
rect 13872 11092 13878 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 15565 11135 15623 11141
rect 15565 11132 15577 11135
rect 14185 11095 14243 11101
rect 15212 11104 15577 11132
rect 2501 11067 2559 11073
rect 2501 11033 2513 11067
rect 2547 11064 2559 11067
rect 2682 11064 2688 11076
rect 2547 11036 2688 11064
rect 2547 11033 2559 11036
rect 2501 11027 2559 11033
rect 2682 11024 2688 11036
rect 2740 11024 2746 11076
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 8018 11064 8024 11076
rect 4120 11036 8024 11064
rect 4120 11024 4126 11036
rect 8018 11024 8024 11036
rect 8076 11024 8082 11076
rect 11241 11067 11299 11073
rect 11241 11033 11253 11067
rect 11287 11064 11299 11067
rect 12158 11064 12164 11076
rect 11287 11036 12164 11064
rect 11287 11033 11299 11036
rect 11241 11027 11299 11033
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 15212 11008 15240 11104
rect 15565 11101 15577 11104
rect 15611 11101 15623 11135
rect 15565 11095 15623 11101
rect 15672 11064 15700 11172
rect 15749 11169 15761 11203
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 15856 11141 15884 11240
rect 15930 11228 15936 11240
rect 15988 11268 15994 11280
rect 21634 11268 21640 11280
rect 15988 11240 21640 11268
rect 15988 11228 15994 11240
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 21729 11271 21787 11277
rect 21729 11237 21741 11271
rect 21775 11268 21787 11271
rect 21775 11240 23612 11268
rect 21775 11237 21787 11240
rect 21729 11231 21787 11237
rect 21361 11203 21419 11209
rect 21361 11200 21373 11203
rect 20548 11172 21373 11200
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 17586 11092 17592 11144
rect 17644 11132 17650 11144
rect 20548 11141 20576 11172
rect 21361 11169 21373 11172
rect 21407 11169 21419 11203
rect 21361 11163 21419 11169
rect 21560 11172 21772 11200
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 17644 11104 19257 11132
rect 17644 11092 17650 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 20533 11135 20591 11141
rect 20533 11132 20545 11135
rect 19245 11095 19303 11101
rect 19444 11104 20545 11132
rect 18598 11064 18604 11076
rect 15672 11036 18604 11064
rect 18598 11024 18604 11036
rect 18656 11024 18662 11076
rect 19444 11008 19472 11104
rect 20533 11101 20545 11104
rect 20579 11101 20591 11135
rect 20533 11095 20591 11101
rect 20622 11092 20628 11144
rect 20680 11132 20686 11144
rect 21560 11141 21588 11172
rect 21545 11135 21603 11141
rect 20680 11104 21404 11132
rect 20680 11092 20686 11104
rect 20254 11024 20260 11076
rect 20312 11064 20318 11076
rect 20349 11067 20407 11073
rect 20349 11064 20361 11067
rect 20312 11036 20361 11064
rect 20312 11024 20318 11036
rect 20349 11033 20361 11036
rect 20395 11064 20407 11067
rect 21269 11067 21327 11073
rect 21269 11064 21281 11067
rect 20395 11036 21281 11064
rect 20395 11033 20407 11036
rect 20349 11027 20407 11033
rect 21269 11033 21281 11036
rect 21315 11033 21327 11067
rect 21376 11064 21404 11104
rect 21545 11101 21557 11135
rect 21591 11101 21603 11135
rect 21744 11132 21772 11172
rect 22002 11160 22008 11212
rect 22060 11200 22066 11212
rect 22281 11203 22339 11209
rect 22281 11200 22293 11203
rect 22060 11172 22293 11200
rect 22060 11160 22066 11172
rect 22281 11169 22293 11172
rect 22327 11169 22339 11203
rect 22281 11163 22339 11169
rect 23584 11141 23612 11240
rect 24964 11209 24992 11308
rect 25958 11296 25964 11308
rect 26016 11336 26022 11348
rect 28629 11339 28687 11345
rect 28629 11336 28641 11339
rect 26016 11308 28641 11336
rect 26016 11296 26022 11308
rect 28629 11305 28641 11308
rect 28675 11336 28687 11339
rect 30282 11336 30288 11348
rect 28675 11308 30288 11336
rect 28675 11305 28687 11308
rect 28629 11299 28687 11305
rect 30282 11296 30288 11308
rect 30340 11296 30346 11348
rect 32861 11339 32919 11345
rect 32861 11305 32873 11339
rect 32907 11336 32919 11339
rect 33870 11336 33876 11348
rect 32907 11308 33876 11336
rect 32907 11305 32919 11308
rect 32861 11299 32919 11305
rect 33870 11296 33876 11308
rect 33928 11336 33934 11348
rect 34698 11336 34704 11348
rect 33928 11308 34704 11336
rect 33928 11296 33934 11308
rect 34698 11296 34704 11308
rect 34756 11296 34762 11348
rect 30098 11228 30104 11280
rect 30156 11268 30162 11280
rect 30745 11271 30803 11277
rect 30745 11268 30757 11271
rect 30156 11240 30757 11268
rect 30156 11228 30162 11240
rect 30745 11237 30757 11240
rect 30791 11237 30803 11271
rect 30745 11231 30803 11237
rect 24949 11203 25007 11209
rect 24949 11169 24961 11203
rect 24995 11169 25007 11203
rect 24949 11163 25007 11169
rect 25222 11160 25228 11212
rect 25280 11200 25286 11212
rect 25409 11203 25467 11209
rect 25409 11200 25421 11203
rect 25280 11172 25421 11200
rect 25280 11160 25286 11172
rect 25409 11169 25421 11172
rect 25455 11169 25467 11203
rect 25409 11163 25467 11169
rect 22465 11135 22523 11141
rect 22465 11132 22477 11135
rect 21744 11104 22477 11132
rect 21545 11095 21603 11101
rect 22465 11101 22477 11104
rect 22511 11101 22523 11135
rect 22465 11095 22523 11101
rect 23569 11135 23627 11141
rect 23569 11101 23581 11135
rect 23615 11101 23627 11135
rect 23569 11095 23627 11101
rect 27249 11135 27307 11141
rect 27249 11101 27261 11135
rect 27295 11132 27307 11135
rect 28994 11132 29000 11144
rect 27295 11104 29000 11132
rect 27295 11101 27307 11104
rect 27249 11095 27307 11101
rect 21560 11064 21588 11095
rect 28994 11092 29000 11104
rect 29052 11132 29058 11144
rect 29052 11104 29684 11132
rect 29052 11092 29058 11104
rect 21376 11036 21588 11064
rect 21269 11027 21327 11033
rect 21634 11024 21640 11076
rect 21692 11064 21698 11076
rect 22186 11064 22192 11076
rect 21692 11036 22192 11064
rect 21692 11024 21698 11036
rect 22186 11024 22192 11036
rect 22244 11024 22250 11076
rect 25133 11067 25191 11073
rect 25133 11064 25145 11067
rect 23768 11036 25145 11064
rect 2961 10999 3019 11005
rect 2961 10965 2973 10999
rect 3007 10996 3019 10999
rect 3050 10996 3056 11008
rect 3007 10968 3056 10996
rect 3007 10965 3019 10968
rect 2961 10959 3019 10965
rect 3050 10956 3056 10968
rect 3108 10956 3114 11008
rect 11698 10996 11704 11008
rect 11659 10968 11704 10996
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 13170 10956 13176 11008
rect 13228 10996 13234 11008
rect 14369 10999 14427 11005
rect 14369 10996 14381 10999
rect 13228 10968 14381 10996
rect 13228 10956 13234 10968
rect 14369 10965 14381 10968
rect 14415 10996 14427 10999
rect 15194 10996 15200 11008
rect 14415 10968 15200 10996
rect 14415 10965 14427 10968
rect 14369 10959 14427 10965
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 19426 10996 19432 11008
rect 19387 10968 19432 10996
rect 19426 10956 19432 10968
rect 19484 10956 19490 11008
rect 20806 10996 20812 11008
rect 20767 10968 20812 10996
rect 20806 10956 20812 10968
rect 20864 10956 20870 11008
rect 22646 10996 22652 11008
rect 22607 10968 22652 10996
rect 22646 10956 22652 10968
rect 22704 10956 22710 11008
rect 23768 11005 23796 11036
rect 25133 11033 25145 11036
rect 25179 11033 25191 11067
rect 25133 11027 25191 11033
rect 27154 11024 27160 11076
rect 27212 11064 27218 11076
rect 27494 11067 27552 11073
rect 27494 11064 27506 11067
rect 27212 11036 27506 11064
rect 27212 11024 27218 11036
rect 27494 11033 27506 11036
rect 27540 11033 27552 11067
rect 27494 11027 27552 11033
rect 29656 11005 29684 11104
rect 30374 11092 30380 11144
rect 30432 11132 30438 11144
rect 32677 11135 32735 11141
rect 32677 11132 32689 11135
rect 30432 11104 32689 11132
rect 30432 11092 30438 11104
rect 32677 11101 32689 11104
rect 32723 11101 32735 11135
rect 32677 11095 32735 11101
rect 23753 10999 23811 11005
rect 23753 10965 23765 10999
rect 23799 10965 23811 10999
rect 23753 10959 23811 10965
rect 29641 10999 29699 11005
rect 29641 10965 29653 10999
rect 29687 10996 29699 10999
rect 29914 10996 29920 11008
rect 29687 10968 29920 10996
rect 29687 10965 29699 10968
rect 29641 10959 29699 10965
rect 29914 10956 29920 10968
rect 29972 10956 29978 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 4525 10795 4583 10801
rect 4525 10761 4537 10795
rect 4571 10792 4583 10795
rect 15286 10792 15292 10804
rect 4571 10764 15292 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 16022 10792 16028 10804
rect 15979 10764 16028 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 10686 10684 10692 10736
rect 10744 10724 10750 10736
rect 10781 10727 10839 10733
rect 10781 10724 10793 10727
rect 10744 10696 10793 10724
rect 10744 10684 10750 10696
rect 10781 10693 10793 10696
rect 10827 10724 10839 10727
rect 12158 10724 12164 10736
rect 10827 10696 12164 10724
rect 10827 10693 10839 10696
rect 10781 10687 10839 10693
rect 12158 10684 12164 10696
rect 12216 10724 12222 10736
rect 12529 10727 12587 10733
rect 12529 10724 12541 10727
rect 12216 10696 12541 10724
rect 12216 10684 12222 10696
rect 12529 10693 12541 10696
rect 12575 10693 12587 10727
rect 12529 10687 12587 10693
rect 12894 10684 12900 10736
rect 12952 10724 12958 10736
rect 13449 10727 13507 10733
rect 13449 10724 13461 10727
rect 12952 10696 13461 10724
rect 12952 10684 12958 10696
rect 13449 10693 13461 10696
rect 13495 10724 13507 10727
rect 14921 10727 14979 10733
rect 14921 10724 14933 10727
rect 13495 10696 14933 10724
rect 13495 10693 13507 10696
rect 13449 10687 13507 10693
rect 14921 10693 14933 10696
rect 14967 10724 14979 10727
rect 15010 10724 15016 10736
rect 14967 10696 15016 10724
rect 14967 10693 14979 10696
rect 14921 10687 14979 10693
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 15948 10724 15976 10755
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 22097 10795 22155 10801
rect 22097 10761 22109 10795
rect 22143 10792 22155 10795
rect 22186 10792 22192 10804
rect 22143 10764 22192 10792
rect 22143 10761 22155 10764
rect 22097 10755 22155 10761
rect 22186 10752 22192 10764
rect 22244 10752 22250 10804
rect 30374 10792 30380 10804
rect 30335 10764 30380 10792
rect 30374 10752 30380 10764
rect 30432 10752 30438 10804
rect 31113 10795 31171 10801
rect 31113 10761 31125 10795
rect 31159 10792 31171 10795
rect 31662 10792 31668 10804
rect 31159 10764 31668 10792
rect 31159 10761 31171 10764
rect 31113 10755 31171 10761
rect 31662 10752 31668 10764
rect 31720 10752 31726 10804
rect 18046 10724 18052 10736
rect 15120 10696 15976 10724
rect 17420 10696 18052 10724
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10656 1458 10668
rect 2041 10659 2099 10665
rect 2041 10656 2053 10659
rect 1452 10628 2053 10656
rect 1452 10616 1458 10628
rect 2041 10625 2053 10628
rect 2087 10625 2099 10659
rect 2866 10656 2872 10668
rect 2827 10628 2872 10656
rect 2041 10619 2099 10625
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 2958 10616 2964 10668
rect 3016 10656 3022 10668
rect 3099 10659 3157 10665
rect 3099 10656 3111 10659
rect 3016 10628 3111 10656
rect 3016 10616 3022 10628
rect 3099 10625 3111 10628
rect 3145 10625 3157 10659
rect 3099 10619 3157 10625
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3384 10628 4077 10656
rect 3384 10616 3390 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4614 10656 4620 10668
rect 4387 10628 4620 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 10502 10656 10508 10668
rect 10463 10628 10508 10656
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10656 12311 10659
rect 13170 10656 13176 10668
rect 12299 10628 13176 10656
rect 12299 10625 12311 10628
rect 12253 10619 12311 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 13998 10656 14004 10668
rect 13959 10628 14004 10656
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 15120 10665 15148 10696
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 17420 10665 17448 10696
rect 18046 10684 18052 10696
rect 18104 10684 18110 10736
rect 18598 10684 18604 10736
rect 18656 10724 18662 10736
rect 29733 10727 29791 10733
rect 18656 10696 20208 10724
rect 18656 10684 18662 10696
rect 17405 10659 17463 10665
rect 15252 10628 15297 10656
rect 15252 10616 15258 10628
rect 17405 10625 17417 10659
rect 17451 10625 17463 10659
rect 17586 10656 17592 10668
rect 17547 10628 17592 10656
rect 17405 10619 17463 10625
rect 17586 10616 17592 10628
rect 17644 10616 17650 10668
rect 17862 10656 17868 10668
rect 17823 10628 17868 10656
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 18414 10656 18420 10668
rect 18375 10628 18420 10656
rect 18414 10616 18420 10628
rect 18472 10616 18478 10668
rect 20180 10665 20208 10696
rect 29733 10693 29745 10727
rect 29779 10724 29791 10727
rect 30098 10724 30104 10736
rect 29779 10696 30104 10724
rect 29779 10693 29791 10696
rect 29733 10687 29791 10693
rect 30098 10684 30104 10696
rect 30156 10724 30162 10736
rect 30285 10727 30343 10733
rect 30285 10724 30297 10727
rect 30156 10696 30297 10724
rect 30156 10684 30162 10696
rect 30285 10693 30297 10696
rect 30331 10724 30343 10727
rect 30331 10696 30972 10724
rect 30331 10693 30343 10696
rect 30285 10687 30343 10693
rect 30944 10668 30972 10696
rect 19521 10659 19579 10665
rect 19521 10656 19533 10659
rect 18524 10628 19533 10656
rect 18524 10600 18552 10628
rect 19521 10625 19533 10628
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 20165 10659 20223 10665
rect 20165 10625 20177 10659
rect 20211 10625 20223 10659
rect 20165 10619 20223 10625
rect 20806 10616 20812 10668
rect 20864 10656 20870 10668
rect 23017 10659 23075 10665
rect 23017 10656 23029 10659
rect 20864 10628 23029 10656
rect 20864 10616 20870 10628
rect 23017 10625 23029 10628
rect 23063 10625 23075 10659
rect 30926 10656 30932 10668
rect 30839 10628 30932 10656
rect 23017 10619 23075 10625
rect 30926 10616 30932 10628
rect 30984 10616 30990 10668
rect 34698 10656 34704 10668
rect 34659 10628 34704 10656
rect 34698 10616 34704 10628
rect 34756 10616 34762 10668
rect 34790 10616 34796 10668
rect 34848 10656 34854 10668
rect 34885 10659 34943 10665
rect 34885 10656 34897 10659
rect 34848 10628 34897 10656
rect 34848 10616 34854 10628
rect 34885 10625 34897 10628
rect 34931 10625 34943 10659
rect 34885 10619 34943 10625
rect 1946 10548 1952 10600
rect 2004 10588 2010 10600
rect 3237 10591 3295 10597
rect 3237 10588 3249 10591
rect 2004 10560 3249 10588
rect 2004 10548 2010 10560
rect 3237 10557 3249 10560
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 3970 10548 3976 10600
rect 4028 10588 4034 10600
rect 4157 10591 4215 10597
rect 4157 10588 4169 10591
rect 4028 10560 4169 10588
rect 4028 10548 4034 10560
rect 4157 10557 4169 10560
rect 4203 10557 4215 10591
rect 9306 10588 9312 10600
rect 9267 10560 9312 10588
rect 4157 10551 4215 10557
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10588 10747 10591
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 10735 10560 12449 10588
rect 10735 10557 10747 10560
rect 10689 10551 10747 10557
rect 12437 10557 12449 10560
rect 12483 10588 12495 10591
rect 12526 10588 12532 10600
rect 12483 10560 12532 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 2498 10520 2504 10532
rect 1627 10492 2504 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 2498 10480 2504 10492
rect 2556 10480 2562 10532
rect 3513 10523 3571 10529
rect 3513 10489 3525 10523
rect 3559 10520 3571 10523
rect 4706 10520 4712 10532
rect 3559 10492 4712 10520
rect 3559 10489 3571 10492
rect 3513 10483 3571 10489
rect 4706 10480 4712 10492
rect 4764 10480 4770 10532
rect 9600 10520 9628 10551
rect 12526 10548 12532 10560
rect 12584 10588 12590 10600
rect 13265 10591 13323 10597
rect 13265 10588 13277 10591
rect 12584 10560 13277 10588
rect 12584 10548 12590 10560
rect 13265 10557 13277 10560
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 18506 10588 18512 10600
rect 13872 10560 18512 10588
rect 13872 10548 13878 10560
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 10321 10523 10379 10529
rect 10321 10520 10333 10523
rect 9600 10492 10333 10520
rect 10321 10489 10333 10492
rect 10367 10489 10379 10523
rect 17218 10520 17224 10532
rect 10321 10483 10379 10489
rect 12544 10492 13492 10520
rect 17179 10492 17224 10520
rect 3050 10461 3056 10464
rect 3034 10455 3056 10461
rect 3034 10421 3046 10455
rect 3034 10415 3056 10421
rect 3050 10412 3056 10415
rect 3108 10412 3114 10464
rect 4062 10452 4068 10464
rect 4023 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 10594 10452 10600 10464
rect 10555 10424 10600 10452
rect 10594 10412 10600 10424
rect 10652 10412 10658 10464
rect 12066 10452 12072 10464
rect 12027 10424 12072 10452
rect 12066 10412 12072 10424
rect 12124 10412 12130 10464
rect 12544 10461 12572 10492
rect 12529 10455 12587 10461
rect 12529 10421 12541 10455
rect 12575 10421 12587 10455
rect 12529 10415 12587 10421
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 13464 10461 13492 10492
rect 17218 10480 17224 10492
rect 17276 10480 17282 10532
rect 34330 10480 34336 10532
rect 34388 10520 34394 10532
rect 34701 10523 34759 10529
rect 34701 10520 34713 10523
rect 34388 10492 34713 10520
rect 34388 10480 34394 10492
rect 34701 10489 34713 10492
rect 34747 10489 34759 10523
rect 34701 10483 34759 10489
rect 12989 10455 13047 10461
rect 12989 10452 13001 10455
rect 12768 10424 13001 10452
rect 12768 10412 12774 10424
rect 12989 10421 13001 10424
rect 13035 10421 13047 10455
rect 12989 10415 13047 10421
rect 13449 10455 13507 10461
rect 13449 10421 13461 10455
rect 13495 10452 13507 10455
rect 14185 10455 14243 10461
rect 14185 10452 14197 10455
rect 13495 10424 14197 10452
rect 13495 10421 13507 10424
rect 13449 10415 13507 10421
rect 14185 10421 14197 10424
rect 14231 10452 14243 10455
rect 15102 10452 15108 10464
rect 14231 10424 15108 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 15102 10412 15108 10424
rect 15160 10412 15166 10464
rect 15381 10455 15439 10461
rect 15381 10421 15393 10455
rect 15427 10452 15439 10455
rect 15470 10452 15476 10464
rect 15427 10424 15476 10452
rect 15427 10421 15439 10424
rect 15381 10415 15439 10421
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 19702 10452 19708 10464
rect 19663 10424 19708 10452
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 20346 10452 20352 10464
rect 20307 10424 20352 10452
rect 20346 10412 20352 10424
rect 20404 10412 20410 10464
rect 23201 10455 23259 10461
rect 23201 10421 23213 10455
rect 23247 10452 23259 10455
rect 26050 10452 26056 10464
rect 23247 10424 26056 10452
rect 23247 10421 23259 10424
rect 23201 10415 23259 10421
rect 26050 10412 26056 10424
rect 26108 10412 26114 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1946 10248 1952 10260
rect 1907 10220 1952 10248
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2501 10251 2559 10257
rect 2501 10248 2513 10251
rect 2280 10220 2513 10248
rect 2280 10208 2286 10220
rect 2501 10217 2513 10220
rect 2547 10217 2559 10251
rect 2501 10211 2559 10217
rect 2961 10251 3019 10257
rect 2961 10217 2973 10251
rect 3007 10248 3019 10251
rect 4062 10248 4068 10260
rect 3007 10220 4068 10248
rect 3007 10217 3019 10220
rect 2961 10211 3019 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4706 10208 4712 10260
rect 4764 10248 4770 10260
rect 4764 10220 6316 10248
rect 4764 10208 4770 10220
rect 6288 10180 6316 10220
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 12437 10251 12495 10257
rect 12437 10248 12449 10251
rect 11940 10220 12449 10248
rect 11940 10208 11946 10220
rect 12437 10217 12449 10220
rect 12483 10217 12495 10251
rect 15102 10248 15108 10260
rect 15063 10220 15108 10248
rect 12437 10211 12495 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 16022 10248 16028 10260
rect 15983 10220 16028 10248
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 19705 10251 19763 10257
rect 19705 10217 19717 10251
rect 19751 10248 19763 10251
rect 20346 10248 20352 10260
rect 19751 10220 20352 10248
rect 19751 10217 19763 10220
rect 19705 10211 19763 10217
rect 20346 10208 20352 10220
rect 20404 10248 20410 10260
rect 20625 10251 20683 10257
rect 20625 10248 20637 10251
rect 20404 10220 20637 10248
rect 20404 10208 20410 10220
rect 20625 10217 20637 10220
rect 20671 10248 20683 10251
rect 21269 10251 21327 10257
rect 21269 10248 21281 10251
rect 20671 10220 21281 10248
rect 20671 10217 20683 10220
rect 20625 10211 20683 10217
rect 21269 10217 21281 10220
rect 21315 10217 21327 10251
rect 21269 10211 21327 10217
rect 6288 10152 12434 10180
rect 2590 10112 2596 10124
rect 2551 10084 2596 10112
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 11054 10112 11060 10124
rect 11015 10084 11060 10112
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 2498 10044 2504 10056
rect 2459 10016 2504 10044
rect 1857 10007 1915 10013
rect 1872 9976 1900 10007
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 2832 10016 2877 10044
rect 2832 10004 2838 10016
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 5261 10047 5319 10053
rect 5261 10044 5273 10047
rect 3936 10016 5273 10044
rect 3936 10004 3942 10016
rect 5261 10013 5273 10016
rect 5307 10044 5319 10047
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 5307 10016 7113 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 10134 10044 10140 10056
rect 10095 10016 10140 10044
rect 7101 10007 7159 10013
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 2590 9976 2596 9988
rect 1872 9948 2596 9976
rect 2590 9936 2596 9948
rect 2648 9936 2654 9988
rect 5534 9985 5540 9988
rect 5528 9939 5540 9985
rect 5592 9976 5598 9988
rect 10318 9976 10324 9988
rect 5592 9948 5628 9976
rect 10279 9948 10324 9976
rect 5534 9936 5540 9939
rect 5592 9936 5598 9948
rect 10318 9936 10324 9948
rect 10376 9936 10382 9988
rect 12406 9976 12434 10152
rect 15197 10115 15255 10121
rect 15197 10081 15209 10115
rect 15243 10112 15255 10115
rect 16040 10112 16068 10208
rect 15243 10084 16068 10112
rect 15243 10081 15255 10084
rect 15197 10075 15255 10081
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19521 10115 19579 10121
rect 19521 10112 19533 10115
rect 19484 10084 19533 10112
rect 19484 10072 19490 10084
rect 19521 10081 19533 10084
rect 19567 10112 19579 10115
rect 20441 10115 20499 10121
rect 20441 10112 20453 10115
rect 19567 10084 20453 10112
rect 19567 10081 19579 10084
rect 19521 10075 19579 10081
rect 20441 10081 20453 10084
rect 20487 10112 20499 10115
rect 21361 10115 21419 10121
rect 21361 10112 21373 10115
rect 20487 10084 21373 10112
rect 20487 10081 20499 10084
rect 20441 10075 20499 10081
rect 21361 10081 21373 10084
rect 21407 10081 21419 10115
rect 24394 10112 24400 10124
rect 24355 10084 24400 10112
rect 21361 10075 21419 10081
rect 24394 10072 24400 10084
rect 24452 10072 24458 10124
rect 26050 10112 26056 10124
rect 26011 10084 26056 10112
rect 26050 10072 26056 10084
rect 26108 10072 26114 10124
rect 30282 10072 30288 10124
rect 30340 10112 30346 10124
rect 30469 10115 30527 10121
rect 30469 10112 30481 10115
rect 30340 10084 30481 10112
rect 30340 10072 30346 10084
rect 30469 10081 30481 10084
rect 30515 10081 30527 10115
rect 31294 10112 31300 10124
rect 30469 10075 30527 10081
rect 30944 10084 31300 10112
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10044 12679 10047
rect 13814 10044 13820 10056
rect 12667 10016 13820 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 15010 10044 15016 10056
rect 14971 10016 15016 10044
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 15286 10044 15292 10056
rect 15247 10016 15292 10044
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 19702 10044 19708 10056
rect 19663 10016 19708 10044
rect 19702 10004 19708 10016
rect 19760 10044 19766 10056
rect 20625 10047 20683 10053
rect 20625 10044 20637 10047
rect 19760 10016 20637 10044
rect 19760 10004 19766 10016
rect 20625 10013 20637 10016
rect 20671 10044 20683 10047
rect 20806 10044 20812 10056
rect 20671 10016 20812 10044
rect 20671 10013 20683 10016
rect 20625 10007 20683 10013
rect 20806 10004 20812 10016
rect 20864 10044 20870 10056
rect 21545 10047 21603 10053
rect 21545 10044 21557 10047
rect 20864 10016 21557 10044
rect 20864 10004 20870 10016
rect 21545 10013 21557 10016
rect 21591 10013 21603 10047
rect 21545 10007 21603 10013
rect 26237 10047 26295 10053
rect 26237 10013 26249 10047
rect 26283 10044 26295 10047
rect 30834 10044 30840 10056
rect 26283 10016 30840 10044
rect 26283 10013 26295 10016
rect 26237 10007 26295 10013
rect 30834 10004 30840 10016
rect 30892 10004 30898 10056
rect 30944 10053 30972 10084
rect 31294 10072 31300 10084
rect 31352 10112 31358 10124
rect 31352 10084 31708 10112
rect 31352 10072 31358 10084
rect 30929 10047 30987 10053
rect 30929 10013 30941 10047
rect 30975 10013 30987 10047
rect 31478 10044 31484 10056
rect 31439 10016 31484 10044
rect 30929 10007 30987 10013
rect 31478 10004 31484 10016
rect 31536 10004 31542 10056
rect 31680 10053 31708 10084
rect 31665 10047 31723 10053
rect 31665 10013 31677 10047
rect 31711 10044 31723 10047
rect 34330 10044 34336 10056
rect 31711 10016 34336 10044
rect 31711 10013 31723 10016
rect 31665 10007 31723 10013
rect 34330 10004 34336 10016
rect 34388 10004 34394 10056
rect 34977 10047 35035 10053
rect 34977 10044 34989 10047
rect 34532 10016 34989 10044
rect 16945 9979 17003 9985
rect 16945 9976 16957 9979
rect 12406 9948 16957 9976
rect 16945 9945 16957 9948
rect 16991 9976 17003 9979
rect 17862 9976 17868 9988
rect 16991 9948 17868 9976
rect 16991 9945 17003 9948
rect 16945 9939 17003 9945
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 19429 9979 19487 9985
rect 19429 9945 19441 9979
rect 19475 9976 19487 9979
rect 20254 9976 20260 9988
rect 19475 9948 20260 9976
rect 19475 9945 19487 9948
rect 19429 9939 19487 9945
rect 20254 9936 20260 9948
rect 20312 9936 20318 9988
rect 20349 9979 20407 9985
rect 20349 9945 20361 9979
rect 20395 9976 20407 9979
rect 20438 9976 20444 9988
rect 20395 9948 20444 9976
rect 20395 9945 20407 9948
rect 20349 9939 20407 9945
rect 20438 9936 20444 9948
rect 20496 9976 20502 9988
rect 21269 9979 21327 9985
rect 21269 9976 21281 9979
rect 20496 9948 21281 9976
rect 20496 9936 20502 9948
rect 21269 9945 21281 9948
rect 21315 9945 21327 9979
rect 31386 9976 31392 9988
rect 31347 9948 31392 9976
rect 21269 9939 21327 9945
rect 31386 9936 31392 9948
rect 31444 9936 31450 9988
rect 34532 9920 34560 10016
rect 34977 10013 34989 10016
rect 35023 10013 35035 10047
rect 38102 10044 38108 10056
rect 38063 10016 38108 10044
rect 34977 10007 35035 10013
rect 38102 10004 38108 10016
rect 38160 10004 38166 10056
rect 35066 9936 35072 9988
rect 35124 9976 35130 9988
rect 35222 9979 35280 9985
rect 35222 9976 35234 9979
rect 35124 9948 35234 9976
rect 35124 9936 35130 9948
rect 35222 9945 35234 9948
rect 35268 9945 35280 9979
rect 35222 9939 35280 9945
rect 6546 9868 6552 9920
rect 6604 9908 6610 9920
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 6604 9880 6653 9908
rect 6604 9868 6610 9880
rect 6641 9877 6653 9880
rect 6687 9908 6699 9911
rect 10134 9908 10140 9920
rect 6687 9880 10140 9908
rect 6687 9877 6699 9880
rect 6641 9871 6699 9877
rect 10134 9868 10140 9880
rect 10192 9868 10198 9920
rect 13078 9908 13084 9920
rect 13039 9880 13084 9908
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 15473 9911 15531 9917
rect 15473 9877 15485 9911
rect 15519 9908 15531 9911
rect 15838 9908 15844 9920
rect 15519 9880 15844 9908
rect 15519 9877 15531 9880
rect 15473 9871 15531 9877
rect 15838 9868 15844 9880
rect 15896 9868 15902 9920
rect 18414 9868 18420 9920
rect 18472 9908 18478 9920
rect 18598 9908 18604 9920
rect 18472 9880 18604 9908
rect 18472 9868 18478 9880
rect 18598 9868 18604 9880
rect 18656 9868 18662 9920
rect 19889 9911 19947 9917
rect 19889 9877 19901 9911
rect 19935 9908 19947 9911
rect 19978 9908 19984 9920
rect 19935 9880 19984 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 19978 9868 19984 9880
rect 20036 9868 20042 9920
rect 20809 9911 20867 9917
rect 20809 9877 20821 9911
rect 20855 9908 20867 9911
rect 21542 9908 21548 9920
rect 20855 9880 21548 9908
rect 20855 9877 20867 9880
rect 20809 9871 20867 9877
rect 21542 9868 21548 9880
rect 21600 9868 21606 9920
rect 21726 9908 21732 9920
rect 21687 9880 21732 9908
rect 21726 9868 21732 9880
rect 21784 9868 21790 9920
rect 29914 9908 29920 9920
rect 29875 9880 29920 9908
rect 29914 9868 29920 9880
rect 29972 9868 29978 9920
rect 30742 9908 30748 9920
rect 30703 9880 30748 9908
rect 30742 9868 30748 9880
rect 30800 9868 30806 9920
rect 34149 9911 34207 9917
rect 34149 9877 34161 9911
rect 34195 9908 34207 9911
rect 34514 9908 34520 9920
rect 34195 9880 34520 9908
rect 34195 9877 34207 9880
rect 34149 9871 34207 9877
rect 34514 9868 34520 9880
rect 34572 9868 34578 9920
rect 36354 9908 36360 9920
rect 36315 9880 36360 9908
rect 36354 9868 36360 9880
rect 36412 9868 36418 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 2774 9704 2780 9716
rect 2746 9664 2780 9704
rect 2832 9664 2838 9716
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 2961 9707 3019 9713
rect 2961 9704 2973 9707
rect 2924 9676 2973 9704
rect 2924 9664 2930 9676
rect 2961 9673 2973 9676
rect 3007 9673 3019 9707
rect 2961 9667 3019 9673
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 5810 9704 5816 9716
rect 4120 9676 5816 9704
rect 4120 9664 4126 9676
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 10318 9664 10324 9716
rect 10376 9704 10382 9716
rect 10689 9707 10747 9713
rect 10689 9704 10701 9707
rect 10376 9676 10701 9704
rect 10376 9664 10382 9676
rect 10689 9673 10701 9676
rect 10735 9673 10747 9707
rect 10689 9667 10747 9673
rect 28368 9676 28580 9704
rect 2746 9636 2774 9664
rect 3605 9639 3663 9645
rect 3605 9636 3617 9639
rect 2516 9608 2774 9636
rect 3068 9608 3617 9636
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 2516 9577 2544 9608
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 1596 9540 2513 9568
rect 1596 9441 1624 9540
rect 2501 9537 2513 9540
rect 2547 9537 2559 9571
rect 2501 9531 2559 9537
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9568 2835 9571
rect 3068 9568 3096 9608
rect 3605 9605 3617 9608
rect 3651 9605 3663 9639
rect 3605 9599 3663 9605
rect 3789 9639 3847 9645
rect 3789 9605 3801 9639
rect 3835 9636 3847 9639
rect 4614 9636 4620 9648
rect 3835 9608 4620 9636
rect 3835 9605 3847 9608
rect 3789 9599 3847 9605
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 7837 9639 7895 9645
rect 7837 9605 7849 9639
rect 7883 9636 7895 9639
rect 9306 9636 9312 9648
rect 7883 9608 9312 9636
rect 7883 9605 7895 9608
rect 7837 9599 7895 9605
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 20438 9596 20444 9648
rect 20496 9636 20502 9648
rect 20533 9639 20591 9645
rect 20533 9636 20545 9639
rect 20496 9608 20545 9636
rect 20496 9596 20502 9608
rect 20533 9605 20545 9608
rect 20579 9605 20591 9639
rect 20533 9599 20591 9605
rect 22094 9596 22100 9648
rect 22152 9636 22158 9648
rect 28368 9636 28396 9676
rect 22152 9608 28396 9636
rect 28552 9636 28580 9676
rect 30834 9664 30840 9716
rect 30892 9704 30898 9716
rect 31389 9707 31447 9713
rect 31389 9704 31401 9707
rect 30892 9676 31401 9704
rect 30892 9664 30898 9676
rect 31389 9673 31401 9676
rect 31435 9673 31447 9707
rect 34790 9704 34796 9716
rect 31389 9667 31447 9673
rect 34440 9676 34796 9704
rect 29365 9639 29423 9645
rect 29365 9636 29377 9639
rect 28552 9608 29377 9636
rect 22152 9596 22158 9608
rect 29365 9605 29377 9608
rect 29411 9605 29423 9639
rect 29365 9599 29423 9605
rect 33597 9639 33655 9645
rect 33597 9605 33609 9639
rect 33643 9636 33655 9639
rect 34440 9636 34468 9676
rect 34790 9664 34796 9676
rect 34848 9664 34854 9716
rect 33643 9608 34468 9636
rect 34517 9639 34575 9645
rect 33643 9605 33655 9608
rect 33597 9599 33655 9605
rect 34517 9605 34529 9639
rect 34563 9636 34575 9639
rect 35066 9636 35072 9648
rect 34563 9608 35072 9636
rect 34563 9605 34575 9608
rect 34517 9599 34575 9605
rect 35066 9596 35072 9608
rect 35124 9596 35130 9648
rect 35244 9639 35302 9645
rect 35244 9605 35256 9639
rect 35290 9636 35302 9639
rect 35342 9636 35348 9648
rect 35290 9608 35348 9636
rect 35290 9605 35302 9608
rect 35244 9599 35302 9605
rect 35342 9596 35348 9608
rect 35400 9596 35406 9648
rect 2823 9540 3096 9568
rect 3421 9571 3479 9577
rect 2823 9537 2835 9540
rect 2777 9531 2835 9537
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 5626 9568 5632 9580
rect 5587 9540 5632 9568
rect 3421 9531 3479 9537
rect 2682 9500 2688 9512
rect 2643 9472 2688 9500
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9401 1639 9435
rect 1581 9395 1639 9401
rect 2406 9392 2412 9444
rect 2464 9432 2470 9444
rect 2792 9432 2820 9531
rect 3436 9500 3464 9531
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 10870 9568 10876 9580
rect 10831 9540 10876 9568
rect 10870 9528 10876 9540
rect 10928 9528 10934 9580
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9568 11575 9571
rect 12066 9568 12072 9580
rect 11563 9540 12072 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 12066 9528 12072 9540
rect 12124 9528 12130 9580
rect 15470 9568 15476 9580
rect 15431 9540 15476 9568
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 15838 9528 15844 9580
rect 15896 9568 15902 9580
rect 16117 9571 16175 9577
rect 16117 9568 16129 9571
rect 15896 9540 16129 9568
rect 15896 9528 15902 9540
rect 16117 9537 16129 9540
rect 16163 9537 16175 9571
rect 16117 9531 16175 9537
rect 20622 9528 20628 9580
rect 20680 9568 20686 9580
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 20680 9540 20729 9568
rect 20680 9528 20686 9540
rect 20717 9537 20729 9540
rect 20763 9537 20775 9571
rect 20717 9531 20775 9537
rect 20806 9528 20812 9580
rect 20864 9568 20870 9580
rect 20864 9540 20909 9568
rect 20864 9528 20870 9540
rect 22646 9528 22652 9580
rect 22704 9568 22710 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 22704 9540 23949 9568
rect 22704 9528 22710 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 28626 9568 28632 9580
rect 23937 9531 23995 9537
rect 24044 9540 28488 9568
rect 28587 9540 28632 9568
rect 2464 9404 2820 9432
rect 3068 9472 3464 9500
rect 2464 9392 2470 9404
rect 3068 9376 3096 9472
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 7653 9503 7711 9509
rect 7653 9500 7665 9503
rect 7432 9472 7665 9500
rect 7432 9460 7438 9472
rect 7653 9469 7665 9472
rect 7699 9469 7711 9503
rect 9490 9500 9496 9512
rect 9451 9472 9496 9500
rect 7653 9463 7711 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 11790 9500 11796 9512
rect 11751 9472 11796 9500
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 17402 9460 17408 9512
rect 17460 9500 17466 9512
rect 24044 9500 24072 9540
rect 17460 9472 24072 9500
rect 24213 9503 24271 9509
rect 17460 9460 17466 9472
rect 24213 9469 24225 9503
rect 24259 9500 24271 9503
rect 26602 9500 26608 9512
rect 24259 9472 26608 9500
rect 24259 9469 24271 9472
rect 24213 9463 24271 9469
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 26973 9503 27031 9509
rect 26973 9469 26985 9503
rect 27019 9469 27031 9503
rect 26973 9463 27031 9469
rect 27249 9503 27307 9509
rect 27249 9469 27261 9503
rect 27295 9500 27307 9503
rect 27522 9500 27528 9512
rect 27295 9472 27528 9500
rect 27295 9469 27307 9472
rect 27249 9463 27307 9469
rect 5445 9435 5503 9441
rect 5445 9401 5457 9435
rect 5491 9432 5503 9435
rect 5534 9432 5540 9444
rect 5491 9404 5540 9432
rect 5491 9401 5503 9404
rect 5445 9395 5503 9401
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 5810 9392 5816 9444
rect 5868 9432 5874 9444
rect 11054 9432 11060 9444
rect 5868 9404 11060 9432
rect 5868 9392 5874 9404
rect 11054 9392 11060 9404
rect 11112 9392 11118 9444
rect 20993 9435 21051 9441
rect 20993 9401 21005 9435
rect 21039 9432 21051 9435
rect 26988 9432 27016 9463
rect 27522 9460 27528 9472
rect 27580 9460 27586 9512
rect 21039 9404 27016 9432
rect 21039 9401 21051 9404
rect 20993 9395 21051 9401
rect 2777 9367 2835 9373
rect 2777 9333 2789 9367
rect 2823 9364 2835 9367
rect 3050 9364 3056 9376
rect 2823 9336 3056 9364
rect 2823 9333 2835 9336
rect 2777 9327 2835 9333
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 4890 9324 4896 9376
rect 4948 9364 4954 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 4948 9336 6377 9364
rect 4948 9324 4954 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 15286 9364 15292 9376
rect 15247 9336 15292 9364
rect 6365 9327 6423 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 15933 9367 15991 9373
rect 15933 9364 15945 9367
rect 15620 9336 15945 9364
rect 15620 9324 15626 9336
rect 15933 9333 15945 9336
rect 15979 9333 15991 9367
rect 15933 9327 15991 9333
rect 20346 9324 20352 9376
rect 20404 9364 20410 9376
rect 20533 9367 20591 9373
rect 20533 9364 20545 9367
rect 20404 9336 20545 9364
rect 20404 9324 20410 9336
rect 20533 9333 20545 9336
rect 20579 9333 20591 9367
rect 28460 9364 28488 9540
rect 28626 9528 28632 9540
rect 28684 9528 28690 9580
rect 30265 9571 30323 9577
rect 30265 9568 30277 9571
rect 28828 9540 30277 9568
rect 28828 9441 28856 9540
rect 30265 9537 30277 9540
rect 30311 9537 30323 9571
rect 33321 9571 33379 9577
rect 33321 9568 33333 9571
rect 30265 9531 30323 9537
rect 32784 9540 33333 9568
rect 29362 9460 29368 9512
rect 29420 9500 29426 9512
rect 29549 9503 29607 9509
rect 29549 9500 29561 9503
rect 29420 9472 29561 9500
rect 29420 9460 29426 9472
rect 29549 9469 29561 9472
rect 29595 9500 29607 9503
rect 29914 9500 29920 9512
rect 29595 9472 29920 9500
rect 29595 9469 29607 9472
rect 29549 9463 29607 9469
rect 29914 9460 29920 9472
rect 29972 9500 29978 9512
rect 30009 9503 30067 9509
rect 30009 9500 30021 9503
rect 29972 9472 30021 9500
rect 29972 9460 29978 9472
rect 30009 9469 30021 9472
rect 30055 9469 30067 9503
rect 30009 9463 30067 9469
rect 28813 9435 28871 9441
rect 28813 9401 28825 9435
rect 28859 9401 28871 9435
rect 28813 9395 28871 9401
rect 32784 9373 32812 9540
rect 33321 9537 33333 9540
rect 33367 9537 33379 9571
rect 33321 9531 33379 9537
rect 34057 9571 34115 9577
rect 34057 9537 34069 9571
rect 34103 9537 34115 9571
rect 34238 9568 34244 9580
rect 34199 9540 34244 9568
rect 34057 9531 34115 9537
rect 33413 9435 33471 9441
rect 33413 9401 33425 9435
rect 33459 9432 33471 9435
rect 34072 9432 34100 9531
rect 34238 9528 34244 9540
rect 34296 9528 34302 9580
rect 34422 9568 34428 9580
rect 34383 9540 34428 9568
rect 34422 9528 34428 9540
rect 34480 9528 34486 9580
rect 34330 9500 34336 9512
rect 34291 9472 34336 9500
rect 34330 9460 34336 9472
rect 34388 9460 34394 9512
rect 34514 9460 34520 9512
rect 34572 9500 34578 9512
rect 34977 9503 35035 9509
rect 34977 9500 34989 9503
rect 34572 9472 34989 9500
rect 34572 9460 34578 9472
rect 34977 9469 34989 9472
rect 35023 9469 35035 9503
rect 34977 9463 35035 9469
rect 34606 9432 34612 9444
rect 33459 9404 34008 9432
rect 34072 9404 34612 9432
rect 33459 9401 33471 9404
rect 33413 9395 33471 9401
rect 32769 9367 32827 9373
rect 32769 9364 32781 9367
rect 28460 9336 32781 9364
rect 20533 9327 20591 9333
rect 32769 9333 32781 9336
rect 32815 9333 32827 9367
rect 33502 9364 33508 9376
rect 33463 9336 33508 9364
rect 32769 9327 32827 9333
rect 33502 9324 33508 9336
rect 33560 9324 33566 9376
rect 33980 9364 34008 9404
rect 34606 9392 34612 9404
rect 34664 9392 34670 9444
rect 34698 9364 34704 9376
rect 33980 9336 34704 9364
rect 34698 9324 34704 9336
rect 34756 9364 34762 9376
rect 36357 9367 36415 9373
rect 36357 9364 36369 9367
rect 34756 9336 36369 9364
rect 34756 9324 34762 9336
rect 36357 9333 36369 9336
rect 36403 9333 36415 9367
rect 36357 9327 36415 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2961 9163 3019 9169
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 3326 9160 3332 9172
rect 3007 9132 3332 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 5537 9163 5595 9169
rect 5537 9129 5549 9163
rect 5583 9160 5595 9163
rect 5626 9160 5632 9172
rect 5583 9132 5632 9160
rect 5583 9129 5595 9132
rect 5537 9123 5595 9129
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 20625 9163 20683 9169
rect 20625 9160 20637 9163
rect 20404 9132 20637 9160
rect 20404 9120 20410 9132
rect 20625 9129 20637 9132
rect 20671 9129 20683 9163
rect 20625 9123 20683 9129
rect 28997 9163 29055 9169
rect 28997 9129 29009 9163
rect 29043 9160 29055 9163
rect 29546 9160 29552 9172
rect 29043 9132 29552 9160
rect 29043 9129 29055 9132
rect 28997 9123 29055 9129
rect 29546 9120 29552 9132
rect 29604 9120 29610 9172
rect 29914 9120 29920 9172
rect 29972 9160 29978 9172
rect 34057 9163 34115 9169
rect 34057 9160 34069 9163
rect 29972 9132 34069 9160
rect 29972 9120 29978 9132
rect 34057 9129 34069 9132
rect 34103 9160 34115 9163
rect 34514 9160 34520 9172
rect 34103 9132 34520 9160
rect 34103 9129 34115 9132
rect 34057 9123 34115 9129
rect 34514 9120 34520 9132
rect 34572 9120 34578 9172
rect 1394 9092 1400 9104
rect 1355 9064 1400 9092
rect 1394 9052 1400 9064
rect 1452 9052 1458 9104
rect 5166 9052 5172 9104
rect 5224 9092 5230 9104
rect 9490 9092 9496 9104
rect 5224 9064 9496 9092
rect 5224 9052 5230 9064
rect 9490 9052 9496 9064
rect 9548 9052 9554 9104
rect 31294 9092 31300 9104
rect 31255 9064 31300 9092
rect 31294 9052 31300 9064
rect 31352 9052 31358 9104
rect 34238 9052 34244 9104
rect 34296 9092 34302 9104
rect 35618 9092 35624 9104
rect 34296 9064 35624 9092
rect 34296 9052 34302 9064
rect 35618 9052 35624 9064
rect 35676 9092 35682 9104
rect 35989 9095 36047 9101
rect 35989 9092 36001 9095
rect 35676 9064 36001 9092
rect 35676 9052 35682 9064
rect 35989 9061 36001 9064
rect 36035 9061 36047 9095
rect 35989 9055 36047 9061
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 6549 9027 6607 9033
rect 6549 9024 6561 9027
rect 5776 8996 6561 9024
rect 5776 8984 5782 8996
rect 6549 8993 6561 8996
rect 6595 8993 6607 9027
rect 12710 9024 12716 9036
rect 12671 8996 12716 9024
rect 6549 8987 6607 8993
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 15562 9024 15568 9036
rect 15523 8996 15568 9024
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 16574 9024 16580 9036
rect 16535 8996 16580 9024
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 20622 8984 20628 9036
rect 20680 9024 20686 9036
rect 20717 9027 20775 9033
rect 20717 9024 20729 9027
rect 20680 8996 20729 9024
rect 20680 8984 20686 8996
rect 20717 8993 20729 8996
rect 20763 8993 20775 9027
rect 27062 9024 27068 9036
rect 27023 8996 27068 9024
rect 20717 8987 20775 8993
rect 27062 8984 27068 8996
rect 27120 8984 27126 9036
rect 29086 8984 29092 9036
rect 29144 9024 29150 9036
rect 29733 9027 29791 9033
rect 29733 9024 29745 9027
rect 29144 8996 29745 9024
rect 29144 8984 29150 8996
rect 29733 8993 29745 8996
rect 29779 8993 29791 9027
rect 29733 8987 29791 8993
rect 30742 8984 30748 9036
rect 30800 9024 30806 9036
rect 30800 8996 31524 9024
rect 30800 8984 30806 8996
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 4948 8928 5181 8956
rect 4948 8916 4954 8928
rect 5169 8925 5181 8928
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 5316 8928 5365 8956
rect 5316 8916 5322 8928
rect 5353 8925 5365 8928
rect 5399 8925 5411 8959
rect 10962 8956 10968 8968
rect 10923 8928 10968 8956
rect 5353 8919 5411 8925
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 11756 8928 11897 8956
rect 11756 8916 11762 8928
rect 11885 8925 11897 8928
rect 11931 8925 11943 8959
rect 11885 8919 11943 8925
rect 12618 8916 12624 8968
rect 12676 8956 12682 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12676 8928 13001 8956
rect 12676 8916 12682 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 15378 8956 15384 8968
rect 15339 8928 15384 8956
rect 12989 8919 13047 8925
rect 15378 8916 15384 8928
rect 15436 8916 15442 8968
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 19978 8956 19984 8968
rect 19935 8928 19984 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 19978 8916 19984 8928
rect 20036 8916 20042 8968
rect 20806 8916 20812 8968
rect 20864 8956 20870 8968
rect 20901 8959 20959 8965
rect 20901 8956 20913 8959
rect 20864 8928 20913 8956
rect 20864 8916 20870 8928
rect 20901 8925 20913 8928
rect 20947 8925 20959 8959
rect 25222 8956 25228 8968
rect 25183 8928 25228 8956
rect 20901 8919 20959 8925
rect 25222 8916 25228 8928
rect 25280 8916 25286 8968
rect 29917 8959 29975 8965
rect 29917 8925 29929 8959
rect 29963 8956 29975 8959
rect 30834 8956 30840 8968
rect 29963 8928 30840 8956
rect 29963 8925 29975 8928
rect 29917 8919 29975 8925
rect 30834 8916 30840 8928
rect 30892 8956 30898 8968
rect 31496 8965 31524 8996
rect 34790 8984 34796 9036
rect 34848 9024 34854 9036
rect 35437 9027 35495 9033
rect 35437 9024 35449 9027
rect 34848 8996 35449 9024
rect 34848 8984 34854 8996
rect 35437 8993 35449 8996
rect 35483 9024 35495 9027
rect 35894 9024 35900 9036
rect 35483 8996 35900 9024
rect 35483 8993 35495 8996
rect 35437 8987 35495 8993
rect 35894 8984 35900 8996
rect 35952 9024 35958 9036
rect 36354 9024 36360 9036
rect 35952 8996 36360 9024
rect 35952 8984 35958 8996
rect 31205 8959 31263 8965
rect 31205 8956 31217 8959
rect 30892 8928 31217 8956
rect 30892 8916 30898 8928
rect 31205 8925 31217 8928
rect 31251 8925 31263 8959
rect 31205 8919 31263 8925
rect 31481 8959 31539 8965
rect 31481 8925 31493 8959
rect 31527 8925 31539 8959
rect 31481 8919 31539 8925
rect 34698 8916 34704 8968
rect 34756 8956 34762 8968
rect 35158 8956 35164 8968
rect 34756 8928 35164 8956
rect 34756 8916 34762 8928
rect 35158 8916 35164 8928
rect 35216 8916 35222 8968
rect 35250 8916 35256 8968
rect 35308 8956 35314 8968
rect 36096 8965 36124 8996
rect 36354 8984 36360 8996
rect 36412 8984 36418 9036
rect 35345 8959 35403 8965
rect 35345 8956 35357 8959
rect 35308 8928 35357 8956
rect 35308 8916 35314 8928
rect 35345 8925 35357 8928
rect 35391 8925 35403 8959
rect 35345 8919 35403 8925
rect 36081 8959 36139 8965
rect 36081 8925 36093 8959
rect 36127 8925 36139 8959
rect 36081 8919 36139 8925
rect 2590 8888 2596 8900
rect 2551 8860 2596 8888
rect 2590 8848 2596 8860
rect 2648 8848 2654 8900
rect 2682 8848 2688 8900
rect 2740 8888 2746 8900
rect 2777 8891 2835 8897
rect 2777 8888 2789 8891
rect 2740 8860 2789 8888
rect 2740 8848 2746 8860
rect 2777 8857 2789 8860
rect 2823 8857 2835 8891
rect 2777 8851 2835 8857
rect 6365 8891 6423 8897
rect 6365 8857 6377 8891
rect 6411 8888 6423 8891
rect 6546 8888 6552 8900
rect 6411 8860 6552 8888
rect 6411 8857 6423 8860
rect 6365 8851 6423 8857
rect 6546 8848 6552 8860
rect 6604 8848 6610 8900
rect 20438 8848 20444 8900
rect 20496 8888 20502 8900
rect 20625 8891 20683 8897
rect 20625 8888 20637 8891
rect 20496 8860 20637 8888
rect 20496 8848 20502 8860
rect 20625 8857 20637 8860
rect 20671 8857 20683 8891
rect 20625 8851 20683 8857
rect 24026 8848 24032 8900
rect 24084 8888 24090 8900
rect 25409 8891 25467 8897
rect 25409 8888 25421 8891
rect 24084 8860 25421 8888
rect 24084 8848 24090 8860
rect 25409 8857 25421 8860
rect 25455 8857 25467 8891
rect 25409 8851 25467 8857
rect 29546 8848 29552 8900
rect 29604 8888 29610 8900
rect 30009 8891 30067 8897
rect 30009 8888 30021 8891
rect 29604 8860 30021 8888
rect 29604 8848 29610 8860
rect 30009 8857 30021 8860
rect 30055 8857 30067 8891
rect 30009 8851 30067 8857
rect 34606 8848 34612 8900
rect 34664 8888 34670 8900
rect 35268 8888 35296 8916
rect 34664 8860 35296 8888
rect 34664 8848 34670 8860
rect 5626 8780 5632 8832
rect 5684 8820 5690 8832
rect 5997 8823 6055 8829
rect 5997 8820 6009 8823
rect 5684 8792 6009 8820
rect 5684 8780 5690 8792
rect 5997 8789 6009 8792
rect 6043 8789 6055 8823
rect 5997 8783 6055 8789
rect 6457 8823 6515 8829
rect 6457 8789 6469 8823
rect 6503 8820 6515 8823
rect 6914 8820 6920 8832
rect 6503 8792 6920 8820
rect 6503 8789 6515 8792
rect 6457 8783 6515 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 11146 8820 11152 8832
rect 11107 8792 11152 8820
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 12069 8823 12127 8829
rect 12069 8789 12081 8823
rect 12115 8820 12127 8823
rect 12158 8820 12164 8832
rect 12115 8792 12164 8820
rect 12115 8789 12127 8792
rect 12069 8783 12127 8789
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 19705 8823 19763 8829
rect 19705 8820 19717 8823
rect 19484 8792 19717 8820
rect 19484 8780 19490 8792
rect 19705 8789 19717 8792
rect 19751 8789 19763 8823
rect 19705 8783 19763 8789
rect 21085 8823 21143 8829
rect 21085 8789 21097 8823
rect 21131 8820 21143 8823
rect 23750 8820 23756 8832
rect 21131 8792 23756 8820
rect 21131 8789 21143 8792
rect 21085 8783 21143 8789
rect 23750 8780 23756 8792
rect 23808 8780 23814 8832
rect 30374 8820 30380 8832
rect 30335 8792 30380 8820
rect 30374 8780 30380 8792
rect 30432 8780 30438 8832
rect 31662 8820 31668 8832
rect 31623 8792 31668 8820
rect 31662 8780 31668 8792
rect 31720 8780 31726 8832
rect 34514 8780 34520 8832
rect 34572 8820 34578 8832
rect 34977 8823 35035 8829
rect 34977 8820 34989 8823
rect 34572 8792 34989 8820
rect 34572 8780 34578 8792
rect 34977 8789 34989 8792
rect 35023 8789 35035 8823
rect 34977 8783 35035 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 5258 8616 5264 8628
rect 5219 8588 5264 8616
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5810 8616 5816 8628
rect 5736 8588 5816 8616
rect 5626 8548 5632 8560
rect 5587 8520 5632 8548
rect 5626 8508 5632 8520
rect 5684 8508 5690 8560
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 5445 8483 5503 8489
rect 5445 8480 5457 8483
rect 5408 8452 5457 8480
rect 5408 8440 5414 8452
rect 5445 8449 5457 8452
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5736 8480 5764 8588
rect 5810 8576 5816 8588
rect 5868 8616 5874 8628
rect 6365 8619 6423 8625
rect 6365 8616 6377 8619
rect 5868 8588 6377 8616
rect 5868 8576 5874 8588
rect 6365 8585 6377 8588
rect 6411 8585 6423 8619
rect 6914 8616 6920 8628
rect 6875 8588 6920 8616
rect 6365 8579 6423 8585
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 7285 8619 7343 8625
rect 7285 8585 7297 8619
rect 7331 8616 7343 8619
rect 9214 8616 9220 8628
rect 7331 8588 9220 8616
rect 7331 8585 7343 8588
rect 7285 8579 7343 8585
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 25130 8616 25136 8628
rect 13832 8588 25136 8616
rect 9309 8551 9367 8557
rect 9309 8517 9321 8551
rect 9355 8548 9367 8551
rect 11790 8548 11796 8560
rect 9355 8520 11796 8548
rect 9355 8517 9367 8520
rect 9309 8511 9367 8517
rect 11790 8508 11796 8520
rect 11848 8508 11854 8560
rect 12158 8548 12164 8560
rect 12119 8520 12164 8548
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 13722 8508 13728 8560
rect 13780 8548 13786 8560
rect 13832 8557 13860 8588
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 25222 8576 25228 8628
rect 25280 8616 25286 8628
rect 26050 8616 26056 8628
rect 25280 8588 26056 8616
rect 25280 8576 25286 8588
rect 26050 8576 26056 8588
rect 26108 8616 26114 8628
rect 28353 8619 28411 8625
rect 28353 8616 28365 8619
rect 26108 8588 28365 8616
rect 26108 8576 26114 8588
rect 28353 8585 28365 8588
rect 28399 8585 28411 8619
rect 28353 8579 28411 8585
rect 28626 8576 28632 8628
rect 28684 8616 28690 8628
rect 29825 8619 29883 8625
rect 29825 8616 29837 8619
rect 28684 8588 29837 8616
rect 28684 8576 28690 8588
rect 29825 8585 29837 8588
rect 29871 8585 29883 8619
rect 29825 8579 29883 8585
rect 34977 8619 35035 8625
rect 34977 8585 34989 8619
rect 35023 8616 35035 8619
rect 35342 8616 35348 8628
rect 35023 8588 35348 8616
rect 35023 8585 35035 8588
rect 34977 8579 35035 8585
rect 35342 8576 35348 8588
rect 35400 8576 35406 8628
rect 13817 8551 13875 8557
rect 13817 8548 13829 8551
rect 13780 8520 13829 8548
rect 13780 8508 13786 8520
rect 13817 8517 13829 8520
rect 13863 8517 13875 8551
rect 13817 8511 13875 8517
rect 16853 8551 16911 8557
rect 16853 8517 16865 8551
rect 16899 8548 16911 8551
rect 22094 8548 22100 8560
rect 16899 8520 22100 8548
rect 16899 8517 16911 8520
rect 16853 8511 16911 8517
rect 22094 8508 22100 8520
rect 22152 8508 22158 8560
rect 26988 8520 28856 8548
rect 5583 8452 5764 8480
rect 5813 8483 5871 8489
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 8294 8480 8300 8492
rect 5859 8452 8300 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 23750 8480 23756 8492
rect 23711 8452 23756 8480
rect 23750 8440 23756 8452
rect 23808 8440 23814 8492
rect 24026 8480 24032 8492
rect 23987 8452 24032 8480
rect 24026 8440 24032 8452
rect 24084 8440 24090 8492
rect 25133 8483 25191 8489
rect 25133 8480 25145 8483
rect 24872 8452 25145 8480
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 7374 8412 7380 8424
rect 5316 8384 7380 8412
rect 5316 8372 5322 8384
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 8754 8412 8760 8424
rect 8404 8384 8760 8412
rect 4062 8304 4068 8356
rect 4120 8344 4126 8356
rect 5166 8344 5172 8356
rect 4120 8316 5172 8344
rect 4120 8304 4126 8316
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 8404 8276 8432 8384
rect 8754 8372 8760 8384
rect 8812 8412 8818 8424
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 8812 8384 9137 8412
rect 8812 8372 8818 8384
rect 9125 8381 9137 8384
rect 9171 8381 9183 8415
rect 10962 8412 10968 8424
rect 10923 8384 10968 8412
rect 9125 8375 9183 8381
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 11974 8412 11980 8424
rect 11935 8384 11980 8412
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 16666 8344 16672 8356
rect 16627 8316 16672 8344
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 6696 8248 8432 8276
rect 6696 8236 6702 8248
rect 20714 8236 20720 8288
rect 20772 8276 20778 8288
rect 24872 8276 24900 8452
rect 25133 8449 25145 8452
rect 25179 8480 25191 8483
rect 25406 8480 25412 8492
rect 25179 8452 25412 8480
rect 25179 8449 25191 8452
rect 25133 8443 25191 8449
rect 25406 8440 25412 8452
rect 25464 8440 25470 8492
rect 25866 8480 25872 8492
rect 25827 8452 25872 8480
rect 25866 8440 25872 8452
rect 25924 8440 25930 8492
rect 25958 8440 25964 8492
rect 26016 8480 26022 8492
rect 26988 8489 27016 8520
rect 27246 8489 27252 8492
rect 26053 8483 26111 8489
rect 26053 8480 26065 8483
rect 26016 8452 26065 8480
rect 26016 8440 26022 8452
rect 26053 8449 26065 8452
rect 26099 8449 26111 8483
rect 26053 8443 26111 8449
rect 26973 8483 27031 8489
rect 26973 8449 26985 8483
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27240 8443 27252 8489
rect 27304 8480 27310 8492
rect 27304 8452 27340 8480
rect 27246 8440 27252 8443
rect 27304 8440 27310 8452
rect 28828 8356 28856 8520
rect 35158 8508 35164 8560
rect 35216 8548 35222 8560
rect 35526 8548 35532 8560
rect 35216 8520 35532 8548
rect 35216 8508 35222 8520
rect 35526 8508 35532 8520
rect 35584 8508 35590 8560
rect 35713 8551 35771 8557
rect 35713 8517 35725 8551
rect 35759 8548 35771 8551
rect 35894 8548 35900 8560
rect 35759 8520 35900 8548
rect 35759 8517 35771 8520
rect 35713 8511 35771 8517
rect 35894 8508 35900 8520
rect 35952 8508 35958 8560
rect 30009 8483 30067 8489
rect 30009 8449 30021 8483
rect 30055 8480 30067 8483
rect 30374 8480 30380 8492
rect 30055 8452 30380 8480
rect 30055 8449 30067 8452
rect 30009 8443 30067 8449
rect 30374 8440 30380 8452
rect 30432 8440 30438 8492
rect 30837 8483 30895 8489
rect 30837 8449 30849 8483
rect 30883 8480 30895 8483
rect 30926 8480 30932 8492
rect 30883 8452 30932 8480
rect 30883 8449 30895 8452
rect 30837 8443 30895 8449
rect 30926 8440 30932 8452
rect 30984 8480 30990 8492
rect 31297 8483 31355 8489
rect 31297 8480 31309 8483
rect 30984 8452 31309 8480
rect 30984 8440 30990 8452
rect 31297 8449 31309 8452
rect 31343 8449 31355 8483
rect 34514 8480 34520 8492
rect 34475 8452 34520 8480
rect 31297 8443 31355 8449
rect 34514 8440 34520 8452
rect 34572 8440 34578 8492
rect 34793 8483 34851 8489
rect 34793 8449 34805 8483
rect 34839 8449 34851 8483
rect 34793 8443 34851 8449
rect 30193 8415 30251 8421
rect 30193 8381 30205 8415
rect 30239 8412 30251 8415
rect 30466 8412 30472 8424
rect 30239 8384 30472 8412
rect 30239 8381 30251 8384
rect 30193 8375 30251 8381
rect 30466 8372 30472 8384
rect 30524 8372 30530 8424
rect 33502 8372 33508 8424
rect 33560 8412 33566 8424
rect 34146 8412 34152 8424
rect 33560 8384 34152 8412
rect 33560 8372 33566 8384
rect 34146 8372 34152 8384
rect 34204 8412 34210 8424
rect 34609 8415 34667 8421
rect 34609 8412 34621 8415
rect 34204 8384 34621 8412
rect 34204 8372 34210 8384
rect 34609 8381 34621 8384
rect 34655 8381 34667 8415
rect 34609 8375 34667 8381
rect 34808 8412 34836 8443
rect 35342 8440 35348 8492
rect 35400 8480 35406 8492
rect 35437 8483 35495 8489
rect 35437 8480 35449 8483
rect 35400 8452 35449 8480
rect 35400 8440 35406 8452
rect 35437 8449 35449 8452
rect 35483 8449 35495 8483
rect 35437 8443 35495 8449
rect 34808 8384 35480 8412
rect 25038 8304 25044 8356
rect 25096 8344 25102 8356
rect 25317 8347 25375 8353
rect 25317 8344 25329 8347
rect 25096 8316 25329 8344
rect 25096 8304 25102 8316
rect 25317 8313 25329 8316
rect 25363 8313 25375 8347
rect 28810 8344 28816 8356
rect 28771 8316 28816 8344
rect 25317 8307 25375 8313
rect 28810 8304 28816 8316
rect 28868 8344 28874 8356
rect 29362 8344 29368 8356
rect 28868 8316 29368 8344
rect 28868 8304 28874 8316
rect 29362 8304 29368 8316
rect 29420 8304 29426 8356
rect 33594 8304 33600 8356
rect 33652 8344 33658 8356
rect 34057 8347 34115 8353
rect 34057 8344 34069 8347
rect 33652 8316 34069 8344
rect 33652 8304 33658 8316
rect 34057 8313 34069 8316
rect 34103 8344 34115 8347
rect 34808 8344 34836 8384
rect 35452 8356 35480 8384
rect 34103 8316 34836 8344
rect 34103 8313 34115 8316
rect 34057 8307 34115 8313
rect 35434 8304 35440 8356
rect 35492 8304 35498 8356
rect 35710 8344 35716 8356
rect 35671 8316 35716 8344
rect 35710 8304 35716 8316
rect 35768 8304 35774 8356
rect 20772 8248 24900 8276
rect 26237 8279 26295 8285
rect 20772 8236 20778 8248
rect 26237 8245 26249 8279
rect 26283 8276 26295 8279
rect 26970 8276 26976 8288
rect 26283 8248 26976 8276
rect 26283 8245 26295 8248
rect 26237 8239 26295 8245
rect 26970 8236 26976 8248
rect 27028 8236 27034 8288
rect 30742 8276 30748 8288
rect 30703 8248 30748 8276
rect 30742 8236 30748 8248
rect 30800 8236 30806 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 2222 8072 2228 8084
rect 1627 8044 2228 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 19334 8032 19340 8084
rect 19392 8072 19398 8084
rect 28166 8072 28172 8084
rect 19392 8044 28172 8072
rect 19392 8032 19398 8044
rect 3510 7964 3516 8016
rect 3568 8004 3574 8016
rect 3568 7976 11468 8004
rect 3568 7964 3574 7976
rect 11440 7948 11468 7976
rect 19426 7964 19432 8016
rect 19484 8004 19490 8016
rect 19484 7976 19564 8004
rect 19484 7964 19490 7976
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 6638 7936 6644 7948
rect 5868 7908 6644 7936
rect 5868 7896 5874 7908
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 6825 7939 6883 7945
rect 6825 7905 6837 7939
rect 6871 7936 6883 7939
rect 7558 7936 7564 7948
rect 6871 7908 7564 7936
rect 6871 7905 6883 7908
rect 6825 7899 6883 7905
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 11146 7936 11152 7948
rect 11107 7908 11152 7936
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 11422 7936 11428 7948
rect 11335 7908 11428 7936
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 15286 7936 15292 7948
rect 15247 7908 15292 7936
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15746 7936 15752 7948
rect 15707 7908 15752 7936
rect 15746 7896 15752 7908
rect 15804 7896 15810 7948
rect 17126 7896 17132 7948
rect 17184 7936 17190 7948
rect 19536 7945 19564 7976
rect 19812 7945 19840 8044
rect 28166 8032 28172 8044
rect 28224 8032 28230 8084
rect 30377 8075 30435 8081
rect 30377 8041 30389 8075
rect 30423 8072 30435 8075
rect 30466 8072 30472 8084
rect 30423 8044 30472 8072
rect 30423 8041 30435 8044
rect 30377 8035 30435 8041
rect 30466 8032 30472 8044
rect 30524 8032 30530 8084
rect 35345 8075 35403 8081
rect 35345 8041 35357 8075
rect 35391 8072 35403 8075
rect 35526 8072 35532 8084
rect 35391 8044 35532 8072
rect 35391 8041 35403 8044
rect 35345 8035 35403 8041
rect 35526 8032 35532 8044
rect 35584 8032 35590 8084
rect 19337 7939 19395 7945
rect 19337 7936 19349 7939
rect 17184 7908 19349 7936
rect 17184 7896 17190 7908
rect 19337 7905 19349 7908
rect 19383 7905 19395 7939
rect 19337 7899 19395 7905
rect 19521 7939 19579 7945
rect 19521 7905 19533 7939
rect 19567 7905 19579 7939
rect 19521 7899 19579 7905
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7936 19855 7939
rect 19978 7936 19984 7948
rect 19843 7908 19984 7936
rect 19843 7905 19855 7908
rect 19797 7899 19855 7905
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7868 1458 7880
rect 2041 7871 2099 7877
rect 2041 7868 2053 7871
rect 1452 7840 2053 7868
rect 1452 7828 1458 7840
rect 2041 7837 2053 7840
rect 2087 7837 2099 7871
rect 6546 7868 6552 7880
rect 6507 7840 6552 7868
rect 2041 7831 2099 7837
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 10980 7800 11008 7831
rect 14550 7828 14556 7880
rect 14608 7868 14614 7880
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 14608 7840 15117 7868
rect 14608 7828 14614 7840
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7868 17739 7871
rect 18598 7868 18604 7880
rect 17727 7840 18604 7868
rect 17727 7837 17739 7840
rect 17681 7831 17739 7837
rect 16850 7800 16856 7812
rect 10100 7772 16856 7800
rect 10100 7760 10106 7772
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 6181 7735 6239 7741
rect 6181 7732 6193 7735
rect 5500 7704 6193 7732
rect 5500 7692 5506 7704
rect 6181 7701 6193 7704
rect 6227 7701 6239 7735
rect 6181 7695 6239 7701
rect 17865 7735 17923 7741
rect 17865 7701 17877 7735
rect 17911 7732 17923 7735
rect 18322 7732 18328 7744
rect 17911 7704 18328 7732
rect 17911 7701 17923 7704
rect 17865 7695 17923 7701
rect 18322 7692 18328 7704
rect 18380 7692 18386 7744
rect 18524 7741 18552 7840
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 19352 7800 19380 7899
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 21726 7896 21732 7948
rect 21784 7936 21790 7948
rect 22649 7939 22707 7945
rect 22649 7936 22661 7939
rect 21784 7908 22661 7936
rect 21784 7896 21790 7908
rect 22649 7905 22661 7908
rect 22695 7905 22707 7939
rect 25314 7936 25320 7948
rect 25275 7908 25320 7936
rect 22649 7899 22707 7905
rect 25314 7896 25320 7908
rect 25372 7896 25378 7948
rect 26602 7896 26608 7948
rect 26660 7936 26666 7948
rect 26973 7939 27031 7945
rect 26973 7936 26985 7939
rect 26660 7908 26985 7936
rect 26660 7896 26666 7908
rect 26973 7905 26985 7908
rect 27019 7905 27031 7939
rect 26973 7899 27031 7905
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7868 22983 7871
rect 25590 7868 25596 7880
rect 22971 7840 25596 7868
rect 22971 7837 22983 7840
rect 22925 7831 22983 7837
rect 25590 7828 25596 7840
rect 25648 7828 25654 7880
rect 27157 7871 27215 7877
rect 27157 7837 27169 7871
rect 27203 7868 27215 7871
rect 28718 7868 28724 7880
rect 27203 7840 28724 7868
rect 27203 7837 27215 7840
rect 27157 7831 27215 7837
rect 28718 7828 28724 7840
rect 28776 7828 28782 7880
rect 35158 7868 35164 7880
rect 35119 7840 35164 7868
rect 35158 7828 35164 7840
rect 35216 7828 35222 7880
rect 35342 7828 35348 7880
rect 35400 7868 35406 7880
rect 35618 7868 35624 7880
rect 35400 7840 35624 7868
rect 35400 7828 35406 7840
rect 35618 7828 35624 7840
rect 35676 7828 35682 7880
rect 20438 7800 20444 7812
rect 19352 7772 20444 7800
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 21266 7760 21272 7812
rect 21324 7800 21330 7812
rect 21821 7803 21879 7809
rect 21821 7800 21833 7803
rect 21324 7772 21833 7800
rect 21324 7760 21330 7772
rect 21821 7769 21833 7772
rect 21867 7769 21879 7803
rect 21821 7763 21879 7769
rect 22005 7803 22063 7809
rect 22005 7769 22017 7803
rect 22051 7800 22063 7803
rect 25958 7800 25964 7812
rect 22051 7772 25964 7800
rect 22051 7769 22063 7772
rect 22005 7763 22063 7769
rect 25958 7760 25964 7772
rect 26016 7760 26022 7812
rect 18509 7735 18567 7741
rect 18509 7701 18521 7735
rect 18555 7732 18567 7735
rect 20162 7732 20168 7744
rect 18555 7704 20168 7732
rect 18555 7701 18567 7704
rect 18509 7695 18567 7701
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 22189 7735 22247 7741
rect 22189 7701 22201 7735
rect 22235 7732 22247 7735
rect 22278 7732 22284 7744
rect 22235 7704 22284 7732
rect 22235 7701 22247 7704
rect 22189 7695 22247 7701
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 35529 7735 35587 7741
rect 35529 7701 35541 7735
rect 35575 7732 35587 7735
rect 35894 7732 35900 7744
rect 35575 7704 35900 7732
rect 35575 7701 35587 7704
rect 35529 7695 35587 7701
rect 35894 7692 35900 7704
rect 35952 7692 35958 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 5442 7528 5448 7540
rect 5403 7500 5448 7528
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 10042 7528 10048 7540
rect 10003 7500 10048 7528
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10192 7500 10237 7528
rect 10192 7488 10198 7500
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 19334 7528 19340 7540
rect 11480 7500 19340 7528
rect 11480 7488 11486 7500
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 19978 7528 19984 7540
rect 19939 7500 19984 7528
rect 19978 7488 19984 7500
rect 20036 7528 20042 7540
rect 20901 7531 20959 7537
rect 20901 7528 20913 7531
rect 20036 7500 20913 7528
rect 20036 7488 20042 7500
rect 20901 7497 20913 7500
rect 20947 7497 20959 7531
rect 21266 7528 21272 7540
rect 21227 7500 21272 7528
rect 20901 7491 20959 7497
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 23106 7488 23112 7540
rect 23164 7528 23170 7540
rect 23937 7531 23995 7537
rect 23937 7528 23949 7531
rect 23164 7500 23949 7528
rect 23164 7488 23170 7500
rect 23937 7497 23949 7500
rect 23983 7528 23995 7531
rect 24394 7528 24400 7540
rect 23983 7500 24400 7528
rect 23983 7497 23995 7500
rect 23937 7491 23995 7497
rect 24394 7488 24400 7500
rect 24452 7488 24458 7540
rect 25593 7531 25651 7537
rect 25593 7497 25605 7531
rect 25639 7528 25651 7531
rect 25866 7528 25872 7540
rect 25639 7500 25872 7528
rect 25639 7497 25651 7500
rect 25593 7491 25651 7497
rect 25866 7488 25872 7500
rect 25924 7488 25930 7540
rect 26050 7528 26056 7540
rect 26011 7500 26056 7528
rect 26050 7488 26056 7500
rect 26108 7528 26114 7540
rect 27157 7531 27215 7537
rect 26108 7500 26234 7528
rect 26108 7488 26114 7500
rect 12618 7460 12624 7472
rect 12579 7432 12624 7460
rect 12618 7420 12624 7432
rect 12676 7420 12682 7472
rect 14182 7420 14188 7472
rect 14240 7460 14246 7472
rect 14277 7463 14335 7469
rect 14277 7460 14289 7463
rect 14240 7432 14289 7460
rect 14240 7420 14246 7432
rect 14277 7429 14289 7432
rect 14323 7460 14335 7463
rect 25961 7463 26019 7469
rect 25961 7460 25973 7463
rect 14323 7432 25973 7460
rect 14323 7429 14335 7432
rect 14277 7423 14335 7429
rect 25961 7429 25973 7432
rect 26007 7429 26019 7463
rect 26206 7460 26234 7500
rect 27157 7497 27169 7531
rect 27203 7528 27215 7531
rect 27246 7528 27252 7540
rect 27203 7500 27252 7528
rect 27203 7497 27215 7500
rect 27157 7491 27215 7497
rect 27246 7488 27252 7500
rect 27304 7488 27310 7540
rect 30653 7531 30711 7537
rect 27356 7500 30236 7528
rect 27356 7460 27384 7500
rect 26206 7432 27384 7460
rect 25961 7423 26019 7429
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 5316 7364 5365 7392
rect 5316 7352 5322 7364
rect 5353 7361 5365 7364
rect 5399 7392 5411 7395
rect 5442 7392 5448 7404
rect 5399 7364 5448 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 15286 7392 15292 7404
rect 15247 7364 15292 7392
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7392 15439 7395
rect 15562 7392 15568 7404
rect 15427 7364 15568 7392
rect 15427 7361 15439 7364
rect 15381 7355 15439 7361
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 17126 7352 17132 7404
rect 17184 7392 17190 7404
rect 17221 7395 17279 7401
rect 17221 7392 17233 7395
rect 17184 7364 17233 7392
rect 17184 7352 17190 7364
rect 17221 7361 17233 7364
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 20622 7352 20628 7404
rect 20680 7392 20686 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20680 7364 20821 7392
rect 20680 7352 20686 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 21542 7352 21548 7404
rect 21600 7392 21606 7404
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 21600 7364 21833 7392
rect 21600 7352 21606 7364
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 23106 7392 23112 7404
rect 23067 7364 23112 7392
rect 21821 7355 21879 7361
rect 23106 7352 23112 7364
rect 23164 7352 23170 7404
rect 25976 7392 26004 7423
rect 27522 7420 27528 7472
rect 27580 7460 27586 7472
rect 27985 7463 28043 7469
rect 27985 7460 27997 7463
rect 27580 7432 27997 7460
rect 27580 7420 27586 7432
rect 27985 7429 27997 7432
rect 28031 7429 28043 7463
rect 27985 7423 28043 7429
rect 29178 7420 29184 7472
rect 29236 7460 29242 7472
rect 29638 7460 29644 7472
rect 29236 7432 29644 7460
rect 29236 7420 29242 7432
rect 29638 7420 29644 7432
rect 29696 7420 29702 7472
rect 26602 7392 26608 7404
rect 25976 7364 26608 7392
rect 26602 7352 26608 7364
rect 26660 7392 26666 7404
rect 26970 7392 26976 7404
rect 26660 7364 26740 7392
rect 26931 7364 26976 7392
rect 26660 7352 26666 7364
rect 5626 7324 5632 7336
rect 5587 7296 5632 7324
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 10321 7327 10379 7333
rect 10321 7293 10333 7327
rect 10367 7293 10379 7327
rect 10321 7287 10379 7293
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 10336 7256 10364 7287
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 15473 7327 15531 7333
rect 12492 7296 12537 7324
rect 12492 7284 12498 7296
rect 15473 7293 15485 7327
rect 15519 7293 15531 7327
rect 20714 7324 20720 7336
rect 20675 7296 20720 7324
rect 15473 7287 15531 7293
rect 15488 7256 15516 7287
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 22094 7324 22100 7336
rect 22055 7296 22100 7324
rect 22094 7284 22100 7296
rect 22152 7284 22158 7336
rect 15562 7256 15568 7268
rect 7616 7228 15568 7256
rect 7616 7216 7622 7228
rect 15562 7216 15568 7228
rect 15620 7256 15626 7268
rect 17037 7259 17095 7265
rect 17037 7256 17049 7259
rect 15620 7228 17049 7256
rect 15620 7216 15626 7228
rect 17037 7225 17049 7228
rect 17083 7225 17095 7259
rect 17037 7219 17095 7225
rect 19334 7216 19340 7268
rect 19392 7256 19398 7268
rect 23124 7256 23152 7352
rect 25406 7284 25412 7336
rect 25464 7324 25470 7336
rect 26145 7327 26203 7333
rect 26145 7324 26157 7327
rect 25464 7296 26157 7324
rect 25464 7284 25470 7296
rect 26145 7293 26157 7296
rect 26191 7293 26203 7327
rect 26712 7324 26740 7364
rect 26970 7352 26976 7364
rect 27028 7352 27034 7404
rect 29270 7352 29276 7404
rect 29328 7392 29334 7404
rect 30208 7401 30236 7500
rect 30653 7497 30665 7531
rect 30699 7528 30711 7531
rect 35158 7528 35164 7540
rect 30699 7500 35164 7528
rect 30699 7497 30711 7500
rect 30653 7491 30711 7497
rect 35158 7488 35164 7500
rect 35216 7488 35222 7540
rect 33594 7460 33600 7472
rect 33555 7432 33600 7460
rect 33594 7420 33600 7432
rect 33652 7420 33658 7472
rect 30101 7395 30159 7401
rect 30101 7392 30113 7395
rect 29328 7364 30113 7392
rect 29328 7352 29334 7364
rect 30101 7361 30113 7364
rect 30147 7361 30159 7395
rect 30101 7355 30159 7361
rect 30193 7395 30251 7401
rect 30193 7361 30205 7395
rect 30239 7361 30251 7395
rect 30374 7392 30380 7404
rect 30335 7364 30380 7392
rect 30193 7355 30251 7361
rect 30374 7352 30380 7364
rect 30432 7352 30438 7404
rect 30466 7352 30472 7404
rect 30524 7392 30530 7404
rect 30524 7364 30569 7392
rect 30524 7352 30530 7364
rect 30742 7352 30748 7404
rect 30800 7392 30806 7404
rect 32125 7395 32183 7401
rect 32125 7392 32137 7395
rect 30800 7364 32137 7392
rect 30800 7352 30806 7364
rect 32125 7361 32137 7364
rect 32171 7361 32183 7395
rect 32125 7355 32183 7361
rect 27062 7324 27068 7336
rect 26712 7296 27068 7324
rect 26145 7287 26203 7293
rect 27062 7284 27068 7296
rect 27120 7284 27126 7336
rect 27801 7327 27859 7333
rect 27801 7293 27813 7327
rect 27847 7324 27859 7327
rect 28074 7324 28080 7336
rect 27847 7296 28080 7324
rect 27847 7293 27859 7296
rect 27801 7287 27859 7293
rect 28074 7284 28080 7296
rect 28132 7284 28138 7336
rect 19392 7228 23152 7256
rect 32309 7259 32367 7265
rect 19392 7216 19398 7228
rect 32309 7225 32321 7259
rect 32355 7256 32367 7259
rect 33594 7256 33600 7268
rect 32355 7228 33600 7256
rect 32355 7225 32367 7228
rect 32309 7219 32367 7225
rect 33594 7216 33600 7228
rect 33652 7216 33658 7268
rect 4798 7148 4804 7200
rect 4856 7188 4862 7200
rect 4985 7191 5043 7197
rect 4985 7188 4997 7191
rect 4856 7160 4997 7188
rect 4856 7148 4862 7160
rect 4985 7157 4997 7160
rect 5031 7157 5043 7191
rect 9674 7188 9680 7200
rect 9635 7160 9680 7188
rect 4985 7151 5043 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 14918 7188 14924 7200
rect 14879 7160 14924 7188
rect 14918 7148 14924 7160
rect 14976 7148 14982 7200
rect 23290 7188 23296 7200
rect 23251 7160 23296 7188
rect 23290 7148 23296 7160
rect 23348 7148 23354 7200
rect 28626 7148 28632 7200
rect 28684 7188 28690 7200
rect 29546 7188 29552 7200
rect 28684 7160 29552 7188
rect 28684 7148 28690 7160
rect 29546 7148 29552 7160
rect 29604 7148 29610 7200
rect 36170 7188 36176 7200
rect 36131 7160 36176 7188
rect 36170 7148 36176 7160
rect 36228 7148 36234 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 23290 6944 23296 6996
rect 23348 6984 23354 6996
rect 28626 6984 28632 6996
rect 23348 6956 28632 6984
rect 23348 6944 23354 6956
rect 28626 6944 28632 6956
rect 28684 6944 28690 6996
rect 28905 6987 28963 6993
rect 28905 6953 28917 6987
rect 28951 6984 28963 6987
rect 30466 6984 30472 6996
rect 28951 6956 30472 6984
rect 28951 6953 28963 6956
rect 28905 6947 28963 6953
rect 30466 6944 30472 6956
rect 30524 6944 30530 6996
rect 30558 6944 30564 6996
rect 30616 6984 30622 6996
rect 30616 6956 30661 6984
rect 30616 6944 30622 6956
rect 28074 6876 28080 6928
rect 28132 6916 28138 6928
rect 29270 6916 29276 6928
rect 28132 6888 29276 6916
rect 28132 6876 28138 6888
rect 29270 6876 29276 6888
rect 29328 6876 29334 6928
rect 30374 6876 30380 6928
rect 30432 6876 30438 6928
rect 33980 6888 34284 6916
rect 5166 6848 5172 6860
rect 5127 6820 5172 6848
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 9585 6851 9643 6857
rect 7944 6820 8432 6848
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6780 1458 6792
rect 2041 6783 2099 6789
rect 2041 6780 2053 6783
rect 1452 6752 2053 6780
rect 1452 6740 1458 6752
rect 2041 6749 2053 6752
rect 2087 6749 2099 6783
rect 3970 6780 3976 6792
rect 3931 6752 3976 6780
rect 2041 6743 2099 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4172 6712 4200 6743
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 5350 6780 5356 6792
rect 4672 6752 5356 6780
rect 4672 6740 4678 6752
rect 5350 6740 5356 6752
rect 5408 6780 5414 6792
rect 7944 6789 7972 6820
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 5408 6752 7941 6780
rect 5408 6740 5414 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8018 6740 8024 6792
rect 8076 6780 8082 6792
rect 8294 6780 8300 6792
rect 8076 6752 8121 6780
rect 8255 6752 8300 6780
rect 8076 6740 8082 6752
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8113 6715 8171 6721
rect 4172 6684 4752 6712
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2682 6644 2688 6656
rect 1627 6616 2688 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 2866 6604 2872 6656
rect 2924 6644 2930 6656
rect 4724 6653 4752 6684
rect 8113 6681 8125 6715
rect 8159 6681 8171 6715
rect 8404 6712 8432 6820
rect 9585 6817 9597 6851
rect 9631 6848 9643 6851
rect 10226 6848 10232 6860
rect 9631 6820 10232 6848
rect 9631 6817 9643 6820
rect 9585 6811 9643 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 15562 6848 15568 6860
rect 15523 6820 15568 6848
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 16482 6808 16488 6860
rect 16540 6848 16546 6860
rect 16761 6851 16819 6857
rect 16761 6848 16773 6851
rect 16540 6820 16773 6848
rect 16540 6808 16546 6820
rect 16761 6817 16773 6820
rect 16807 6817 16819 6851
rect 26602 6848 26608 6860
rect 16761 6811 16819 6817
rect 18156 6820 19380 6848
rect 26563 6820 26608 6848
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 9674 6780 9680 6792
rect 9447 6752 9680 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 15654 6740 15660 6792
rect 15712 6780 15718 6792
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15712 6752 15853 6780
rect 15712 6740 15718 6752
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 16850 6740 16856 6792
rect 16908 6780 16914 6792
rect 17037 6783 17095 6789
rect 17037 6780 17049 6783
rect 16908 6752 17049 6780
rect 16908 6740 16914 6752
rect 17037 6749 17049 6752
rect 17083 6749 17095 6783
rect 17037 6743 17095 6749
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 18156 6789 18184 6820
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 17276 6752 18061 6780
rect 17276 6740 17282 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6749 18199 6783
rect 18414 6780 18420 6792
rect 18375 6752 18420 6780
rect 18141 6743 18199 6749
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 19352 6789 19380 6820
rect 26602 6808 26608 6820
rect 26660 6808 26666 6860
rect 29917 6851 29975 6857
rect 29917 6817 29929 6851
rect 29963 6848 29975 6851
rect 30392 6848 30420 6876
rect 29963 6820 30420 6848
rect 29963 6817 29975 6820
rect 29917 6811 29975 6817
rect 33318 6808 33324 6860
rect 33376 6848 33382 6860
rect 33980 6848 34008 6888
rect 34146 6848 34152 6860
rect 33376 6820 34008 6848
rect 34107 6820 34152 6848
rect 33376 6808 33382 6820
rect 34146 6808 34152 6820
rect 34204 6808 34210 6860
rect 19337 6783 19395 6789
rect 19337 6749 19349 6783
rect 19383 6780 19395 6783
rect 22186 6780 22192 6792
rect 19383 6752 22094 6780
rect 22147 6752 22192 6780
rect 19383 6749 19395 6752
rect 19337 6743 19395 6749
rect 17236 6712 17264 6740
rect 18233 6715 18291 6721
rect 8404 6684 17264 6712
rect 17420 6684 18092 6712
rect 8113 6675 8171 6681
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 2924 6616 3801 6644
rect 2924 6604 2930 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 3789 6607 3847 6613
rect 4709 6647 4767 6653
rect 4709 6613 4721 6647
rect 4755 6644 4767 6647
rect 4890 6644 4896 6656
rect 4755 6616 4896 6644
rect 4755 6613 4767 6616
rect 4709 6607 4767 6613
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 5721 6647 5779 6653
rect 5721 6644 5733 6647
rect 5592 6616 5733 6644
rect 5592 6604 5598 6616
rect 5721 6613 5733 6616
rect 5767 6613 5779 6647
rect 5721 6607 5779 6613
rect 7745 6647 7803 6653
rect 7745 6613 7757 6647
rect 7791 6644 7803 6647
rect 7926 6644 7932 6656
rect 7791 6616 7932 6644
rect 7791 6613 7803 6616
rect 7745 6607 7803 6613
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8128 6644 8156 6675
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8128 6616 8953 6644
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 9306 6644 9312 6656
rect 9267 6616 9312 6644
rect 8941 6607 8999 6613
rect 9306 6604 9312 6616
rect 9364 6644 9370 6656
rect 11974 6644 11980 6656
rect 9364 6616 11980 6644
rect 9364 6604 9370 6616
rect 11974 6604 11980 6616
rect 12032 6644 12038 6656
rect 15378 6644 15384 6656
rect 12032 6616 15384 6644
rect 12032 6604 12038 6616
rect 15378 6604 15384 6616
rect 15436 6644 15442 6656
rect 17420 6653 17448 6684
rect 15749 6647 15807 6653
rect 15749 6644 15761 6647
rect 15436 6616 15761 6644
rect 15436 6604 15442 6616
rect 15749 6613 15761 6616
rect 15795 6613 15807 6647
rect 15749 6607 15807 6613
rect 16209 6647 16267 6653
rect 16209 6613 16221 6647
rect 16255 6644 16267 6647
rect 16945 6647 17003 6653
rect 16945 6644 16957 6647
rect 16255 6616 16957 6644
rect 16255 6613 16267 6616
rect 16209 6607 16267 6613
rect 16945 6613 16957 6616
rect 16991 6613 17003 6647
rect 16945 6607 17003 6613
rect 17405 6647 17463 6653
rect 17405 6613 17417 6647
rect 17451 6613 17463 6647
rect 17862 6644 17868 6656
rect 17823 6616 17868 6644
rect 17405 6607 17463 6613
rect 17862 6604 17868 6616
rect 17920 6604 17926 6656
rect 18064 6644 18092 6684
rect 18233 6681 18245 6715
rect 18279 6681 18291 6715
rect 20162 6712 20168 6724
rect 20075 6684 20168 6712
rect 18233 6675 18291 6681
rect 18248 6644 18276 6675
rect 20162 6672 20168 6684
rect 20220 6712 20226 6724
rect 20714 6712 20720 6724
rect 20220 6684 20720 6712
rect 20220 6672 20226 6684
rect 20714 6672 20720 6684
rect 20772 6672 20778 6724
rect 21818 6672 21824 6724
rect 21876 6712 21882 6724
rect 21922 6715 21980 6721
rect 21922 6712 21934 6715
rect 21876 6684 21934 6712
rect 21876 6672 21882 6684
rect 21922 6681 21934 6684
rect 21968 6681 21980 6715
rect 22066 6712 22094 6752
rect 22186 6740 22192 6752
rect 22244 6740 22250 6792
rect 26142 6780 26148 6792
rect 26103 6752 26148 6780
rect 26142 6740 26148 6752
rect 26200 6740 26206 6792
rect 27706 6740 27712 6792
rect 27764 6780 27770 6792
rect 28718 6780 28724 6792
rect 27764 6752 28724 6780
rect 27764 6740 27770 6752
rect 28718 6740 28724 6752
rect 28776 6780 28782 6792
rect 28813 6783 28871 6789
rect 28813 6780 28825 6783
rect 28776 6752 28825 6780
rect 28776 6740 28782 6752
rect 28813 6749 28825 6752
rect 28859 6749 28871 6783
rect 28813 6743 28871 6749
rect 28997 6783 29055 6789
rect 28997 6749 29009 6783
rect 29043 6780 29055 6783
rect 29733 6783 29791 6789
rect 29733 6780 29745 6783
rect 29043 6752 29745 6780
rect 29043 6749 29055 6752
rect 28997 6743 29055 6749
rect 29733 6749 29745 6752
rect 29779 6749 29791 6783
rect 30374 6780 30380 6792
rect 30287 6752 30380 6780
rect 29733 6743 29791 6749
rect 23290 6712 23296 6724
rect 22066 6684 23296 6712
rect 21922 6675 21980 6681
rect 23290 6672 23296 6684
rect 23348 6672 23354 6724
rect 28828 6712 28856 6743
rect 29549 6715 29607 6721
rect 29549 6712 29561 6715
rect 28828 6684 29561 6712
rect 29549 6681 29561 6684
rect 29595 6681 29607 6715
rect 29748 6712 29776 6743
rect 30374 6740 30380 6752
rect 30432 6780 30438 6792
rect 30742 6780 30748 6792
rect 30432 6752 30748 6780
rect 30432 6740 30438 6752
rect 30742 6740 30748 6752
rect 30800 6740 30806 6792
rect 31389 6783 31447 6789
rect 31389 6749 31401 6783
rect 31435 6780 31447 6783
rect 31754 6780 31760 6792
rect 31435 6752 31760 6780
rect 31435 6749 31447 6752
rect 31389 6743 31447 6749
rect 31754 6740 31760 6752
rect 31812 6780 31818 6792
rect 33229 6783 33287 6789
rect 33229 6780 33241 6783
rect 31812 6752 33241 6780
rect 31812 6740 31818 6752
rect 33229 6749 33241 6752
rect 33275 6749 33287 6783
rect 33229 6743 33287 6749
rect 32858 6712 32864 6724
rect 29748 6684 32864 6712
rect 29549 6675 29607 6681
rect 32858 6672 32864 6684
rect 32916 6672 32922 6724
rect 32984 6715 33042 6721
rect 32984 6681 32996 6715
rect 33030 6712 33042 6715
rect 33244 6712 33272 6743
rect 33594 6740 33600 6792
rect 33652 6780 33658 6792
rect 33873 6783 33931 6789
rect 33873 6780 33885 6783
rect 33652 6752 33885 6780
rect 33652 6740 33658 6752
rect 33873 6749 33885 6752
rect 33919 6749 33931 6783
rect 34054 6780 34060 6792
rect 34015 6752 34060 6780
rect 33873 6743 33931 6749
rect 34054 6740 34060 6752
rect 34112 6740 34118 6792
rect 34256 6780 34284 6888
rect 35710 6848 35716 6860
rect 35671 6820 35716 6848
rect 35710 6808 35716 6820
rect 35768 6808 35774 6860
rect 35894 6848 35900 6860
rect 35855 6820 35900 6848
rect 35894 6808 35900 6820
rect 35952 6808 35958 6860
rect 36004 6820 36492 6848
rect 35618 6780 35624 6792
rect 34256 6752 35624 6780
rect 35618 6740 35624 6752
rect 35676 6780 35682 6792
rect 36004 6780 36032 6820
rect 35676 6752 36032 6780
rect 36357 6783 36415 6789
rect 35676 6740 35682 6752
rect 36357 6749 36369 6783
rect 36403 6749 36415 6783
rect 36464 6780 36492 6820
rect 36464 6752 36768 6780
rect 36357 6743 36415 6749
rect 36170 6712 36176 6724
rect 33030 6684 33180 6712
rect 33244 6684 36176 6712
rect 33030 6681 33042 6684
rect 32984 6675 33042 6681
rect 20070 6644 20076 6656
rect 18064 6616 18276 6644
rect 20031 6616 20076 6644
rect 20070 6604 20076 6616
rect 20128 6604 20134 6656
rect 20438 6604 20444 6656
rect 20496 6644 20502 6656
rect 20809 6647 20867 6653
rect 20809 6644 20821 6647
rect 20496 6616 20821 6644
rect 20496 6604 20502 6616
rect 20809 6613 20821 6616
rect 20855 6613 20867 6647
rect 25958 6644 25964 6656
rect 25919 6616 25964 6644
rect 20809 6607 20867 6613
rect 25958 6604 25964 6616
rect 26016 6604 26022 6656
rect 31849 6647 31907 6653
rect 31849 6613 31861 6647
rect 31895 6644 31907 6647
rect 32214 6644 32220 6656
rect 31895 6616 32220 6644
rect 31895 6613 31907 6616
rect 31849 6607 31907 6613
rect 32214 6604 32220 6616
rect 32272 6604 32278 6656
rect 33152 6644 33180 6684
rect 36170 6672 36176 6684
rect 36228 6712 36234 6724
rect 36372 6712 36400 6743
rect 36228 6684 36400 6712
rect 36228 6672 36234 6684
rect 36446 6672 36452 6724
rect 36504 6712 36510 6724
rect 36602 6715 36660 6721
rect 36602 6712 36614 6715
rect 36504 6684 36614 6712
rect 36504 6672 36510 6684
rect 36602 6681 36614 6684
rect 36648 6681 36660 6715
rect 36602 6675 36660 6681
rect 33689 6647 33747 6653
rect 33689 6644 33701 6647
rect 33152 6616 33701 6644
rect 33689 6613 33701 6616
rect 33735 6613 33747 6647
rect 33689 6607 33747 6613
rect 35897 6647 35955 6653
rect 35897 6613 35909 6647
rect 35943 6644 35955 6647
rect 35986 6644 35992 6656
rect 35943 6616 35992 6644
rect 35943 6613 35955 6616
rect 35897 6607 35955 6613
rect 35986 6604 35992 6616
rect 36044 6604 36050 6656
rect 36740 6644 36768 6752
rect 37737 6647 37795 6653
rect 37737 6644 37749 6647
rect 36740 6616 37749 6644
rect 37737 6613 37749 6616
rect 37783 6613 37795 6647
rect 37737 6607 37795 6613
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 3605 6443 3663 6449
rect 3605 6409 3617 6443
rect 3651 6440 3663 6443
rect 5810 6440 5816 6452
rect 3651 6412 5816 6440
rect 3651 6409 3663 6412
rect 3605 6403 3663 6409
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8389 6443 8447 6449
rect 8389 6440 8401 6443
rect 8076 6412 8401 6440
rect 8076 6400 8082 6412
rect 8389 6409 8401 6412
rect 8435 6440 8447 6443
rect 13722 6440 13728 6452
rect 8435 6412 13728 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 14550 6440 14556 6452
rect 14511 6412 14556 6440
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 14645 6443 14703 6449
rect 14645 6409 14657 6443
rect 14691 6440 14703 6443
rect 14918 6440 14924 6452
rect 14691 6412 14924 6440
rect 14691 6409 14703 6412
rect 14645 6403 14703 6409
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 15749 6443 15807 6449
rect 15749 6440 15761 6443
rect 15712 6412 15761 6440
rect 15712 6400 15718 6412
rect 15749 6409 15761 6412
rect 15795 6409 15807 6443
rect 21818 6440 21824 6452
rect 21779 6412 21824 6440
rect 15749 6403 15807 6409
rect 21818 6400 21824 6412
rect 21876 6400 21882 6452
rect 33413 6443 33471 6449
rect 22066 6412 26234 6440
rect 3878 6372 3884 6384
rect 2240 6344 3884 6372
rect 2240 6313 2268 6344
rect 3878 6332 3884 6344
rect 3936 6332 3942 6384
rect 4798 6372 4804 6384
rect 4759 6344 4804 6372
rect 4798 6332 4804 6344
rect 4856 6332 4862 6384
rect 5166 6372 5172 6384
rect 4908 6344 5172 6372
rect 2498 6313 2504 6316
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2492 6267 2504 6313
rect 2556 6304 2562 6316
rect 4614 6304 4620 6316
rect 2556 6276 2592 6304
rect 4575 6276 4620 6304
rect 2498 6264 2504 6267
rect 2556 6264 2562 6276
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6304 4767 6307
rect 4908 6304 4936 6344
rect 5166 6332 5172 6344
rect 5224 6332 5230 6384
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 14366 6372 14372 6384
rect 8352 6344 14372 6372
rect 8352 6332 8358 6344
rect 14366 6332 14372 6344
rect 14424 6372 14430 6384
rect 18414 6372 18420 6384
rect 14424 6344 18420 6372
rect 14424 6332 14430 6344
rect 18414 6332 18420 6344
rect 18472 6332 18478 6384
rect 20070 6332 20076 6384
rect 20128 6372 20134 6384
rect 22066 6372 22094 6412
rect 25590 6372 25596 6384
rect 20128 6344 22094 6372
rect 25551 6344 25596 6372
rect 20128 6332 20134 6344
rect 25590 6332 25596 6344
rect 25648 6332 25654 6384
rect 26206 6372 26234 6412
rect 33413 6409 33425 6443
rect 33459 6440 33471 6443
rect 34054 6440 34060 6452
rect 33459 6412 34060 6440
rect 33459 6409 33471 6412
rect 33413 6403 33471 6409
rect 34054 6400 34060 6412
rect 34112 6400 34118 6452
rect 35618 6400 35624 6452
rect 35676 6440 35682 6452
rect 36446 6440 36452 6452
rect 35676 6412 36216 6440
rect 36407 6412 36452 6440
rect 35676 6400 35682 6412
rect 33965 6375 34023 6381
rect 33965 6372 33977 6375
rect 26206 6344 33977 6372
rect 4755 6276 4936 6304
rect 4985 6307 5043 6313
rect 4755 6273 4767 6276
rect 4709 6267 4767 6273
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5534 6304 5540 6316
rect 5031 6276 5540 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 17218 6304 17224 6316
rect 17179 6276 17224 6304
rect 17218 6264 17224 6276
rect 17276 6264 17282 6316
rect 22005 6307 22063 6313
rect 22005 6273 22017 6307
rect 22051 6304 22063 6307
rect 22278 6304 22284 6316
rect 22051 6276 22284 6304
rect 22051 6273 22063 6276
rect 22005 6267 22063 6273
rect 22278 6264 22284 6276
rect 22336 6264 22342 6316
rect 23934 6304 23940 6316
rect 23895 6276 23940 6304
rect 23934 6264 23940 6276
rect 23992 6264 23998 6316
rect 32214 6304 32220 6316
rect 32175 6276 32220 6304
rect 32214 6264 32220 6276
rect 32272 6264 32278 6316
rect 33336 6313 33364 6344
rect 33965 6341 33977 6344
rect 34011 6341 34023 6375
rect 33965 6335 34023 6341
rect 35894 6332 35900 6384
rect 35952 6372 35958 6384
rect 35952 6344 36124 6372
rect 35952 6332 35958 6344
rect 33321 6307 33379 6313
rect 33321 6273 33333 6307
rect 33367 6273 33379 6307
rect 33321 6267 33379 6273
rect 33505 6307 33563 6313
rect 33505 6273 33517 6307
rect 33551 6304 33563 6307
rect 34790 6304 34796 6316
rect 33551 6276 34796 6304
rect 33551 6273 33563 6276
rect 33505 6267 33563 6273
rect 34790 6264 34796 6276
rect 34848 6304 34854 6316
rect 35342 6304 35348 6316
rect 34848 6276 35348 6304
rect 34848 6264 34854 6276
rect 35342 6264 35348 6276
rect 35400 6264 35406 6316
rect 35805 6307 35863 6313
rect 35805 6273 35817 6307
rect 35851 6273 35863 6307
rect 35986 6304 35992 6316
rect 35947 6276 35992 6304
rect 35805 6267 35863 6273
rect 10226 6196 10232 6248
rect 10284 6236 10290 6248
rect 14829 6239 14887 6245
rect 14829 6236 14841 6239
rect 10284 6208 14841 6236
rect 10284 6196 10290 6208
rect 14829 6205 14841 6208
rect 14875 6236 14887 6239
rect 15562 6236 15568 6248
rect 14875 6208 15568 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 15562 6196 15568 6208
rect 15620 6236 15626 6248
rect 16482 6236 16488 6248
rect 15620 6208 16488 6236
rect 15620 6196 15626 6208
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 4154 6128 4160 6180
rect 4212 6168 4218 6180
rect 4706 6168 4712 6180
rect 4212 6140 4712 6168
rect 4212 6128 4218 6140
rect 4706 6128 4712 6140
rect 4764 6168 4770 6180
rect 5537 6171 5595 6177
rect 5537 6168 5549 6171
rect 4764 6140 5549 6168
rect 4764 6128 4770 6140
rect 5537 6137 5549 6140
rect 5583 6168 5595 6171
rect 10962 6168 10968 6180
rect 5583 6140 10968 6168
rect 5583 6137 5595 6140
rect 5537 6131 5595 6137
rect 10962 6128 10968 6140
rect 11020 6128 11026 6180
rect 14458 6128 14464 6180
rect 14516 6168 14522 6180
rect 17034 6168 17040 6180
rect 14516 6140 17040 6168
rect 14516 6128 14522 6140
rect 17034 6128 17040 6140
rect 17092 6128 17098 6180
rect 21082 6128 21088 6180
rect 21140 6168 21146 6180
rect 22186 6168 22192 6180
rect 21140 6140 22192 6168
rect 21140 6128 21146 6140
rect 22186 6128 22192 6140
rect 22244 6128 22250 6180
rect 23952 6168 23980 6264
rect 25777 6239 25835 6245
rect 25777 6205 25789 6239
rect 25823 6236 25835 6239
rect 30282 6236 30288 6248
rect 25823 6208 30288 6236
rect 25823 6205 25835 6208
rect 25777 6199 25835 6205
rect 30282 6196 30288 6208
rect 30340 6236 30346 6248
rect 32490 6236 32496 6248
rect 30340 6208 32496 6236
rect 30340 6196 30346 6208
rect 32490 6196 32496 6208
rect 32548 6196 32554 6248
rect 33594 6196 33600 6248
rect 33652 6236 33658 6248
rect 35253 6239 35311 6245
rect 35253 6236 35265 6239
rect 33652 6208 35265 6236
rect 33652 6196 33658 6208
rect 35253 6205 35265 6208
rect 35299 6236 35311 6239
rect 35820 6236 35848 6267
rect 35986 6264 35992 6276
rect 36044 6264 36050 6316
rect 36096 6313 36124 6344
rect 36188 6313 36216 6412
rect 36446 6400 36452 6412
rect 36504 6400 36510 6452
rect 36081 6307 36139 6313
rect 36081 6273 36093 6307
rect 36127 6273 36139 6307
rect 36081 6267 36139 6273
rect 36173 6307 36231 6313
rect 36173 6273 36185 6307
rect 36219 6273 36231 6307
rect 37826 6304 37832 6316
rect 37787 6276 37832 6304
rect 36173 6267 36231 6273
rect 37826 6264 37832 6276
rect 37884 6264 37890 6316
rect 35299 6208 35848 6236
rect 35299 6205 35311 6208
rect 35253 6199 35311 6205
rect 29822 6168 29828 6180
rect 23952 6140 29828 6168
rect 29822 6128 29828 6140
rect 29880 6128 29886 6180
rect 4433 6103 4491 6109
rect 4433 6069 4445 6103
rect 4479 6100 4491 6103
rect 4614 6100 4620 6112
rect 4479 6072 4620 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 14185 6103 14243 6109
rect 14185 6069 14197 6103
rect 14231 6100 14243 6103
rect 14274 6100 14280 6112
rect 14231 6072 14280 6100
rect 14231 6069 14243 6072
rect 14185 6063 14243 6069
rect 14274 6060 14280 6072
rect 14332 6060 14338 6112
rect 20441 6103 20499 6109
rect 20441 6069 20453 6103
rect 20487 6100 20499 6103
rect 20714 6100 20720 6112
rect 20487 6072 20720 6100
rect 20487 6069 20499 6072
rect 20441 6063 20499 6069
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 20898 6100 20904 6112
rect 20859 6072 20904 6100
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 32214 6100 32220 6112
rect 32175 6072 32220 6100
rect 32214 6060 32220 6072
rect 32272 6060 32278 6112
rect 38010 6100 38016 6112
rect 37971 6072 38016 6100
rect 38010 6060 38016 6072
rect 38068 6060 38074 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 2498 5856 2504 5908
rect 2556 5896 2562 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 2556 5868 2697 5896
rect 2556 5856 2562 5868
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4341 5899 4399 5905
rect 4341 5896 4353 5899
rect 4028 5868 4353 5896
rect 4028 5856 4034 5868
rect 4341 5865 4353 5868
rect 4387 5865 4399 5899
rect 4341 5859 4399 5865
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 19702 5896 19708 5908
rect 11020 5868 19708 5896
rect 11020 5856 11026 5868
rect 19702 5856 19708 5868
rect 19760 5856 19766 5908
rect 25958 5896 25964 5908
rect 19812 5868 25964 5896
rect 4522 5788 4528 5840
rect 4580 5828 4586 5840
rect 4890 5828 4896 5840
rect 4580 5800 4896 5828
rect 4580 5788 4586 5800
rect 4890 5788 4896 5800
rect 4948 5828 4954 5840
rect 9033 5831 9091 5837
rect 9033 5828 9045 5831
rect 4948 5800 9045 5828
rect 4948 5788 4954 5800
rect 4706 5760 4712 5772
rect 4448 5732 4712 5760
rect 2866 5692 2872 5704
rect 2827 5664 2872 5692
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 4448 5624 4476 5732
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 5626 5720 5632 5772
rect 5684 5760 5690 5772
rect 8128 5769 8156 5800
rect 9033 5797 9045 5800
rect 9079 5828 9091 5831
rect 19812 5828 19840 5868
rect 25958 5856 25964 5868
rect 26016 5856 26022 5908
rect 9079 5800 19840 5828
rect 9079 5797 9091 5800
rect 9033 5791 9091 5797
rect 20714 5788 20720 5840
rect 20772 5828 20778 5840
rect 32214 5828 32220 5840
rect 20772 5800 32220 5828
rect 20772 5788 20778 5800
rect 32214 5788 32220 5800
rect 32272 5788 32278 5840
rect 5997 5763 6055 5769
rect 5997 5760 6009 5763
rect 5684 5732 6009 5760
rect 5684 5720 5690 5732
rect 5997 5729 6009 5732
rect 6043 5729 6055 5763
rect 5997 5723 6055 5729
rect 8113 5763 8171 5769
rect 8113 5729 8125 5763
rect 8159 5729 8171 5763
rect 8113 5723 8171 5729
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4893 5695 4951 5701
rect 4571 5664 4844 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4617 5627 4675 5633
rect 4617 5624 4629 5627
rect 4448 5596 4629 5624
rect 4617 5593 4629 5596
rect 4663 5593 4675 5627
rect 4617 5587 4675 5593
rect 4709 5627 4767 5633
rect 4709 5593 4721 5627
rect 4755 5593 4767 5627
rect 4816 5624 4844 5664
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 5534 5692 5540 5704
rect 4939 5664 5540 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5692 5779 5695
rect 5810 5692 5816 5704
rect 5767 5664 5816 5692
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 5166 5624 5172 5636
rect 4816 5596 5172 5624
rect 4709 5587 4767 5593
rect 3878 5556 3884 5568
rect 3839 5528 3884 5556
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 4724 5556 4752 5587
rect 5166 5584 5172 5596
rect 5224 5584 5230 5636
rect 6012 5624 6040 5723
rect 15654 5720 15660 5772
rect 15712 5760 15718 5772
rect 16301 5763 16359 5769
rect 16301 5760 16313 5763
rect 15712 5732 16313 5760
rect 15712 5720 15718 5732
rect 16301 5729 16313 5732
rect 16347 5729 16359 5763
rect 16301 5723 16359 5729
rect 19426 5720 19432 5772
rect 19484 5760 19490 5772
rect 19797 5763 19855 5769
rect 19797 5760 19809 5763
rect 19484 5732 19809 5760
rect 19484 5720 19490 5732
rect 19797 5729 19809 5732
rect 19843 5729 19855 5763
rect 19797 5723 19855 5729
rect 7926 5692 7932 5704
rect 7887 5664 7932 5692
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 10226 5692 10232 5704
rect 10187 5664 10232 5692
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 14274 5692 14280 5704
rect 14235 5664 14280 5692
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 14366 5652 14372 5704
rect 14424 5692 14430 5704
rect 14645 5695 14703 5701
rect 14424 5664 14469 5692
rect 14424 5652 14430 5664
rect 14645 5661 14657 5695
rect 14691 5692 14703 5695
rect 14691 5664 15240 5692
rect 14691 5661 14703 5664
rect 14645 5655 14703 5661
rect 6730 5624 6736 5636
rect 6012 5596 6736 5624
rect 6730 5584 6736 5596
rect 6788 5624 6794 5636
rect 6788 5596 10364 5624
rect 6788 5584 6794 5596
rect 10336 5568 10364 5596
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 14516 5596 14561 5624
rect 14516 5584 14522 5596
rect 15212 5568 15240 5664
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 19702 5692 19708 5704
rect 19392 5664 19708 5692
rect 19392 5652 19398 5664
rect 19702 5652 19708 5664
rect 19760 5652 19766 5704
rect 5353 5559 5411 5565
rect 5353 5556 5365 5559
rect 4724 5528 5365 5556
rect 5353 5525 5365 5528
rect 5399 5525 5411 5559
rect 5353 5519 5411 5525
rect 5810 5516 5816 5568
rect 5868 5556 5874 5568
rect 6638 5556 6644 5568
rect 5868 5528 5913 5556
rect 6599 5528 6644 5556
rect 5868 5516 5874 5528
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 7745 5559 7803 5565
rect 7745 5525 7757 5559
rect 7791 5556 7803 5559
rect 7926 5556 7932 5568
rect 7791 5528 7932 5556
rect 7791 5525 7803 5528
rect 7745 5519 7803 5525
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 10318 5556 10324 5568
rect 10279 5528 10324 5556
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 14093 5559 14151 5565
rect 14093 5525 14105 5559
rect 14139 5556 14151 5559
rect 14274 5556 14280 5568
rect 14139 5528 14280 5556
rect 14139 5525 14151 5528
rect 14093 5519 14151 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 15194 5556 15200 5568
rect 15155 5528 15200 5556
rect 15194 5516 15200 5528
rect 15252 5516 15258 5568
rect 19242 5556 19248 5568
rect 19203 5528 19248 5556
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19613 5559 19671 5565
rect 19613 5556 19625 5559
rect 19392 5528 19625 5556
rect 19392 5516 19398 5528
rect 19613 5525 19625 5528
rect 19659 5525 19671 5559
rect 19812 5556 19840 5723
rect 19886 5720 19892 5772
rect 19944 5760 19950 5772
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 19944 5732 22477 5760
rect 19944 5720 19950 5732
rect 22465 5729 22477 5732
rect 22511 5760 22523 5763
rect 23750 5760 23756 5772
rect 22511 5732 23756 5760
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 23750 5720 23756 5732
rect 23808 5720 23814 5772
rect 26142 5720 26148 5772
rect 26200 5760 26206 5772
rect 26697 5763 26755 5769
rect 26697 5760 26709 5763
rect 26200 5732 26709 5760
rect 26200 5720 26206 5732
rect 26697 5729 26709 5732
rect 26743 5760 26755 5763
rect 26743 5732 28580 5760
rect 26743 5729 26755 5732
rect 26697 5723 26755 5729
rect 20438 5692 20444 5704
rect 20399 5664 20444 5692
rect 20438 5652 20444 5664
rect 20496 5652 20502 5704
rect 22005 5695 22063 5701
rect 22005 5661 22017 5695
rect 22051 5661 22063 5695
rect 22005 5655 22063 5661
rect 19886 5584 19892 5636
rect 19944 5624 19950 5636
rect 20714 5624 20720 5636
rect 19944 5596 20720 5624
rect 19944 5584 19950 5596
rect 20714 5584 20720 5596
rect 20772 5584 20778 5636
rect 22020 5624 22048 5655
rect 26786 5652 26792 5704
rect 26844 5692 26850 5704
rect 26973 5695 27031 5701
rect 26973 5692 26985 5695
rect 26844 5664 26985 5692
rect 26844 5652 26850 5664
rect 26973 5661 26985 5664
rect 27019 5661 27031 5695
rect 28552 5692 28580 5732
rect 29086 5720 29092 5772
rect 29144 5760 29150 5772
rect 30101 5763 30159 5769
rect 30101 5760 30113 5763
rect 29144 5732 30113 5760
rect 29144 5720 29150 5732
rect 30101 5729 30113 5732
rect 30147 5729 30159 5763
rect 30282 5760 30288 5772
rect 30243 5732 30288 5760
rect 30101 5723 30159 5729
rect 30282 5720 30288 5732
rect 30340 5720 30346 5772
rect 30558 5720 30564 5772
rect 30616 5760 30622 5772
rect 31573 5763 31631 5769
rect 31573 5760 31585 5763
rect 30616 5732 31585 5760
rect 30616 5720 30622 5732
rect 31573 5729 31585 5732
rect 31619 5729 31631 5763
rect 31573 5723 31631 5729
rect 30374 5692 30380 5704
rect 28552 5664 30380 5692
rect 26973 5655 27031 5661
rect 30374 5652 30380 5664
rect 30432 5652 30438 5704
rect 31389 5695 31447 5701
rect 31389 5692 31401 5695
rect 30760 5664 31401 5692
rect 22020 5596 22140 5624
rect 20622 5556 20628 5568
rect 19812 5528 20628 5556
rect 19613 5519 19671 5525
rect 20622 5516 20628 5528
rect 20680 5516 20686 5568
rect 22112 5556 22140 5596
rect 22186 5584 22192 5636
rect 22244 5624 22250 5636
rect 22244 5596 22289 5624
rect 22244 5584 22250 5596
rect 24762 5584 24768 5636
rect 24820 5624 24826 5636
rect 27798 5624 27804 5636
rect 24820 5596 27804 5624
rect 24820 5584 24826 5596
rect 27798 5584 27804 5596
rect 27856 5584 27862 5636
rect 29822 5584 29828 5636
rect 29880 5624 29886 5636
rect 30650 5624 30656 5636
rect 29880 5596 30656 5624
rect 29880 5584 29886 5596
rect 23474 5556 23480 5568
rect 22112 5528 23480 5556
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 30392 5565 30420 5596
rect 30650 5584 30656 5596
rect 30708 5584 30714 5636
rect 30760 5565 30788 5664
rect 31389 5661 31401 5664
rect 31435 5661 31447 5695
rect 31389 5655 31447 5661
rect 30377 5559 30435 5565
rect 30377 5525 30389 5559
rect 30423 5525 30435 5559
rect 30377 5519 30435 5525
rect 30745 5559 30803 5565
rect 30745 5525 30757 5559
rect 30791 5525 30803 5559
rect 30745 5519 30803 5525
rect 31018 5516 31024 5568
rect 31076 5556 31082 5568
rect 31205 5559 31263 5565
rect 31205 5556 31217 5559
rect 31076 5528 31217 5556
rect 31076 5516 31082 5528
rect 31205 5525 31217 5528
rect 31251 5525 31263 5559
rect 31205 5519 31263 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 2590 5352 2596 5364
rect 1627 5324 2596 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 4522 5352 4528 5364
rect 4483 5324 4528 5352
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 6917 5355 6975 5361
rect 6917 5321 6929 5355
rect 6963 5352 6975 5355
rect 8389 5355 8447 5361
rect 8389 5352 8401 5355
rect 6963 5324 8401 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 8389 5321 8401 5324
rect 8435 5321 8447 5355
rect 8754 5352 8760 5364
rect 8715 5324 8760 5352
rect 8389 5315 8447 5321
rect 5353 5287 5411 5293
rect 5353 5253 5365 5287
rect 5399 5284 5411 5287
rect 6472 5284 6500 5315
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 10505 5355 10563 5361
rect 10505 5321 10517 5355
rect 10551 5352 10563 5355
rect 11885 5355 11943 5361
rect 11885 5352 11897 5355
rect 10551 5324 11897 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 11885 5321 11897 5324
rect 11931 5321 11943 5355
rect 11885 5315 11943 5321
rect 12345 5355 12403 5361
rect 12345 5321 12357 5355
rect 12391 5352 12403 5355
rect 14550 5352 14556 5364
rect 12391 5324 14556 5352
rect 12391 5321 12403 5324
rect 12345 5315 12403 5321
rect 14550 5312 14556 5324
rect 14608 5312 14614 5364
rect 15470 5352 15476 5364
rect 15431 5324 15476 5352
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 19426 5352 19432 5364
rect 18340 5324 19432 5352
rect 18340 5284 18368 5324
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 20714 5352 20720 5364
rect 20675 5324 20720 5352
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 26326 5352 26332 5364
rect 26287 5324 26332 5352
rect 26326 5312 26332 5324
rect 26384 5352 26390 5364
rect 27617 5355 27675 5361
rect 27617 5352 27629 5355
rect 26384 5324 27629 5352
rect 26384 5312 26390 5324
rect 27617 5321 27629 5324
rect 27663 5321 27675 5355
rect 28442 5352 28448 5364
rect 28403 5324 28448 5352
rect 27617 5315 27675 5321
rect 28442 5312 28448 5324
rect 28500 5312 28506 5364
rect 29822 5352 29828 5364
rect 29783 5324 29828 5352
rect 29822 5312 29828 5324
rect 29880 5312 29886 5364
rect 30558 5312 30564 5364
rect 30616 5352 30622 5364
rect 31021 5355 31079 5361
rect 31021 5352 31033 5355
rect 30616 5324 31033 5352
rect 30616 5312 30622 5324
rect 31021 5321 31033 5324
rect 31067 5321 31079 5355
rect 31021 5315 31079 5321
rect 5399 5256 6500 5284
rect 9048 5256 18368 5284
rect 18417 5287 18475 5293
rect 5399 5253 5411 5256
rect 5353 5247 5411 5253
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5216 1458 5228
rect 2041 5219 2099 5225
rect 2041 5216 2053 5219
rect 1452 5188 2053 5216
rect 1452 5176 1458 5188
rect 2041 5185 2053 5188
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5216 3847 5219
rect 4614 5216 4620 5228
rect 3835 5188 4620 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 5166 5216 5172 5228
rect 5127 5188 5172 5216
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5185 5319 5219
rect 5534 5216 5540 5228
rect 5447 5188 5540 5216
rect 5261 5179 5319 5185
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 3988 5080 4016 5111
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 5276 5148 5304 5179
rect 5534 5176 5540 5188
rect 5592 5216 5598 5228
rect 6638 5216 6644 5228
rect 5592 5188 6644 5216
rect 5592 5176 5598 5188
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 6822 5216 6828 5228
rect 6783 5188 6828 5216
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 9048 5160 9076 5256
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 10643 5188 10732 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 5718 5148 5724 5160
rect 4212 5120 5724 5148
rect 4212 5108 4218 5120
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 7009 5151 7067 5157
rect 7009 5148 7021 5151
rect 6788 5120 7021 5148
rect 6788 5108 6794 5120
rect 7009 5117 7021 5120
rect 7055 5117 7067 5151
rect 7009 5111 7067 5117
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 4522 5080 4528 5092
rect 3988 5052 4528 5080
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 8864 5080 8892 5111
rect 9030 5108 9036 5160
rect 9088 5148 9094 5160
rect 10318 5148 10324 5160
rect 9088 5120 9181 5148
rect 10279 5120 10324 5148
rect 9088 5108 9094 5120
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 9766 5080 9772 5092
rect 8864 5052 9772 5080
rect 9766 5040 9772 5052
rect 9824 5080 9830 5092
rect 10704 5080 10732 5188
rect 10778 5176 10784 5228
rect 10836 5216 10842 5228
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 10836 5188 12265 5216
rect 10836 5176 10842 5188
rect 12253 5185 12265 5188
rect 12299 5216 12311 5219
rect 12526 5216 12532 5228
rect 12299 5188 12532 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12636 5148 12664 5256
rect 18417 5253 18429 5287
rect 18463 5284 18475 5287
rect 19242 5284 19248 5296
rect 18463 5256 19248 5284
rect 18463 5253 18475 5256
rect 18417 5247 18475 5253
rect 19242 5244 19248 5256
rect 19300 5244 19306 5296
rect 19334 5244 19340 5296
rect 19392 5284 19398 5296
rect 20073 5287 20131 5293
rect 20073 5284 20085 5287
rect 19392 5256 20085 5284
rect 19392 5244 19398 5256
rect 20073 5253 20085 5256
rect 20119 5284 20131 5287
rect 20254 5284 20260 5296
rect 20119 5256 20260 5284
rect 20119 5253 20131 5256
rect 20073 5247 20131 5253
rect 20254 5244 20260 5256
rect 20312 5244 20318 5296
rect 15565 5219 15623 5225
rect 15304 5188 15516 5216
rect 15304 5157 15332 5188
rect 12483 5120 12664 5148
rect 15289 5151 15347 5157
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 15289 5117 15301 5151
rect 15335 5117 15347 5151
rect 15488 5148 15516 5188
rect 15565 5185 15577 5219
rect 15611 5216 15623 5219
rect 15838 5216 15844 5228
rect 15611 5188 15844 5216
rect 15611 5185 15623 5188
rect 15565 5179 15623 5185
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 17034 5176 17040 5228
rect 17092 5216 17098 5228
rect 18233 5219 18291 5225
rect 18233 5216 18245 5219
rect 17092 5188 18245 5216
rect 17092 5176 17098 5188
rect 18233 5185 18245 5188
rect 18279 5185 18291 5219
rect 18506 5216 18512 5228
rect 18467 5188 18512 5216
rect 18233 5179 18291 5185
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 18601 5219 18659 5225
rect 18601 5185 18613 5219
rect 18647 5216 18659 5219
rect 19702 5216 19708 5228
rect 18647 5188 19708 5216
rect 18647 5185 18659 5188
rect 18601 5179 18659 5185
rect 19702 5176 19708 5188
rect 19760 5176 19766 5228
rect 26206 5188 27936 5216
rect 15654 5148 15660 5160
rect 15488 5120 15660 5148
rect 15289 5111 15347 5117
rect 15654 5108 15660 5120
rect 15712 5108 15718 5160
rect 25038 5108 25044 5160
rect 25096 5148 25102 5160
rect 26206 5148 26234 5188
rect 27706 5148 27712 5160
rect 25096 5120 26234 5148
rect 27667 5120 27712 5148
rect 25096 5108 25102 5120
rect 27706 5108 27712 5120
rect 27764 5108 27770 5160
rect 27908 5157 27936 5188
rect 27893 5151 27951 5157
rect 27893 5117 27905 5151
rect 27939 5148 27951 5151
rect 29086 5148 29092 5160
rect 27939 5120 29092 5148
rect 27939 5117 27951 5120
rect 27893 5111 27951 5117
rect 29086 5108 29092 5120
rect 29144 5108 29150 5160
rect 9824 5052 12434 5080
rect 9824 5040 9830 5052
rect 3234 4972 3240 5024
rect 3292 5012 3298 5024
rect 3605 5015 3663 5021
rect 3605 5012 3617 5015
rect 3292 4984 3617 5012
rect 3292 4972 3298 4984
rect 3605 4981 3617 4984
rect 3651 4981 3663 5015
rect 4982 5012 4988 5024
rect 4943 4984 4988 5012
rect 3605 4975 3663 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 10744 4984 10977 5012
rect 10744 4972 10750 4984
rect 10965 4981 10977 4984
rect 11011 4981 11023 5015
rect 12406 5012 12434 5052
rect 15194 5040 15200 5092
rect 15252 5080 15258 5092
rect 26326 5080 26332 5092
rect 15252 5052 26332 5080
rect 15252 5040 15258 5052
rect 26326 5040 26332 5052
rect 26384 5040 26390 5092
rect 15286 5012 15292 5024
rect 12406 4984 15292 5012
rect 10965 4975 11023 4981
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 15930 5012 15936 5024
rect 15891 4984 15936 5012
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 18785 5015 18843 5021
rect 18785 4981 18797 5015
rect 18831 5012 18843 5015
rect 19150 5012 19156 5024
rect 18831 4984 19156 5012
rect 18831 4981 18843 4984
rect 18785 4975 18843 4981
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 26970 4972 26976 5024
rect 27028 5012 27034 5024
rect 27249 5015 27307 5021
rect 27249 5012 27261 5015
rect 27028 4984 27261 5012
rect 27028 4972 27034 4984
rect 27249 4981 27261 4984
rect 27295 4981 27307 5015
rect 34698 5012 34704 5024
rect 34659 4984 34704 5012
rect 27249 4975 27307 4981
rect 34698 4972 34704 4984
rect 34756 4972 34762 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 4893 4811 4951 4817
rect 4893 4808 4905 4811
rect 4672 4780 4905 4808
rect 4672 4768 4678 4780
rect 4893 4777 4905 4780
rect 4939 4777 4951 4811
rect 4893 4771 4951 4777
rect 5810 4768 5816 4820
rect 5868 4808 5874 4820
rect 6825 4811 6883 4817
rect 6825 4808 6837 4811
rect 5868 4780 6837 4808
rect 5868 4768 5874 4780
rect 6825 4777 6837 4780
rect 6871 4777 6883 4811
rect 14458 4808 14464 4820
rect 6825 4771 6883 4777
rect 10888 4780 14464 4808
rect 4065 4675 4123 4681
rect 4065 4641 4077 4675
rect 4111 4672 4123 4675
rect 4632 4672 4660 4768
rect 5166 4700 5172 4752
rect 5224 4740 5230 4752
rect 10888 4740 10916 4780
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 15838 4808 15844 4820
rect 15799 4780 15844 4808
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 19702 4808 19708 4820
rect 19663 4780 19708 4808
rect 19702 4768 19708 4780
rect 19760 4768 19766 4820
rect 23750 4808 23756 4820
rect 23711 4780 23756 4808
rect 23750 4768 23756 4780
rect 23808 4808 23814 4820
rect 24762 4808 24768 4820
rect 23808 4780 24768 4808
rect 23808 4768 23814 4780
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 35253 4811 35311 4817
rect 35253 4777 35265 4811
rect 35299 4808 35311 4811
rect 35894 4808 35900 4820
rect 35299 4780 35900 4808
rect 35299 4777 35311 4780
rect 35253 4771 35311 4777
rect 35894 4768 35900 4780
rect 35952 4808 35958 4820
rect 36357 4811 36415 4817
rect 36357 4808 36369 4811
rect 35952 4780 36369 4808
rect 35952 4768 35958 4780
rect 36357 4777 36369 4780
rect 36403 4777 36415 4811
rect 36357 4771 36415 4777
rect 5224 4712 10916 4740
rect 5224 4700 5230 4712
rect 4111 4644 4660 4672
rect 6273 4675 6331 4681
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 6638 4672 6644 4684
rect 6319 4644 6644 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6638 4632 6644 4644
rect 6696 4672 6702 4684
rect 7374 4672 7380 4684
rect 6696 4644 7380 4672
rect 6696 4632 6702 4644
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4672 7527 4675
rect 9030 4672 9036 4684
rect 7515 4644 9036 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 9030 4632 9036 4644
rect 9088 4632 9094 4684
rect 10778 4672 10784 4684
rect 10428 4644 10784 4672
rect 3234 4604 3240 4616
rect 3195 4576 3240 4604
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 4982 4604 4988 4616
rect 4295 4576 4988 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5718 4604 5724 4616
rect 5679 4576 5724 4604
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 7282 4564 7288 4616
rect 7340 4604 7346 4616
rect 10428 4604 10456 4644
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 7340 4576 10456 4604
rect 7340 4564 7346 4576
rect 10502 4564 10508 4616
rect 10560 4604 10566 4616
rect 10686 4604 10692 4616
rect 10560 4576 10605 4604
rect 10647 4576 10692 4604
rect 10560 4564 10566 4576
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 10888 4613 10916 4712
rect 11057 4743 11115 4749
rect 11057 4709 11069 4743
rect 11103 4709 11115 4743
rect 11057 4703 11115 4709
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 11072 4604 11100 4703
rect 12434 4700 12440 4752
rect 12492 4740 12498 4752
rect 17126 4740 17132 4752
rect 12492 4712 12537 4740
rect 15212 4712 17132 4740
rect 12492 4700 12498 4712
rect 15212 4684 15240 4712
rect 17126 4700 17132 4712
rect 17184 4700 17190 4752
rect 37734 4740 37740 4752
rect 26206 4712 37740 4740
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4672 14519 4675
rect 14642 4672 14648 4684
rect 14507 4644 14648 4672
rect 14507 4641 14519 4644
rect 14461 4635 14519 4641
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 15194 4672 15200 4684
rect 15155 4644 15200 4672
rect 15194 4632 15200 4644
rect 15252 4632 15258 4684
rect 15930 4632 15936 4684
rect 15988 4672 15994 4684
rect 20165 4675 20223 4681
rect 20165 4672 20177 4675
rect 15988 4644 20177 4672
rect 15988 4632 15994 4644
rect 20165 4641 20177 4644
rect 20211 4641 20223 4675
rect 20165 4635 20223 4641
rect 20349 4675 20407 4681
rect 20349 4641 20361 4675
rect 20395 4672 20407 4675
rect 22922 4672 22928 4684
rect 20395 4644 22928 4672
rect 20395 4641 20407 4644
rect 20349 4635 20407 4641
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 25038 4672 25044 4684
rect 24999 4644 25044 4672
rect 25038 4632 25044 4644
rect 25096 4632 25102 4684
rect 11701 4607 11759 4613
rect 11701 4604 11713 4607
rect 11072 4576 11713 4604
rect 10873 4567 10931 4573
rect 11701 4573 11713 4576
rect 11747 4573 11759 4607
rect 11882 4604 11888 4616
rect 11843 4576 11888 4604
rect 11701 4567 11759 4573
rect 11882 4564 11888 4576
rect 11940 4564 11946 4616
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14550 4564 14556 4616
rect 14608 4604 14614 4616
rect 15473 4607 15531 4613
rect 15473 4604 15485 4607
rect 14608 4576 15485 4604
rect 14608 4564 14614 4576
rect 15473 4573 15485 4576
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 17862 4564 17868 4616
rect 17920 4604 17926 4616
rect 18049 4607 18107 4613
rect 18049 4604 18061 4607
rect 17920 4576 18061 4604
rect 17920 4564 17926 4576
rect 18049 4573 18061 4576
rect 18095 4573 18107 4607
rect 18230 4604 18236 4616
rect 18191 4576 18236 4604
rect 18049 4567 18107 4573
rect 18230 4564 18236 4576
rect 18288 4564 18294 4616
rect 20073 4607 20131 4613
rect 20073 4573 20085 4607
rect 20119 4604 20131 4607
rect 20990 4604 20996 4616
rect 20119 4576 20996 4604
rect 20119 4573 20131 4576
rect 20073 4567 20131 4573
rect 20990 4564 20996 4576
rect 21048 4604 21054 4616
rect 26206 4604 26234 4712
rect 37734 4700 37740 4712
rect 37792 4700 37798 4752
rect 26786 4672 26792 4684
rect 26747 4644 26792 4672
rect 26786 4632 26792 4644
rect 26844 4632 26850 4684
rect 28074 4672 28080 4684
rect 28035 4644 28080 4672
rect 28074 4632 28080 4644
rect 28132 4632 28138 4684
rect 28261 4675 28319 4681
rect 28261 4641 28273 4675
rect 28307 4672 28319 4675
rect 29086 4672 29092 4684
rect 28307 4644 29092 4672
rect 28307 4641 28319 4644
rect 28261 4635 28319 4641
rect 29086 4632 29092 4644
rect 29144 4632 29150 4684
rect 34606 4632 34612 4684
rect 34664 4672 34670 4684
rect 35345 4675 35403 4681
rect 35345 4672 35357 4675
rect 34664 4644 35357 4672
rect 34664 4632 34670 4644
rect 35345 4641 35357 4644
rect 35391 4672 35403 4675
rect 35391 4644 37044 4672
rect 35391 4641 35403 4644
rect 35345 4635 35403 4641
rect 26970 4604 26976 4616
rect 21048 4576 26234 4604
rect 26931 4576 26976 4604
rect 21048 4564 21054 4576
rect 26970 4564 26976 4576
rect 27028 4564 27034 4616
rect 27157 4607 27215 4613
rect 27157 4573 27169 4607
rect 27203 4604 27215 4607
rect 28813 4607 28871 4613
rect 28813 4604 28825 4607
rect 27203 4576 28825 4604
rect 27203 4573 27215 4576
rect 27157 4567 27215 4573
rect 28813 4573 28825 4576
rect 28859 4573 28871 4607
rect 31018 4604 31024 4616
rect 30979 4576 31024 4604
rect 28813 4567 28871 4573
rect 31018 4564 31024 4576
rect 31076 4564 31082 4616
rect 34790 4564 34796 4616
rect 34848 4613 34854 4616
rect 37016 4613 37044 4644
rect 34848 4607 34884 4613
rect 34872 4604 34884 4607
rect 35930 4607 35988 4613
rect 35930 4604 35942 4607
rect 34872 4576 35942 4604
rect 34872 4573 34884 4576
rect 34848 4567 34884 4573
rect 35930 4573 35942 4576
rect 35976 4573 35988 4607
rect 35930 4567 35988 4573
rect 36449 4607 36507 4613
rect 36449 4573 36461 4607
rect 36495 4604 36507 4607
rect 36909 4607 36967 4613
rect 36909 4604 36921 4607
rect 36495 4576 36921 4604
rect 36495 4573 36507 4576
rect 36449 4567 36507 4573
rect 36909 4573 36921 4576
rect 36955 4573 36967 4607
rect 36909 4567 36967 4573
rect 37001 4607 37059 4613
rect 37001 4573 37013 4607
rect 37047 4573 37059 4607
rect 37001 4567 37059 4573
rect 34848 4564 34854 4567
rect 5442 4496 5448 4548
rect 5500 4536 5506 4548
rect 5500 4508 7236 4536
rect 5500 4496 5506 4508
rect 3053 4471 3111 4477
rect 3053 4437 3065 4471
rect 3099 4468 3111 4471
rect 3142 4468 3148 4480
rect 3099 4440 3148 4468
rect 3099 4437 3111 4440
rect 3053 4431 3111 4437
rect 3142 4428 3148 4440
rect 3200 4428 3206 4480
rect 4430 4468 4436 4480
rect 4391 4440 4436 4468
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 7208 4477 7236 4508
rect 7374 4496 7380 4548
rect 7432 4536 7438 4548
rect 10520 4536 10548 4564
rect 10778 4536 10784 4548
rect 7432 4508 10548 4536
rect 10739 4508 10784 4536
rect 7432 4496 7438 4508
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 15381 4539 15439 4545
rect 15381 4505 15393 4539
rect 15427 4536 15439 4539
rect 16390 4536 16396 4548
rect 15427 4508 16396 4536
rect 15427 4505 15439 4508
rect 15381 4499 15439 4505
rect 16390 4496 16396 4508
rect 16448 4536 16454 4548
rect 16850 4536 16856 4548
rect 16448 4508 16856 4536
rect 16448 4496 16454 4508
rect 16850 4496 16856 4508
rect 16908 4496 16914 4548
rect 23474 4496 23480 4548
rect 23532 4536 23538 4548
rect 24857 4539 24915 4545
rect 24857 4536 24869 4539
rect 23532 4508 24869 4536
rect 23532 4496 23538 4508
rect 24857 4505 24869 4508
rect 24903 4505 24915 4539
rect 24857 4499 24915 4505
rect 27985 4539 28043 4545
rect 27985 4505 27997 4539
rect 28031 4536 28043 4539
rect 29178 4536 29184 4548
rect 28031 4508 29184 4536
rect 28031 4505 28043 4508
rect 27985 4499 28043 4505
rect 29178 4496 29184 4508
rect 29236 4496 29242 4548
rect 7193 4471 7251 4477
rect 7193 4437 7205 4471
rect 7239 4437 7251 4471
rect 11514 4468 11520 4480
rect 11475 4440 11520 4468
rect 7193 4431 7251 4437
rect 11514 4428 11520 4440
rect 11572 4428 11578 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14093 4471 14151 4477
rect 14093 4468 14105 4471
rect 13872 4440 14105 4468
rect 13872 4428 13878 4440
rect 14093 4437 14105 4440
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 17310 4428 17316 4480
rect 17368 4468 17374 4480
rect 17865 4471 17923 4477
rect 17865 4468 17877 4471
rect 17368 4440 17877 4468
rect 17368 4428 17374 4440
rect 17865 4437 17877 4440
rect 17911 4437 17923 4471
rect 17865 4431 17923 4437
rect 24397 4471 24455 4477
rect 24397 4437 24409 4471
rect 24443 4468 24455 4471
rect 24670 4468 24676 4480
rect 24443 4440 24676 4468
rect 24443 4437 24455 4440
rect 24397 4431 24455 4437
rect 24670 4428 24676 4440
rect 24728 4428 24734 4480
rect 24762 4428 24768 4480
rect 24820 4468 24826 4480
rect 27614 4468 27620 4480
rect 24820 4440 24865 4468
rect 27575 4440 27620 4468
rect 24820 4428 24826 4440
rect 27614 4428 27620 4440
rect 27672 4428 27678 4480
rect 28997 4471 29055 4477
rect 28997 4437 29009 4471
rect 29043 4468 29055 4471
rect 29086 4468 29092 4480
rect 29043 4440 29092 4468
rect 29043 4437 29055 4440
rect 28997 4431 29055 4437
rect 29086 4428 29092 4440
rect 29144 4428 29150 4480
rect 31202 4468 31208 4480
rect 31163 4440 31208 4468
rect 31202 4428 31208 4440
rect 31260 4428 31266 4480
rect 34514 4428 34520 4480
rect 34572 4468 34578 4480
rect 34701 4471 34759 4477
rect 34701 4468 34713 4471
rect 34572 4440 34713 4468
rect 34572 4428 34578 4440
rect 34701 4437 34713 4440
rect 34747 4437 34759 4471
rect 34701 4431 34759 4437
rect 34790 4428 34796 4480
rect 34848 4468 34854 4480
rect 34885 4471 34943 4477
rect 34885 4468 34897 4471
rect 34848 4440 34897 4468
rect 34848 4428 34854 4440
rect 34885 4437 34897 4440
rect 34931 4437 34943 4471
rect 35802 4468 35808 4480
rect 35763 4440 35808 4468
rect 34885 4431 34943 4437
rect 35802 4428 35808 4440
rect 35860 4428 35866 4480
rect 35989 4471 36047 4477
rect 35989 4437 36001 4471
rect 36035 4468 36047 4471
rect 36262 4468 36268 4480
rect 36035 4440 36268 4468
rect 36035 4437 36047 4440
rect 35989 4431 36047 4437
rect 36262 4428 36268 4440
rect 36320 4428 36326 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 4249 4267 4307 4273
rect 4249 4233 4261 4267
rect 4295 4264 4307 4267
rect 5442 4264 5448 4276
rect 4295 4236 5448 4264
rect 4295 4233 4307 4236
rect 4249 4227 4307 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 11517 4267 11575 4273
rect 11517 4264 11529 4267
rect 10796 4236 11529 4264
rect 10796 4208 10824 4236
rect 11517 4233 11529 4236
rect 11563 4264 11575 4267
rect 11606 4264 11612 4276
rect 11563 4236 11612 4264
rect 11563 4233 11575 4236
rect 11517 4227 11575 4233
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 11882 4224 11888 4276
rect 11940 4264 11946 4276
rect 12069 4267 12127 4273
rect 12069 4264 12081 4267
rect 11940 4236 12081 4264
rect 11940 4224 11946 4236
rect 12069 4233 12081 4236
rect 12115 4264 12127 4267
rect 14642 4264 14648 4276
rect 12115 4236 14648 4264
rect 12115 4233 12127 4236
rect 12069 4227 12127 4233
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 15470 4224 15476 4276
rect 15528 4264 15534 4276
rect 15841 4267 15899 4273
rect 15841 4264 15853 4267
rect 15528 4236 15853 4264
rect 15528 4224 15534 4236
rect 15841 4233 15853 4236
rect 15887 4233 15899 4267
rect 15841 4227 15899 4233
rect 27706 4224 27712 4276
rect 27764 4264 27770 4276
rect 27985 4267 28043 4273
rect 27985 4264 27997 4267
rect 27764 4236 27997 4264
rect 27764 4224 27770 4236
rect 27985 4233 27997 4236
rect 28031 4233 28043 4267
rect 27985 4227 28043 4233
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 10778 4196 10784 4208
rect 4120 4168 10784 4196
rect 4120 4156 4126 4168
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 15286 4156 15292 4208
rect 15344 4196 15350 4208
rect 15344 4168 15516 4196
rect 15344 4156 15350 4168
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4128 1458 4140
rect 3142 4137 3148 4140
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 1452 4100 2053 4128
rect 1452 4088 1458 4100
rect 2041 4097 2053 4100
rect 2087 4097 2099 4131
rect 3136 4128 3148 4137
rect 3103 4100 3148 4128
rect 2041 4091 2099 4097
rect 3136 4091 3148 4100
rect 3142 4088 3148 4091
rect 3200 4088 3206 4140
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 4488 4100 4905 4128
rect 4488 4088 4494 4100
rect 4893 4097 4905 4100
rect 4939 4097 4951 4131
rect 7926 4128 7932 4140
rect 7887 4100 7932 4128
rect 4893 4091 4951 4097
rect 7926 4088 7932 4100
rect 7984 4088 7990 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 11514 4128 11520 4140
rect 10551 4100 11520 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 13814 4128 13820 4140
rect 13775 4100 13820 4128
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 15378 4128 15384 4140
rect 15339 4100 15384 4128
rect 15378 4088 15384 4100
rect 15436 4088 15442 4140
rect 15488 4137 15516 4168
rect 28966 4168 29224 4196
rect 15473 4131 15531 4137
rect 15473 4097 15485 4131
rect 15519 4097 15531 4131
rect 17310 4128 17316 4140
rect 17271 4100 17316 4128
rect 15473 4091 15531 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 19150 4128 19156 4140
rect 19111 4100 19156 4128
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 19337 4131 19395 4137
rect 19337 4097 19349 4131
rect 19383 4128 19395 4131
rect 19797 4131 19855 4137
rect 19797 4128 19809 4131
rect 19383 4100 19809 4128
rect 19383 4097 19395 4100
rect 19337 4091 19395 4097
rect 19797 4097 19809 4100
rect 19843 4097 19855 4131
rect 23474 4128 23480 4140
rect 19797 4091 19855 4097
rect 22112 4100 23152 4128
rect 23435 4100 23480 4128
rect 2866 4060 2872 4072
rect 2827 4032 2872 4060
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 15194 4060 15200 4072
rect 15155 4032 15200 4060
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 18969 4063 19027 4069
rect 18969 4060 18981 4063
rect 18288 4032 18981 4060
rect 18288 4020 18294 4032
rect 18969 4029 18981 4032
rect 19015 4060 19027 4063
rect 22112 4060 22140 4100
rect 19015 4032 22140 4060
rect 23017 4063 23075 4069
rect 19015 4029 19027 4032
rect 18969 4023 19027 4029
rect 23017 4029 23029 4063
rect 23063 4029 23075 4063
rect 23017 4023 23075 4029
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 2406 3992 2412 4004
rect 1627 3964 2412 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 2406 3952 2412 3964
rect 2464 3952 2470 4004
rect 15654 3952 15660 4004
rect 15712 3992 15718 4004
rect 23032 3992 23060 4023
rect 15712 3964 23060 3992
rect 23124 3992 23152 4100
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 23658 4128 23664 4140
rect 23619 4100 23664 4128
rect 23658 4088 23664 4100
rect 23716 4088 23722 4140
rect 24670 4128 24676 4140
rect 24631 4100 24676 4128
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 26786 4128 26792 4140
rect 26206 4100 26792 4128
rect 23750 4060 23756 4072
rect 23711 4032 23756 4060
rect 23750 4020 23756 4032
rect 23808 4020 23814 4072
rect 24857 4063 24915 4069
rect 24857 4029 24869 4063
rect 24903 4060 24915 4063
rect 26206 4060 26234 4100
rect 26786 4088 26792 4100
rect 26844 4128 26850 4140
rect 27157 4131 27215 4137
rect 27157 4128 27169 4131
rect 26844 4100 27169 4128
rect 26844 4088 26850 4100
rect 27157 4097 27169 4100
rect 27203 4097 27215 4131
rect 27157 4091 27215 4097
rect 27341 4131 27399 4137
rect 27341 4097 27353 4131
rect 27387 4128 27399 4131
rect 27614 4128 27620 4140
rect 27387 4100 27620 4128
rect 27387 4097 27399 4100
rect 27341 4091 27399 4097
rect 27614 4088 27620 4100
rect 27672 4088 27678 4140
rect 28810 4088 28816 4140
rect 28868 4128 28874 4140
rect 28966 4128 28994 4168
rect 29086 4128 29092 4140
rect 29144 4137 29150 4140
rect 28868 4100 28994 4128
rect 29056 4100 29092 4128
rect 28868 4088 28874 4100
rect 29086 4088 29092 4100
rect 29144 4091 29156 4137
rect 29196 4128 29224 4168
rect 29365 4131 29423 4137
rect 29365 4128 29377 4131
rect 29196 4100 29377 4128
rect 29365 4097 29377 4100
rect 29411 4128 29423 4131
rect 29638 4128 29644 4140
rect 29411 4100 29644 4128
rect 29411 4097 29423 4100
rect 29365 4091 29423 4097
rect 29144 4088 29150 4091
rect 29638 4088 29644 4100
rect 29696 4128 29702 4140
rect 29825 4131 29883 4137
rect 29825 4128 29837 4131
rect 29696 4100 29837 4128
rect 29696 4088 29702 4100
rect 29825 4097 29837 4100
rect 29871 4097 29883 4131
rect 33870 4128 33876 4140
rect 33831 4100 33876 4128
rect 29825 4091 29883 4097
rect 33870 4088 33876 4100
rect 33928 4088 33934 4140
rect 34057 4131 34115 4137
rect 34057 4097 34069 4131
rect 34103 4128 34115 4131
rect 34514 4128 34520 4140
rect 34103 4100 34520 4128
rect 34103 4097 34115 4100
rect 34057 4091 34115 4097
rect 34514 4088 34520 4100
rect 34572 4088 34578 4140
rect 35152 4131 35210 4137
rect 35152 4097 35164 4131
rect 35198 4128 35210 4131
rect 35434 4128 35440 4140
rect 35198 4100 35440 4128
rect 35198 4097 35210 4100
rect 35152 4091 35210 4097
rect 35434 4088 35440 4100
rect 35492 4088 35498 4140
rect 24903 4032 26234 4060
rect 24903 4029 24915 4032
rect 24857 4023 24915 4029
rect 24872 3992 24900 4023
rect 31110 4020 31116 4072
rect 31168 4060 31174 4072
rect 31754 4060 31760 4072
rect 31168 4032 31760 4060
rect 31168 4020 31174 4032
rect 31754 4020 31760 4032
rect 31812 4060 31818 4072
rect 34698 4060 34704 4072
rect 31812 4032 34704 4060
rect 31812 4020 31818 4032
rect 34698 4020 34704 4032
rect 34756 4060 34762 4072
rect 34885 4063 34943 4069
rect 34885 4060 34897 4063
rect 34756 4032 34897 4060
rect 34756 4020 34762 4032
rect 34885 4029 34897 4032
rect 34931 4029 34943 4063
rect 34885 4023 34943 4029
rect 23124 3964 24900 3992
rect 15712 3952 15718 3964
rect 4706 3924 4712 3936
rect 4667 3896 4712 3924
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 5445 3927 5503 3933
rect 5445 3893 5457 3927
rect 5491 3924 5503 3927
rect 5718 3924 5724 3936
rect 5491 3896 5724 3924
rect 5491 3893 5503 3896
rect 5445 3887 5503 3893
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 7742 3924 7748 3936
rect 7703 3896 7748 3924
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 10689 3927 10747 3933
rect 10689 3893 10701 3927
rect 10735 3924 10747 3927
rect 10870 3924 10876 3936
rect 10735 3896 10876 3924
rect 10735 3893 10747 3896
rect 10689 3887 10747 3893
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 13633 3927 13691 3933
rect 13633 3924 13645 3927
rect 13504 3896 13645 3924
rect 13504 3884 13510 3896
rect 13633 3893 13645 3896
rect 13679 3893 13691 3927
rect 17494 3924 17500 3936
rect 17455 3896 17500 3924
rect 13633 3887 13691 3893
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 19886 3884 19892 3936
rect 19944 3924 19950 3936
rect 19981 3927 20039 3933
rect 19981 3924 19993 3927
rect 19944 3896 19993 3924
rect 19944 3884 19950 3896
rect 19981 3893 19993 3896
rect 20027 3893 20039 3927
rect 19981 3887 20039 3893
rect 24489 3927 24547 3933
rect 24489 3893 24501 3927
rect 24535 3924 24547 3927
rect 24578 3924 24584 3936
rect 24535 3896 24584 3924
rect 24535 3893 24547 3896
rect 24489 3887 24547 3893
rect 24578 3884 24584 3896
rect 24636 3884 24642 3936
rect 27525 3927 27583 3933
rect 27525 3893 27537 3927
rect 27571 3924 27583 3927
rect 27614 3924 27620 3936
rect 27571 3896 27620 3924
rect 27571 3893 27583 3896
rect 27525 3887 27583 3893
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 34054 3924 34060 3936
rect 34015 3896 34060 3924
rect 34054 3884 34060 3896
rect 34112 3884 34118 3936
rect 36262 3924 36268 3936
rect 36223 3896 36268 3924
rect 36262 3884 36268 3896
rect 36320 3884 36326 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 2823 3692 11192 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 5169 3655 5227 3661
rect 5169 3621 5181 3655
rect 5215 3652 5227 3655
rect 6822 3652 6828 3664
rect 5215 3624 6828 3652
rect 5215 3621 5227 3624
rect 5169 3615 5227 3621
rect 6822 3612 6828 3624
rect 6880 3612 6886 3664
rect 9766 3652 9772 3664
rect 9727 3624 9772 3652
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 2041 3587 2099 3593
rect 2041 3584 2053 3587
rect 1412 3556 2053 3584
rect 1412 3528 1440 3556
rect 2041 3553 2053 3556
rect 2087 3553 2099 3587
rect 11164 3584 11192 3692
rect 11238 3680 11244 3732
rect 11296 3720 11302 3732
rect 15746 3720 15752 3732
rect 11296 3692 15752 3720
rect 11296 3680 11302 3692
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 16390 3720 16396 3732
rect 16351 3692 16396 3720
rect 16390 3680 16396 3692
rect 16448 3680 16454 3732
rect 19334 3720 19340 3732
rect 16868 3692 19340 3720
rect 15764 3652 15792 3680
rect 16868 3652 16896 3692
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 20990 3720 20996 3732
rect 20951 3692 20996 3720
rect 20990 3680 20996 3692
rect 21048 3680 21054 3732
rect 22922 3720 22928 3732
rect 22883 3692 22928 3720
rect 22922 3680 22928 3692
rect 22980 3680 22986 3732
rect 29638 3720 29644 3732
rect 27632 3692 29644 3720
rect 23750 3652 23756 3664
rect 15764 3624 16896 3652
rect 23400 3624 23756 3652
rect 13078 3584 13084 3596
rect 11164 3556 13084 3584
rect 2041 3547 2099 3553
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 23400 3593 23428 3624
rect 23750 3612 23756 3624
rect 23808 3652 23814 3664
rect 23808 3624 26234 3652
rect 23808 3612 23814 3624
rect 23385 3587 23443 3593
rect 23385 3553 23397 3587
rect 23431 3553 23443 3587
rect 23385 3547 23443 3553
rect 23474 3544 23480 3596
rect 23532 3584 23538 3596
rect 23532 3556 23577 3584
rect 23532 3544 23538 3556
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 1596 3488 2697 3516
rect 1596 3389 1624 3488
rect 2685 3485 2697 3488
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 2924 3488 3801 3516
rect 2924 3476 2930 3488
rect 3789 3485 3801 3488
rect 3835 3516 3847 3519
rect 3878 3516 3884 3528
rect 3835 3488 3884 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 3878 3476 3884 3488
rect 3936 3516 3942 3528
rect 5718 3516 5724 3528
rect 3936 3488 5724 3516
rect 3936 3476 3942 3488
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 10870 3476 10876 3528
rect 10928 3525 10934 3528
rect 10928 3516 10940 3525
rect 11149 3519 11207 3525
rect 10928 3488 10973 3516
rect 10928 3479 10940 3488
rect 11149 3485 11161 3519
rect 11195 3516 11207 3519
rect 11195 3488 11744 3516
rect 11195 3485 11207 3488
rect 11149 3479 11207 3485
rect 10928 3476 10934 3479
rect 4056 3451 4114 3457
rect 4056 3417 4068 3451
rect 4102 3448 4114 3451
rect 4706 3448 4712 3460
rect 4102 3420 4712 3448
rect 4102 3417 4114 3420
rect 4056 3411 4114 3417
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 11238 3448 11244 3460
rect 4816 3420 11244 3448
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 3970 3340 3976 3392
rect 4028 3380 4034 3392
rect 4816 3380 4844 3420
rect 11238 3408 11244 3420
rect 11296 3408 11302 3460
rect 11716 3392 11744 3488
rect 17494 3476 17500 3528
rect 17552 3525 17558 3528
rect 17552 3516 17564 3525
rect 17770 3516 17776 3528
rect 17552 3488 17597 3516
rect 17731 3488 17776 3516
rect 17552 3479 17564 3488
rect 17552 3476 17558 3479
rect 17770 3476 17776 3488
rect 17828 3516 17834 3528
rect 19886 3525 19892 3528
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 17828 3488 18245 3516
rect 17828 3476 17834 3488
rect 18233 3485 18245 3488
rect 18279 3516 18291 3519
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 18279 3488 19625 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 19613 3485 19625 3488
rect 19659 3485 19671 3519
rect 19880 3516 19892 3525
rect 19847 3488 19892 3516
rect 19613 3479 19671 3485
rect 19880 3479 19892 3488
rect 19886 3476 19892 3479
rect 19944 3476 19950 3528
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 26206 3516 26234 3624
rect 27632 3593 27660 3692
rect 29638 3680 29644 3692
rect 29696 3720 29702 3732
rect 30561 3723 30619 3729
rect 30561 3720 30573 3723
rect 29696 3692 30573 3720
rect 29696 3680 29702 3692
rect 30561 3689 30573 3692
rect 30607 3689 30619 3723
rect 32490 3720 32496 3732
rect 32451 3692 32496 3720
rect 30561 3683 30619 3689
rect 28997 3655 29055 3661
rect 28997 3621 29009 3655
rect 29043 3652 29055 3655
rect 29270 3652 29276 3664
rect 29043 3624 29276 3652
rect 29043 3621 29055 3624
rect 28997 3615 29055 3621
rect 29270 3612 29276 3624
rect 29328 3612 29334 3664
rect 27617 3587 27675 3593
rect 27617 3553 27629 3587
rect 27663 3553 27675 3587
rect 30576 3584 30604 3683
rect 32490 3680 32496 3692
rect 32548 3720 32554 3732
rect 34606 3720 34612 3732
rect 32548 3692 34612 3720
rect 32548 3680 32554 3692
rect 34606 3680 34612 3692
rect 34664 3680 34670 3732
rect 35161 3723 35219 3729
rect 35161 3689 35173 3723
rect 35207 3720 35219 3723
rect 35434 3720 35440 3732
rect 35207 3692 35440 3720
rect 35207 3689 35219 3692
rect 35161 3683 35219 3689
rect 35434 3680 35440 3692
rect 35492 3680 35498 3732
rect 31110 3584 31116 3596
rect 30576 3556 31116 3584
rect 27617 3547 27675 3553
rect 31110 3544 31116 3556
rect 31168 3544 31174 3596
rect 36262 3584 36268 3596
rect 34900 3556 36268 3584
rect 34900 3516 34928 3556
rect 36262 3544 36268 3556
rect 36320 3544 36326 3596
rect 26206 3488 34928 3516
rect 34977 3519 35035 3525
rect 34977 3485 34989 3519
rect 35023 3485 35035 3519
rect 34977 3479 35035 3485
rect 35161 3519 35219 3525
rect 35161 3485 35173 3519
rect 35207 3516 35219 3519
rect 35802 3516 35808 3528
rect 35207 3488 35808 3516
rect 35207 3485 35219 3488
rect 35161 3479 35219 3485
rect 23293 3451 23351 3457
rect 23293 3417 23305 3451
rect 23339 3448 23351 3451
rect 23658 3448 23664 3460
rect 23339 3420 23664 3448
rect 23339 3417 23351 3420
rect 23293 3411 23351 3417
rect 23658 3408 23664 3420
rect 23716 3448 23722 3460
rect 27890 3457 27896 3460
rect 23716 3420 26234 3448
rect 23716 3408 23722 3420
rect 5718 3380 5724 3392
rect 4028 3352 4844 3380
rect 5679 3352 5724 3380
rect 4028 3340 4034 3352
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 11698 3380 11704 3392
rect 11659 3352 11704 3380
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 24394 3380 24400 3392
rect 24355 3352 24400 3380
rect 24394 3340 24400 3352
rect 24452 3340 24458 3392
rect 26206 3380 26234 3420
rect 27884 3411 27896 3457
rect 27948 3448 27954 3460
rect 27948 3420 27984 3448
rect 27890 3408 27896 3411
rect 27948 3408 27954 3420
rect 31202 3408 31208 3460
rect 31260 3448 31266 3460
rect 31358 3451 31416 3457
rect 31358 3448 31370 3451
rect 31260 3420 31370 3448
rect 31260 3408 31266 3420
rect 31358 3417 31370 3420
rect 31404 3417 31416 3451
rect 34698 3448 34704 3460
rect 31358 3411 31416 3417
rect 31726 3420 34704 3448
rect 31726 3380 31754 3420
rect 34698 3408 34704 3420
rect 34756 3408 34762 3460
rect 26206 3352 31754 3380
rect 33870 3340 33876 3392
rect 33928 3380 33934 3392
rect 34992 3380 35020 3479
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 33928 3352 35020 3380
rect 33928 3340 33934 3352
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 8849 3179 8907 3185
rect 8849 3145 8861 3179
rect 8895 3176 8907 3179
rect 9306 3176 9312 3188
rect 8895 3148 9312 3176
rect 8895 3145 8907 3148
rect 8849 3139 8907 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 14550 3176 14556 3188
rect 14511 3148 14556 3176
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 22833 3179 22891 3185
rect 22833 3176 22845 3179
rect 22066 3148 22845 3176
rect 5718 3068 5724 3120
rect 5776 3108 5782 3120
rect 9493 3111 9551 3117
rect 9493 3108 9505 3111
rect 5776 3080 9505 3108
rect 5776 3068 5782 3080
rect 7484 3049 7512 3080
rect 9493 3077 9505 3080
rect 9539 3108 9551 3111
rect 11698 3108 11704 3120
rect 9539 3080 11704 3108
rect 9539 3077 9551 3080
rect 9493 3071 9551 3077
rect 11698 3068 11704 3080
rect 11756 3108 11762 3120
rect 15013 3111 15071 3117
rect 15013 3108 15025 3111
rect 11756 3080 15025 3108
rect 11756 3068 11762 3080
rect 7742 3049 7748 3052
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 7469 3043 7527 3049
rect 1719 3012 3740 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 1489 2907 1547 2913
rect 1489 2873 1501 2907
rect 1535 2904 1547 2907
rect 2774 2904 2780 2916
rect 1535 2876 2780 2904
rect 1535 2873 1547 2876
rect 1489 2867 1547 2873
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 2593 2839 2651 2845
rect 2593 2805 2605 2839
rect 2639 2836 2651 2839
rect 2682 2836 2688 2848
rect 2639 2808 2688 2836
rect 2639 2805 2651 2808
rect 2593 2799 2651 2805
rect 2682 2796 2688 2808
rect 2740 2796 2746 2848
rect 2958 2796 2964 2848
rect 3016 2836 3022 2848
rect 3712 2845 3740 3012
rect 7469 3009 7481 3043
rect 7515 3009 7527 3043
rect 7736 3040 7748 3049
rect 7703 3012 7748 3040
rect 7469 3003 7527 3009
rect 7736 3003 7748 3012
rect 7742 3000 7748 3003
rect 7800 3000 7806 3052
rect 13188 3049 13216 3080
rect 15013 3077 15025 3080
rect 15059 3108 15071 3111
rect 16666 3108 16672 3120
rect 15059 3080 16672 3108
rect 15059 3077 15071 3080
rect 15013 3071 15071 3077
rect 16666 3068 16672 3080
rect 16724 3108 16730 3120
rect 17770 3108 17776 3120
rect 16724 3080 17776 3108
rect 16724 3068 16730 3080
rect 17770 3068 17776 3080
rect 17828 3108 17834 3120
rect 19429 3111 19487 3117
rect 19429 3108 19441 3111
rect 17828 3080 19441 3108
rect 17828 3068 17834 3080
rect 19429 3077 19441 3080
rect 19475 3108 19487 3111
rect 20898 3108 20904 3120
rect 19475 3080 20904 3108
rect 19475 3077 19487 3080
rect 19429 3071 19487 3077
rect 20898 3068 20904 3080
rect 20956 3108 20962 3120
rect 22066 3108 22094 3148
rect 22833 3145 22845 3148
rect 22879 3145 22891 3179
rect 22833 3139 22891 3145
rect 20956 3080 22094 3108
rect 20956 3068 20962 3080
rect 13446 3049 13452 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3009 13231 3043
rect 13440 3040 13452 3049
rect 13407 3012 13452 3040
rect 13173 3003 13231 3009
rect 13440 3003 13452 3012
rect 13446 3000 13452 3003
rect 13504 3000 13510 3052
rect 22848 3040 22876 3139
rect 23474 3136 23480 3188
rect 23532 3176 23538 3188
rect 24765 3179 24823 3185
rect 24765 3176 24777 3179
rect 23532 3148 24777 3176
rect 23532 3136 23538 3148
rect 24765 3145 24777 3148
rect 24811 3145 24823 3179
rect 24765 3139 24823 3145
rect 27801 3179 27859 3185
rect 27801 3145 27813 3179
rect 27847 3176 27859 3179
rect 27890 3176 27896 3188
rect 27847 3148 27896 3176
rect 27847 3145 27859 3148
rect 27801 3139 27859 3145
rect 27890 3136 27896 3148
rect 27948 3136 27954 3188
rect 31110 3136 31116 3188
rect 31168 3176 31174 3188
rect 32769 3179 32827 3185
rect 32769 3176 32781 3179
rect 31168 3148 32781 3176
rect 31168 3136 31174 3148
rect 32769 3145 32781 3148
rect 32815 3145 32827 3179
rect 34698 3176 34704 3188
rect 34659 3148 34704 3176
rect 32769 3139 32827 3145
rect 23652 3111 23710 3117
rect 23652 3077 23664 3111
rect 23698 3108 23710 3111
rect 24394 3108 24400 3120
rect 23698 3080 24400 3108
rect 23698 3077 23710 3080
rect 23652 3071 23710 3077
rect 24394 3068 24400 3080
rect 24452 3068 24458 3120
rect 31386 3108 31392 3120
rect 26206 3080 31392 3108
rect 23385 3043 23443 3049
rect 23385 3040 23397 3043
rect 22848 3012 23397 3040
rect 23385 3009 23397 3012
rect 23431 3009 23443 3043
rect 26206 3040 26234 3080
rect 31386 3068 31392 3080
rect 31444 3068 31450 3120
rect 27614 3040 27620 3052
rect 23385 3003 23443 3009
rect 23492 3012 26234 3040
rect 27575 3012 27620 3040
rect 23492 2972 23520 3012
rect 27614 3000 27620 3012
rect 27672 3000 27678 3052
rect 32784 3040 32812 3139
rect 34698 3136 34704 3148
rect 34756 3136 34762 3188
rect 33588 3111 33646 3117
rect 33588 3077 33600 3111
rect 33634 3108 33646 3111
rect 34054 3108 34060 3120
rect 33634 3080 34060 3108
rect 33634 3077 33646 3080
rect 33588 3071 33646 3077
rect 34054 3068 34060 3080
rect 34112 3068 34118 3120
rect 33321 3043 33379 3049
rect 33321 3040 33333 3043
rect 32784 3012 33333 3040
rect 33321 3009 33333 3012
rect 33367 3009 33379 3043
rect 33321 3003 33379 3009
rect 22066 2944 23520 2972
rect 22066 2904 22094 2944
rect 8404 2876 12434 2904
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 3016 2808 3065 2836
rect 3016 2796 3022 2808
rect 3053 2805 3065 2808
rect 3099 2805 3111 2839
rect 3053 2799 3111 2805
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 8404 2836 8432 2876
rect 3743 2808 8432 2836
rect 12406 2836 12434 2876
rect 14476 2876 22094 2904
rect 14476 2836 14504 2876
rect 12406 2808 14504 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 3050 2632 3056 2644
rect 2915 2604 3056 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 2958 2496 2964 2508
rect 1872 2468 2964 2496
rect 1872 2372 1900 2468
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 2682 2428 2688 2440
rect 2643 2400 2688 2428
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 34606 2388 34612 2440
rect 34664 2428 34670 2440
rect 37829 2431 37887 2437
rect 37829 2428 37841 2431
rect 34664 2400 37841 2428
rect 34664 2388 34670 2400
rect 37829 2397 37841 2400
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 2225 2363 2283 2369
rect 2225 2329 2237 2363
rect 2271 2360 2283 2363
rect 13354 2360 13360 2372
rect 2271 2332 13360 2360
rect 2271 2329 2283 2332
rect 2225 2323 2283 2329
rect 13354 2320 13360 2332
rect 13412 2320 13418 2372
rect 38010 2292 38016 2304
rect 37971 2264 38016 2292
rect 38010 2252 38016 2264
rect 38068 2252 38074 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 38016 37451 38068 37460
rect 38016 37417 38025 37451
rect 38025 37417 38059 37451
rect 38059 37417 38068 37451
rect 38016 37408 38068 37417
rect 29920 37204 29972 37256
rect 37832 37247 37884 37256
rect 37832 37213 37841 37247
rect 37841 37213 37875 37247
rect 37875 37213 37884 37247
rect 37832 37204 37884 37213
rect 30196 37111 30248 37120
rect 30196 37077 30205 37111
rect 30205 37077 30239 37111
rect 30239 37077 30248 37111
rect 30196 37068 30248 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 29920 36907 29972 36916
rect 29920 36873 29929 36907
rect 29929 36873 29963 36907
rect 29963 36873 29972 36907
rect 29920 36864 29972 36873
rect 3976 36796 4028 36848
rect 12348 36771 12400 36780
rect 12348 36737 12357 36771
rect 12357 36737 12391 36771
rect 12391 36737 12400 36771
rect 12348 36728 12400 36737
rect 16396 36660 16448 36712
rect 17500 36703 17552 36712
rect 17500 36669 17509 36703
rect 17509 36669 17543 36703
rect 17543 36669 17552 36703
rect 17500 36660 17552 36669
rect 17960 36660 18012 36712
rect 18052 36703 18104 36712
rect 18052 36669 18061 36703
rect 18061 36669 18095 36703
rect 18095 36669 18104 36703
rect 18052 36660 18104 36669
rect 4068 36592 4120 36644
rect 15200 36592 15252 36644
rect 24584 36703 24636 36712
rect 24584 36669 24593 36703
rect 24593 36669 24627 36703
rect 24627 36669 24636 36703
rect 24584 36660 24636 36669
rect 24768 36703 24820 36712
rect 24768 36669 24777 36703
rect 24777 36669 24811 36703
rect 24811 36669 24820 36703
rect 24768 36660 24820 36669
rect 27620 36592 27672 36644
rect 3148 36567 3200 36576
rect 3148 36533 3157 36567
rect 3157 36533 3191 36567
rect 3191 36533 3200 36567
rect 3148 36524 3200 36533
rect 3884 36567 3936 36576
rect 3884 36533 3893 36567
rect 3893 36533 3927 36567
rect 3927 36533 3936 36567
rect 3884 36524 3936 36533
rect 4712 36567 4764 36576
rect 4712 36533 4721 36567
rect 4721 36533 4755 36567
rect 4755 36533 4764 36567
rect 4712 36524 4764 36533
rect 8944 36524 8996 36576
rect 9128 36567 9180 36576
rect 9128 36533 9137 36567
rect 9137 36533 9171 36567
rect 9171 36533 9180 36567
rect 9128 36524 9180 36533
rect 12624 36524 12676 36576
rect 19432 36524 19484 36576
rect 26608 36524 26660 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 12532 36363 12584 36372
rect 12532 36329 12541 36363
rect 12541 36329 12575 36363
rect 12575 36329 12584 36363
rect 12532 36320 12584 36329
rect 17500 36363 17552 36372
rect 17500 36329 17509 36363
rect 17509 36329 17543 36363
rect 17543 36329 17552 36363
rect 17500 36320 17552 36329
rect 17960 36363 18012 36372
rect 17960 36329 17969 36363
rect 17969 36329 18003 36363
rect 18003 36329 18012 36363
rect 17960 36320 18012 36329
rect 24584 36320 24636 36372
rect 3792 36252 3844 36304
rect 5264 36227 5316 36236
rect 5264 36193 5273 36227
rect 5273 36193 5307 36227
rect 5307 36193 5316 36227
rect 5264 36184 5316 36193
rect 8944 36227 8996 36236
rect 8944 36193 8953 36227
rect 8953 36193 8987 36227
rect 8987 36193 8996 36227
rect 8944 36184 8996 36193
rect 9772 36227 9824 36236
rect 9772 36193 9781 36227
rect 9781 36193 9815 36227
rect 9815 36193 9824 36227
rect 9772 36184 9824 36193
rect 12440 36184 12492 36236
rect 13820 36184 13872 36236
rect 19432 36227 19484 36236
rect 19432 36193 19441 36227
rect 19441 36193 19475 36227
rect 19475 36193 19484 36227
rect 19432 36184 19484 36193
rect 20904 36227 20956 36236
rect 20904 36193 20913 36227
rect 20913 36193 20947 36227
rect 20947 36193 20956 36227
rect 20904 36184 20956 36193
rect 23572 36184 23624 36236
rect 26608 36227 26660 36236
rect 26608 36193 26617 36227
rect 26617 36193 26651 36227
rect 26651 36193 26660 36227
rect 26608 36184 26660 36193
rect 27620 36227 27672 36236
rect 27620 36193 27629 36227
rect 27629 36193 27663 36227
rect 27663 36193 27672 36227
rect 27620 36184 27672 36193
rect 7564 36116 7616 36168
rect 12808 36116 12860 36168
rect 3332 36048 3384 36100
rect 11980 36048 12032 36100
rect 12716 35980 12768 36032
rect 14096 36159 14148 36168
rect 14096 36125 14105 36159
rect 14105 36125 14139 36159
rect 14139 36125 14148 36159
rect 14096 36116 14148 36125
rect 16028 36159 16080 36168
rect 16028 36125 16037 36159
rect 16037 36125 16071 36159
rect 16071 36125 16080 36159
rect 16028 36116 16080 36125
rect 18144 36159 18196 36168
rect 18144 36125 18153 36159
rect 18153 36125 18187 36159
rect 18187 36125 18196 36159
rect 18144 36116 18196 36125
rect 21732 36159 21784 36168
rect 21732 36125 21741 36159
rect 21741 36125 21775 36159
rect 21775 36125 21784 36159
rect 21732 36116 21784 36125
rect 24308 36116 24360 36168
rect 26148 36159 26200 36168
rect 26148 36125 26157 36159
rect 26157 36125 26191 36159
rect 26191 36125 26200 36159
rect 26148 36116 26200 36125
rect 21916 36091 21968 36100
rect 13544 36023 13596 36032
rect 13544 35989 13553 36023
rect 13553 35989 13587 36023
rect 13587 35989 13596 36023
rect 13544 35980 13596 35989
rect 19432 35980 19484 36032
rect 21916 36057 21925 36091
rect 21925 36057 21959 36091
rect 21959 36057 21968 36091
rect 21916 36048 21968 36057
rect 26792 36091 26844 36100
rect 26792 36057 26801 36091
rect 26801 36057 26835 36091
rect 26835 36057 26844 36091
rect 26792 36048 26844 36057
rect 20904 35980 20956 36032
rect 25596 35980 25648 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 5264 35751 5316 35760
rect 5264 35717 5273 35751
rect 5273 35717 5307 35751
rect 5307 35717 5316 35751
rect 5264 35708 5316 35717
rect 16856 35776 16908 35828
rect 19432 35776 19484 35828
rect 21916 35776 21968 35828
rect 12624 35751 12676 35760
rect 12624 35717 12633 35751
rect 12633 35717 12667 35751
rect 12667 35717 12676 35751
rect 12624 35708 12676 35717
rect 15200 35708 15252 35760
rect 20904 35708 20956 35760
rect 7564 35683 7616 35692
rect 7564 35649 7573 35683
rect 7573 35649 7607 35683
rect 7607 35649 7616 35683
rect 7564 35640 7616 35649
rect 11520 35640 11572 35692
rect 12440 35683 12492 35692
rect 3792 35572 3844 35624
rect 8024 35572 8076 35624
rect 9772 35572 9824 35624
rect 11888 35615 11940 35624
rect 11888 35581 11897 35615
rect 11897 35581 11931 35615
rect 11931 35581 11940 35615
rect 11888 35572 11940 35581
rect 12440 35649 12449 35683
rect 12449 35649 12483 35683
rect 12483 35649 12492 35683
rect 12440 35640 12492 35649
rect 15936 35683 15988 35692
rect 15936 35649 15945 35683
rect 15945 35649 15979 35683
rect 15979 35649 15988 35683
rect 15936 35640 15988 35649
rect 16028 35640 16080 35692
rect 18972 35640 19024 35692
rect 20628 35683 20680 35692
rect 20628 35649 20637 35683
rect 20637 35649 20671 35683
rect 20671 35649 20680 35683
rect 20628 35640 20680 35649
rect 21732 35640 21784 35692
rect 29552 35640 29604 35692
rect 30288 35683 30340 35692
rect 30288 35649 30322 35683
rect 30322 35649 30340 35683
rect 30288 35640 30340 35649
rect 32220 35640 32272 35692
rect 12808 35572 12860 35624
rect 18236 35615 18288 35624
rect 4068 35504 4120 35556
rect 9312 35436 9364 35488
rect 10140 35436 10192 35488
rect 12532 35436 12584 35488
rect 18236 35581 18245 35615
rect 18245 35581 18279 35615
rect 18279 35581 18288 35615
rect 18236 35572 18288 35581
rect 23112 35615 23164 35624
rect 23112 35581 23121 35615
rect 23121 35581 23155 35615
rect 23155 35581 23164 35615
rect 23112 35572 23164 35581
rect 23296 35615 23348 35624
rect 23296 35581 23305 35615
rect 23305 35581 23339 35615
rect 23339 35581 23348 35615
rect 23296 35572 23348 35581
rect 23756 35615 23808 35624
rect 23756 35581 23765 35615
rect 23765 35581 23799 35615
rect 23799 35581 23808 35615
rect 23756 35572 23808 35581
rect 27160 35615 27212 35624
rect 27160 35581 27169 35615
rect 27169 35581 27203 35615
rect 27203 35581 27212 35615
rect 27160 35572 27212 35581
rect 27620 35572 27672 35624
rect 28356 35615 28408 35624
rect 28356 35581 28365 35615
rect 28365 35581 28399 35615
rect 28399 35581 28408 35615
rect 28356 35572 28408 35581
rect 32128 35615 32180 35624
rect 32128 35581 32137 35615
rect 32137 35581 32171 35615
rect 32171 35581 32180 35615
rect 32128 35572 32180 35581
rect 14280 35436 14332 35488
rect 18052 35436 18104 35488
rect 18328 35436 18380 35488
rect 21916 35436 21968 35488
rect 29920 35436 29972 35488
rect 33508 35479 33560 35488
rect 33508 35445 33517 35479
rect 33517 35445 33551 35479
rect 33551 35445 33560 35479
rect 33508 35436 33560 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3332 35232 3384 35284
rect 3792 35275 3844 35284
rect 3792 35241 3801 35275
rect 3801 35241 3835 35275
rect 3835 35241 3844 35275
rect 3792 35232 3844 35241
rect 8024 35275 8076 35284
rect 8024 35241 8033 35275
rect 8033 35241 8067 35275
rect 8067 35241 8076 35275
rect 8024 35232 8076 35241
rect 12348 35232 12400 35284
rect 16396 35275 16448 35284
rect 10140 35164 10192 35216
rect 12532 35164 12584 35216
rect 16396 35241 16405 35275
rect 16405 35241 16439 35275
rect 16439 35241 16448 35275
rect 16396 35232 16448 35241
rect 17776 35275 17828 35284
rect 17776 35241 17785 35275
rect 17785 35241 17819 35275
rect 17819 35241 17828 35275
rect 17776 35232 17828 35241
rect 20628 35232 20680 35284
rect 26792 35232 26844 35284
rect 32220 35232 32272 35284
rect 6000 35096 6052 35148
rect 9128 35139 9180 35148
rect 9128 35105 9137 35139
rect 9137 35105 9171 35139
rect 9171 35105 9180 35139
rect 9128 35096 9180 35105
rect 9312 35139 9364 35148
rect 9312 35105 9321 35139
rect 9321 35105 9355 35139
rect 9355 35105 9364 35139
rect 9312 35096 9364 35105
rect 11980 35139 12032 35148
rect 6736 35071 6788 35080
rect 4344 34960 4396 35012
rect 4712 34960 4764 35012
rect 6736 35037 6745 35071
rect 6745 35037 6779 35071
rect 6779 35037 6788 35071
rect 6736 35028 6788 35037
rect 8116 35028 8168 35080
rect 11980 35105 11989 35139
rect 11989 35105 12023 35139
rect 12023 35105 12032 35139
rect 11980 35096 12032 35105
rect 13820 35164 13872 35216
rect 14648 35164 14700 35216
rect 12440 35028 12492 35080
rect 4068 34892 4120 34944
rect 11796 34960 11848 35012
rect 14096 35139 14148 35148
rect 14096 35105 14105 35139
rect 14105 35105 14139 35139
rect 14139 35105 14148 35139
rect 14096 35096 14148 35105
rect 15200 35139 15252 35148
rect 15200 35105 15209 35139
rect 15209 35105 15243 35139
rect 15243 35105 15252 35139
rect 15200 35096 15252 35105
rect 17960 35139 18012 35148
rect 12808 35028 12860 35080
rect 16580 35071 16632 35080
rect 16580 35037 16589 35071
rect 16589 35037 16623 35071
rect 16623 35037 16632 35071
rect 16580 35028 16632 35037
rect 16672 35071 16724 35080
rect 16672 35037 16681 35071
rect 16681 35037 16715 35071
rect 16715 35037 16724 35071
rect 16672 35028 16724 35037
rect 16856 35071 16908 35080
rect 16856 35037 16865 35071
rect 16865 35037 16899 35071
rect 16899 35037 16908 35071
rect 17960 35105 17969 35139
rect 17969 35105 18003 35139
rect 18003 35105 18012 35139
rect 17960 35096 18012 35105
rect 21916 35139 21968 35148
rect 21916 35105 21925 35139
rect 21925 35105 21959 35139
rect 21959 35105 21968 35139
rect 21916 35096 21968 35105
rect 23756 35139 23808 35148
rect 23756 35105 23765 35139
rect 23765 35105 23799 35139
rect 23799 35105 23808 35139
rect 23756 35096 23808 35105
rect 24584 35096 24636 35148
rect 24768 35096 24820 35148
rect 26148 35096 26200 35148
rect 28356 35139 28408 35148
rect 28356 35105 28365 35139
rect 28365 35105 28399 35139
rect 28399 35105 28408 35139
rect 28356 35096 28408 35105
rect 29552 35139 29604 35148
rect 29552 35105 29561 35139
rect 29561 35105 29595 35139
rect 29595 35105 29604 35139
rect 29552 35096 29604 35105
rect 16856 35028 16908 35037
rect 17868 35028 17920 35080
rect 18788 35028 18840 35080
rect 23480 35028 23532 35080
rect 25872 35071 25924 35080
rect 25872 35037 25881 35071
rect 25881 35037 25915 35071
rect 25915 35037 25924 35071
rect 25872 35028 25924 35037
rect 31944 35071 31996 35080
rect 31944 35037 31953 35071
rect 31953 35037 31987 35071
rect 31987 35037 31996 35071
rect 31944 35028 31996 35037
rect 12716 34960 12768 35012
rect 13544 34960 13596 35012
rect 17316 34960 17368 35012
rect 21180 34960 21232 35012
rect 26884 35003 26936 35012
rect 26884 34969 26893 35003
rect 26893 34969 26927 35003
rect 26927 34969 26936 35003
rect 26884 34960 26936 34969
rect 29828 35003 29880 35012
rect 29828 34969 29862 35003
rect 29862 34969 29880 35003
rect 29828 34960 29880 34969
rect 18236 34892 18288 34944
rect 30104 34892 30156 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 6736 34731 6788 34740
rect 6736 34697 6745 34731
rect 6745 34697 6779 34731
rect 6779 34697 6788 34731
rect 6736 34688 6788 34697
rect 8116 34731 8168 34740
rect 8116 34697 8125 34731
rect 8125 34697 8159 34731
rect 8159 34697 8168 34731
rect 8116 34688 8168 34697
rect 11520 34731 11572 34740
rect 11520 34697 11529 34731
rect 11529 34697 11563 34731
rect 11563 34697 11572 34731
rect 11520 34688 11572 34697
rect 12440 34731 12492 34740
rect 12440 34697 12449 34731
rect 12449 34697 12483 34731
rect 12483 34697 12492 34731
rect 12440 34688 12492 34697
rect 3884 34620 3936 34672
rect 8024 34620 8076 34672
rect 3148 34595 3200 34604
rect 3148 34561 3157 34595
rect 3157 34561 3191 34595
rect 3191 34561 3200 34595
rect 3148 34552 3200 34561
rect 7472 34552 7524 34604
rect 11796 34595 11848 34604
rect 11796 34561 11805 34595
rect 11805 34561 11839 34595
rect 11839 34561 11848 34595
rect 11796 34552 11848 34561
rect 11980 34595 12032 34604
rect 11980 34561 11989 34595
rect 11989 34561 12023 34595
rect 12023 34561 12032 34595
rect 12808 34620 12860 34672
rect 15936 34688 15988 34740
rect 16856 34688 16908 34740
rect 18052 34731 18104 34740
rect 18052 34697 18061 34731
rect 18061 34697 18095 34731
rect 18095 34697 18104 34731
rect 18972 34731 19024 34740
rect 18052 34688 18104 34697
rect 18972 34697 18981 34731
rect 18981 34697 19015 34731
rect 19015 34697 19024 34731
rect 18972 34688 19024 34697
rect 21180 34731 21232 34740
rect 21180 34697 21189 34731
rect 21189 34697 21223 34731
rect 21223 34697 21232 34731
rect 21180 34688 21232 34697
rect 29828 34731 29880 34740
rect 29828 34697 29837 34731
rect 29837 34697 29871 34731
rect 29871 34697 29880 34731
rect 29828 34688 29880 34697
rect 30288 34731 30340 34740
rect 30288 34697 30297 34731
rect 30297 34697 30331 34731
rect 30331 34697 30340 34731
rect 30288 34688 30340 34697
rect 11980 34552 12032 34561
rect 12900 34595 12952 34604
rect 12900 34561 12909 34595
rect 12909 34561 12943 34595
rect 12943 34561 12952 34595
rect 12900 34552 12952 34561
rect 13544 34595 13596 34604
rect 13544 34561 13553 34595
rect 13553 34561 13587 34595
rect 13587 34561 13596 34595
rect 15936 34595 15988 34604
rect 13544 34552 13596 34561
rect 15936 34561 15945 34595
rect 15945 34561 15979 34595
rect 15979 34561 15988 34595
rect 15936 34552 15988 34561
rect 16120 34552 16172 34604
rect 16580 34552 16632 34604
rect 32128 34620 32180 34672
rect 4344 34527 4396 34536
rect 4344 34493 4353 34527
rect 4353 34493 4387 34527
rect 4387 34493 4396 34527
rect 4344 34484 4396 34493
rect 4620 34484 4672 34536
rect 4068 34416 4120 34468
rect 11888 34484 11940 34536
rect 16672 34484 16724 34536
rect 16948 34527 17000 34536
rect 16948 34493 16957 34527
rect 16957 34493 16991 34527
rect 16991 34493 17000 34527
rect 16948 34484 17000 34493
rect 17684 34527 17736 34536
rect 17684 34493 17693 34527
rect 17693 34493 17727 34527
rect 17727 34493 17736 34527
rect 17684 34484 17736 34493
rect 17868 34595 17920 34604
rect 17868 34561 17893 34595
rect 17893 34561 17920 34595
rect 17868 34552 17920 34561
rect 18052 34484 18104 34536
rect 18144 34484 18196 34536
rect 18788 34595 18840 34604
rect 18788 34561 18797 34595
rect 18797 34561 18831 34595
rect 18831 34561 18840 34595
rect 18788 34552 18840 34561
rect 20168 34552 20220 34604
rect 24308 34595 24360 34604
rect 24308 34561 24317 34595
rect 24317 34561 24351 34595
rect 24351 34561 24360 34595
rect 24308 34552 24360 34561
rect 29644 34595 29696 34604
rect 29644 34561 29653 34595
rect 29653 34561 29687 34595
rect 29687 34561 29696 34595
rect 29644 34552 29696 34561
rect 30472 34595 30524 34604
rect 30472 34561 30481 34595
rect 30481 34561 30515 34595
rect 30515 34561 30524 34595
rect 30472 34552 30524 34561
rect 34796 34620 34848 34672
rect 33232 34595 33284 34604
rect 33232 34561 33266 34595
rect 33266 34561 33284 34595
rect 33232 34552 33284 34561
rect 18604 34527 18656 34536
rect 18604 34493 18613 34527
rect 18613 34493 18647 34527
rect 18647 34493 18656 34527
rect 18604 34484 18656 34493
rect 21824 34527 21876 34536
rect 21824 34493 21833 34527
rect 21833 34493 21867 34527
rect 21867 34493 21876 34527
rect 21824 34484 21876 34493
rect 22008 34527 22060 34536
rect 22008 34493 22017 34527
rect 22017 34493 22051 34527
rect 22051 34493 22060 34527
rect 22008 34484 22060 34493
rect 24492 34527 24544 34536
rect 2780 34348 2832 34400
rect 3700 34348 3752 34400
rect 6276 34348 6328 34400
rect 7656 34391 7708 34400
rect 7656 34357 7665 34391
rect 7665 34357 7699 34391
rect 7699 34357 7708 34391
rect 7656 34348 7708 34357
rect 7932 34416 7984 34468
rect 14464 34416 14516 34468
rect 18420 34416 18472 34468
rect 24492 34493 24501 34527
rect 24501 34493 24535 34527
rect 24535 34493 24544 34527
rect 24492 34484 24544 34493
rect 24584 34484 24636 34536
rect 23664 34416 23716 34468
rect 12532 34348 12584 34400
rect 16120 34391 16172 34400
rect 16120 34357 16129 34391
rect 16129 34357 16163 34391
rect 16163 34357 16172 34391
rect 16120 34348 16172 34357
rect 17132 34391 17184 34400
rect 17132 34357 17141 34391
rect 17141 34357 17175 34391
rect 17175 34357 17184 34391
rect 17132 34348 17184 34357
rect 17776 34348 17828 34400
rect 19340 34348 19392 34400
rect 34336 34391 34388 34400
rect 34336 34357 34345 34391
rect 34345 34357 34379 34391
rect 34379 34357 34388 34391
rect 34336 34348 34388 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 6000 34144 6052 34196
rect 7748 34187 7800 34196
rect 7748 34153 7757 34187
rect 7757 34153 7791 34187
rect 7791 34153 7800 34187
rect 7748 34144 7800 34153
rect 12532 34144 12584 34196
rect 18604 34144 18656 34196
rect 21824 34187 21876 34196
rect 21824 34153 21833 34187
rect 21833 34153 21867 34187
rect 21867 34153 21876 34187
rect 21824 34144 21876 34153
rect 23112 34144 23164 34196
rect 29644 34144 29696 34196
rect 30472 34144 30524 34196
rect 31944 34144 31996 34196
rect 33232 34144 33284 34196
rect 17132 34076 17184 34128
rect 4620 34051 4672 34060
rect 4620 34017 4629 34051
rect 4629 34017 4663 34051
rect 4663 34017 4672 34051
rect 4620 34008 4672 34017
rect 6276 34051 6328 34060
rect 6276 34017 6285 34051
rect 6285 34017 6319 34051
rect 6319 34017 6328 34051
rect 6276 34008 6328 34017
rect 7932 34008 7984 34060
rect 16212 34008 16264 34060
rect 17960 34008 18012 34060
rect 18788 34008 18840 34060
rect 22008 34076 22060 34128
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 7472 33983 7524 33992
rect 7472 33949 7481 33983
rect 7481 33949 7515 33983
rect 7515 33949 7524 33983
rect 7472 33940 7524 33949
rect 12348 33983 12400 33992
rect 6092 33915 6144 33924
rect 6092 33881 6101 33915
rect 6101 33881 6135 33915
rect 6135 33881 6144 33915
rect 6092 33872 6144 33881
rect 8024 33872 8076 33924
rect 2688 33804 2740 33856
rect 11152 33847 11204 33856
rect 11152 33813 11161 33847
rect 11161 33813 11195 33847
rect 11195 33813 11204 33847
rect 11152 33804 11204 33813
rect 12348 33949 12357 33983
rect 12357 33949 12391 33983
rect 12391 33949 12400 33983
rect 12348 33940 12400 33949
rect 15660 33940 15712 33992
rect 17224 33940 17276 33992
rect 12716 33872 12768 33924
rect 17316 33915 17368 33924
rect 17316 33881 17325 33915
rect 17325 33881 17359 33915
rect 17359 33881 17368 33915
rect 17316 33872 17368 33881
rect 19340 33872 19392 33924
rect 13268 33804 13320 33856
rect 13544 33804 13596 33856
rect 16672 33804 16724 33856
rect 24492 34008 24544 34060
rect 26884 34008 26936 34060
rect 31576 34008 31628 34060
rect 24400 33940 24452 33992
rect 26056 33983 26108 33992
rect 26056 33949 26065 33983
rect 26065 33949 26099 33983
rect 26099 33949 26108 33983
rect 26056 33940 26108 33949
rect 27160 33940 27212 33992
rect 25872 33872 25924 33924
rect 23480 33804 23532 33856
rect 23572 33804 23624 33856
rect 29000 33940 29052 33992
rect 30748 33983 30800 33992
rect 30748 33949 30757 33983
rect 30757 33949 30791 33983
rect 30791 33949 30800 33983
rect 30748 33940 30800 33949
rect 31668 33983 31720 33992
rect 31668 33949 31677 33983
rect 31677 33949 31711 33983
rect 31711 33949 31720 33983
rect 31668 33940 31720 33949
rect 32496 33940 32548 33992
rect 38108 33983 38160 33992
rect 38108 33949 38117 33983
rect 38117 33949 38151 33983
rect 38151 33949 38160 33983
rect 38108 33940 38160 33949
rect 37740 33804 37792 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4620 33575 4672 33584
rect 4620 33541 4629 33575
rect 4629 33541 4663 33575
rect 4663 33541 4672 33575
rect 4620 33532 4672 33541
rect 8024 33575 8076 33584
rect 8024 33541 8033 33575
rect 8033 33541 8067 33575
rect 8067 33541 8076 33575
rect 11980 33600 12032 33652
rect 16212 33600 16264 33652
rect 20168 33600 20220 33652
rect 32496 33643 32548 33652
rect 32496 33609 32505 33643
rect 32505 33609 32539 33643
rect 32539 33609 32548 33643
rect 32496 33600 32548 33609
rect 8024 33532 8076 33541
rect 7472 33464 7524 33516
rect 2780 33439 2832 33448
rect 2780 33405 2789 33439
rect 2789 33405 2823 33439
rect 2823 33405 2832 33439
rect 2964 33439 3016 33448
rect 2780 33396 2832 33405
rect 2964 33405 2973 33439
rect 2973 33405 3007 33439
rect 3007 33405 3016 33439
rect 2964 33396 3016 33405
rect 7932 33439 7984 33448
rect 7932 33405 7941 33439
rect 7941 33405 7975 33439
rect 7975 33405 7984 33439
rect 7932 33396 7984 33405
rect 10508 33464 10560 33516
rect 12716 33464 12768 33516
rect 16672 33507 16724 33516
rect 16672 33473 16681 33507
rect 16681 33473 16715 33507
rect 16715 33473 16724 33507
rect 16672 33464 16724 33473
rect 11152 33396 11204 33448
rect 7748 33328 7800 33380
rect 7104 33303 7156 33312
rect 7104 33269 7113 33303
rect 7113 33269 7147 33303
rect 7147 33269 7156 33303
rect 7104 33260 7156 33269
rect 7564 33303 7616 33312
rect 7564 33269 7573 33303
rect 7573 33269 7607 33303
rect 7607 33269 7616 33303
rect 7564 33260 7616 33269
rect 11060 33328 11112 33380
rect 10508 33260 10560 33312
rect 16948 33439 17000 33448
rect 16948 33405 16957 33439
rect 16957 33405 16991 33439
rect 16991 33405 17000 33439
rect 16948 33396 17000 33405
rect 17224 33464 17276 33516
rect 18696 33507 18748 33516
rect 18696 33473 18705 33507
rect 18705 33473 18739 33507
rect 18739 33473 18748 33507
rect 18696 33464 18748 33473
rect 19340 33507 19392 33516
rect 19340 33473 19349 33507
rect 19349 33473 19383 33507
rect 19383 33473 19392 33507
rect 19340 33464 19392 33473
rect 18144 33396 18196 33448
rect 32312 33507 32364 33516
rect 32312 33473 32321 33507
rect 32321 33473 32355 33507
rect 32355 33473 32364 33507
rect 32312 33464 32364 33473
rect 24492 33439 24544 33448
rect 24492 33405 24501 33439
rect 24501 33405 24535 33439
rect 24535 33405 24544 33439
rect 24492 33396 24544 33405
rect 24676 33439 24728 33448
rect 24676 33405 24685 33439
rect 24685 33405 24719 33439
rect 24719 33405 24728 33439
rect 24676 33396 24728 33405
rect 25596 33439 25648 33448
rect 25596 33405 25605 33439
rect 25605 33405 25639 33439
rect 25639 33405 25648 33439
rect 25596 33396 25648 33405
rect 31576 33396 31628 33448
rect 18420 33303 18472 33312
rect 18420 33269 18429 33303
rect 18429 33269 18463 33303
rect 18463 33269 18472 33303
rect 18420 33260 18472 33269
rect 18604 33303 18656 33312
rect 18604 33269 18613 33303
rect 18613 33269 18647 33303
rect 18647 33269 18656 33303
rect 18604 33260 18656 33269
rect 19984 33260 20036 33312
rect 27160 33303 27212 33312
rect 27160 33269 27169 33303
rect 27169 33269 27203 33303
rect 27203 33269 27212 33303
rect 27160 33260 27212 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 11060 33056 11112 33108
rect 12348 33056 12400 33108
rect 17224 33099 17276 33108
rect 17224 33065 17233 33099
rect 17233 33065 17267 33099
rect 17267 33065 17276 33099
rect 17224 33056 17276 33065
rect 18696 33056 18748 33108
rect 24492 33056 24544 33108
rect 2964 32920 3016 32972
rect 11888 32920 11940 32972
rect 14556 32920 14608 32972
rect 17960 32920 18012 32972
rect 18328 32920 18380 32972
rect 23296 32920 23348 32972
rect 25596 32963 25648 32972
rect 25596 32929 25605 32963
rect 25605 32929 25639 32963
rect 25639 32929 25648 32963
rect 25596 32920 25648 32929
rect 27160 32920 27212 32972
rect 3792 32895 3844 32904
rect 3792 32861 3801 32895
rect 3801 32861 3835 32895
rect 3835 32861 3844 32895
rect 3792 32852 3844 32861
rect 7564 32852 7616 32904
rect 11152 32852 11204 32904
rect 12440 32895 12492 32904
rect 12440 32861 12449 32895
rect 12449 32861 12483 32895
rect 12483 32861 12492 32895
rect 14648 32895 14700 32904
rect 12440 32852 12492 32861
rect 14648 32861 14657 32895
rect 14657 32861 14691 32895
rect 14691 32861 14700 32895
rect 14648 32852 14700 32861
rect 15936 32852 15988 32904
rect 18144 32895 18196 32904
rect 18144 32861 18153 32895
rect 18153 32861 18187 32895
rect 18187 32861 18196 32895
rect 18144 32852 18196 32861
rect 22560 32895 22612 32904
rect 22560 32861 22569 32895
rect 22569 32861 22603 32895
rect 22603 32861 22612 32895
rect 22560 32852 22612 32861
rect 27252 32827 27304 32836
rect 7380 32716 7432 32768
rect 11520 32716 11572 32768
rect 27252 32793 27261 32827
rect 27261 32793 27295 32827
rect 27295 32793 27304 32827
rect 27252 32784 27304 32793
rect 12900 32716 12952 32768
rect 17040 32716 17092 32768
rect 19984 32716 20036 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 27252 32512 27304 32564
rect 5264 32444 5316 32496
rect 7380 32487 7432 32496
rect 7380 32453 7389 32487
rect 7389 32453 7423 32487
rect 7423 32453 7432 32487
rect 7380 32444 7432 32453
rect 15200 32444 15252 32496
rect 1400 32419 1452 32428
rect 1400 32385 1409 32419
rect 1409 32385 1443 32419
rect 1443 32385 1452 32419
rect 1400 32376 1452 32385
rect 7104 32376 7156 32428
rect 14280 32419 14332 32428
rect 14280 32385 14289 32419
rect 14289 32385 14323 32419
rect 14323 32385 14332 32419
rect 14280 32376 14332 32385
rect 18052 32376 18104 32428
rect 18788 32376 18840 32428
rect 24676 32376 24728 32428
rect 25412 32419 25464 32428
rect 25412 32385 25421 32419
rect 25421 32385 25455 32419
rect 25455 32385 25464 32419
rect 25412 32376 25464 32385
rect 2872 32351 2924 32360
rect 2872 32317 2881 32351
rect 2881 32317 2915 32351
rect 2915 32317 2924 32351
rect 2872 32308 2924 32317
rect 3056 32351 3108 32360
rect 3056 32317 3065 32351
rect 3065 32317 3099 32351
rect 3099 32317 3108 32351
rect 3056 32308 3108 32317
rect 9036 32351 9088 32360
rect 9036 32317 9045 32351
rect 9045 32317 9079 32351
rect 9079 32317 9088 32351
rect 9036 32308 9088 32317
rect 12440 32351 12492 32360
rect 12440 32317 12449 32351
rect 12449 32317 12483 32351
rect 12483 32317 12492 32351
rect 12440 32308 12492 32317
rect 19340 32351 19392 32360
rect 19340 32317 19349 32351
rect 19349 32317 19383 32351
rect 19383 32317 19392 32351
rect 19340 32308 19392 32317
rect 22100 32308 22152 32360
rect 1584 32215 1636 32224
rect 1584 32181 1593 32215
rect 1593 32181 1627 32215
rect 1627 32181 1636 32215
rect 1584 32172 1636 32181
rect 5816 32172 5868 32224
rect 18880 32215 18932 32224
rect 18880 32181 18889 32215
rect 18889 32181 18923 32215
rect 18923 32181 18932 32215
rect 18880 32172 18932 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2872 32011 2924 32020
rect 2872 31977 2881 32011
rect 2881 31977 2915 32011
rect 2915 31977 2924 32011
rect 2872 31968 2924 31977
rect 18604 31968 18656 32020
rect 24400 32011 24452 32020
rect 24400 31977 24409 32011
rect 24409 31977 24443 32011
rect 24443 31977 24452 32011
rect 24400 31968 24452 31977
rect 24492 31968 24544 32020
rect 16396 31900 16448 31952
rect 18236 31900 18288 31952
rect 37648 31943 37700 31952
rect 37648 31909 37657 31943
rect 37657 31909 37691 31943
rect 37691 31909 37700 31943
rect 37648 31900 37700 31909
rect 4160 31832 4212 31884
rect 5264 31875 5316 31884
rect 5264 31841 5273 31875
rect 5273 31841 5307 31875
rect 5307 31841 5316 31875
rect 5264 31832 5316 31841
rect 5816 31875 5868 31884
rect 5816 31841 5825 31875
rect 5825 31841 5859 31875
rect 5859 31841 5868 31875
rect 5816 31832 5868 31841
rect 6092 31832 6144 31884
rect 11520 31875 11572 31884
rect 11520 31841 11529 31875
rect 11529 31841 11563 31875
rect 11563 31841 11572 31875
rect 11520 31832 11572 31841
rect 16580 31875 16632 31884
rect 16580 31841 16589 31875
rect 16589 31841 16623 31875
rect 16623 31841 16632 31875
rect 16580 31832 16632 31841
rect 29828 31832 29880 31884
rect 33600 31875 33652 31884
rect 33600 31841 33609 31875
rect 33609 31841 33643 31875
rect 33643 31841 33652 31875
rect 33600 31832 33652 31841
rect 9864 31764 9916 31816
rect 11336 31764 11388 31816
rect 12440 31764 12492 31816
rect 13084 31764 13136 31816
rect 18420 31764 18472 31816
rect 20076 31764 20128 31816
rect 24584 31807 24636 31816
rect 24584 31773 24593 31807
rect 24593 31773 24627 31807
rect 24627 31773 24636 31807
rect 24584 31764 24636 31773
rect 5540 31696 5592 31748
rect 7932 31696 7984 31748
rect 14740 31696 14792 31748
rect 16304 31739 16356 31748
rect 16304 31705 16313 31739
rect 16313 31705 16347 31739
rect 16347 31705 16356 31739
rect 16304 31696 16356 31705
rect 24492 31696 24544 31748
rect 35256 31764 35308 31816
rect 12992 31671 13044 31680
rect 12992 31637 13001 31671
rect 13001 31637 13035 31671
rect 13035 31637 13044 31671
rect 12992 31628 13044 31637
rect 22836 31628 22888 31680
rect 29920 31739 29972 31748
rect 29920 31705 29929 31739
rect 29929 31705 29963 31739
rect 29963 31705 29972 31739
rect 29920 31696 29972 31705
rect 33140 31696 33192 31748
rect 33324 31739 33376 31748
rect 33324 31705 33333 31739
rect 33333 31705 33367 31739
rect 33367 31705 33376 31739
rect 33324 31696 33376 31705
rect 34060 31696 34112 31748
rect 34336 31696 34388 31748
rect 36176 31696 36228 31748
rect 25596 31628 25648 31680
rect 29552 31671 29604 31680
rect 29552 31637 29561 31671
rect 29561 31637 29595 31671
rect 29595 31637 29604 31671
rect 29552 31628 29604 31637
rect 30012 31671 30064 31680
rect 30012 31637 30021 31671
rect 30021 31637 30055 31671
rect 30055 31637 30064 31671
rect 30012 31628 30064 31637
rect 31392 31628 31444 31680
rect 31760 31671 31812 31680
rect 31760 31637 31769 31671
rect 31769 31637 31803 31671
rect 31803 31637 31812 31671
rect 31760 31628 31812 31637
rect 32220 31671 32272 31680
rect 32220 31637 32229 31671
rect 32229 31637 32263 31671
rect 32263 31637 32272 31671
rect 32220 31628 32272 31637
rect 32404 31628 32456 31680
rect 33416 31671 33468 31680
rect 33416 31637 33425 31671
rect 33425 31637 33459 31671
rect 33459 31637 33468 31671
rect 33416 31628 33468 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 3056 31424 3108 31476
rect 1584 31356 1636 31408
rect 3608 31356 3660 31408
rect 9036 31356 9088 31408
rect 12072 31356 12124 31408
rect 12992 31399 13044 31408
rect 1400 31331 1452 31340
rect 1400 31297 1409 31331
rect 1409 31297 1443 31331
rect 1443 31297 1452 31331
rect 1400 31288 1452 31297
rect 3884 31331 3936 31340
rect 3884 31297 3893 31331
rect 3893 31297 3927 31331
rect 3927 31297 3936 31331
rect 3884 31288 3936 31297
rect 4804 31288 4856 31340
rect 5540 31331 5592 31340
rect 5540 31297 5549 31331
rect 5549 31297 5583 31331
rect 5583 31297 5592 31331
rect 5540 31288 5592 31297
rect 12164 31331 12216 31340
rect 12164 31297 12173 31331
rect 12173 31297 12207 31331
rect 12207 31297 12216 31331
rect 12164 31288 12216 31297
rect 5816 31263 5868 31272
rect 5816 31229 5825 31263
rect 5825 31229 5859 31263
rect 5859 31229 5868 31263
rect 5816 31220 5868 31229
rect 7472 31263 7524 31272
rect 7472 31229 7481 31263
rect 7481 31229 7515 31263
rect 7515 31229 7524 31263
rect 7472 31220 7524 31229
rect 4068 31152 4120 31204
rect 8300 31152 8352 31204
rect 9036 31152 9088 31204
rect 12164 31152 12216 31204
rect 12992 31365 13001 31399
rect 13001 31365 13035 31399
rect 13035 31365 13044 31399
rect 12992 31356 13044 31365
rect 16580 31356 16632 31408
rect 17040 31399 17092 31408
rect 17040 31365 17049 31399
rect 17049 31365 17083 31399
rect 17083 31365 17092 31399
rect 17040 31356 17092 31365
rect 17960 31356 18012 31408
rect 18880 31356 18932 31408
rect 23572 31424 23624 31476
rect 26056 31467 26108 31476
rect 26056 31433 26065 31467
rect 26065 31433 26099 31467
rect 26099 31433 26108 31467
rect 26056 31424 26108 31433
rect 31668 31424 31720 31476
rect 32220 31424 32272 31476
rect 33324 31424 33376 31476
rect 23756 31356 23808 31408
rect 24492 31356 24544 31408
rect 13084 31220 13136 31272
rect 20076 31288 20128 31340
rect 21548 31288 21600 31340
rect 22192 31288 22244 31340
rect 25596 31331 25648 31340
rect 25596 31297 25605 31331
rect 25605 31297 25639 31331
rect 25639 31297 25648 31331
rect 25596 31288 25648 31297
rect 19340 31220 19392 31272
rect 21916 31263 21968 31272
rect 21916 31229 21925 31263
rect 21925 31229 21959 31263
rect 21959 31229 21968 31263
rect 21916 31220 21968 31229
rect 23296 31263 23348 31272
rect 23296 31229 23305 31263
rect 23305 31229 23339 31263
rect 23339 31229 23348 31263
rect 23296 31220 23348 31229
rect 23756 31263 23808 31272
rect 22836 31152 22888 31204
rect 22928 31152 22980 31204
rect 23756 31229 23765 31263
rect 23765 31229 23799 31263
rect 23799 31229 23808 31263
rect 23756 31220 23808 31229
rect 25044 31220 25096 31272
rect 24584 31152 24636 31204
rect 30104 31288 30156 31340
rect 31760 31356 31812 31408
rect 31300 31331 31352 31340
rect 29644 31263 29696 31272
rect 29644 31229 29653 31263
rect 29653 31229 29687 31263
rect 29687 31229 29696 31263
rect 29644 31220 29696 31229
rect 29828 31263 29880 31272
rect 29828 31229 29837 31263
rect 29837 31229 29871 31263
rect 29871 31229 29880 31263
rect 29828 31220 29880 31229
rect 31300 31297 31309 31331
rect 31309 31297 31343 31331
rect 31343 31297 31352 31331
rect 31300 31288 31352 31297
rect 31392 31331 31444 31340
rect 31392 31297 31401 31331
rect 31401 31297 31435 31331
rect 31435 31297 31444 31331
rect 34336 31331 34388 31340
rect 31392 31288 31444 31297
rect 34336 31297 34345 31331
rect 34345 31297 34379 31331
rect 34379 31297 34388 31331
rect 34336 31288 34388 31297
rect 32496 31220 32548 31272
rect 33140 31263 33192 31272
rect 29920 31152 29972 31204
rect 33140 31229 33149 31263
rect 33149 31229 33183 31263
rect 33183 31229 33192 31263
rect 33140 31220 33192 31229
rect 34796 31220 34848 31272
rect 35256 31263 35308 31272
rect 35256 31229 35265 31263
rect 35265 31229 35299 31263
rect 35299 31229 35308 31263
rect 35256 31220 35308 31229
rect 2688 31127 2740 31136
rect 2688 31093 2712 31127
rect 2712 31093 2740 31127
rect 2688 31084 2740 31093
rect 2780 31127 2832 31136
rect 2780 31093 2789 31127
rect 2789 31093 2823 31127
rect 2823 31093 2832 31127
rect 2780 31084 2832 31093
rect 3608 31084 3660 31136
rect 3976 31084 4028 31136
rect 11980 31127 12032 31136
rect 11980 31093 11989 31127
rect 11989 31093 12023 31127
rect 12023 31093 12032 31127
rect 11980 31084 12032 31093
rect 15384 31084 15436 31136
rect 21640 31084 21692 31136
rect 24400 31084 24452 31136
rect 28632 31084 28684 31136
rect 36544 31084 36596 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 7472 30923 7524 30932
rect 7472 30889 7481 30923
rect 7481 30889 7515 30923
rect 7515 30889 7524 30923
rect 7472 30880 7524 30889
rect 1400 30855 1452 30864
rect 1400 30821 1409 30855
rect 1409 30821 1443 30855
rect 1443 30821 1452 30855
rect 1400 30812 1452 30821
rect 5816 30812 5868 30864
rect 9864 30923 9916 30932
rect 9864 30889 9873 30923
rect 9873 30889 9907 30923
rect 9907 30889 9916 30923
rect 9864 30880 9916 30889
rect 15200 30923 15252 30932
rect 15200 30889 15209 30923
rect 15209 30889 15243 30923
rect 15243 30889 15252 30923
rect 15200 30880 15252 30889
rect 21640 30923 21692 30932
rect 21640 30889 21649 30923
rect 21649 30889 21683 30923
rect 21683 30889 21692 30923
rect 21640 30880 21692 30889
rect 22100 30880 22152 30932
rect 22928 30923 22980 30932
rect 22928 30889 22937 30923
rect 22937 30889 22971 30923
rect 22971 30889 22980 30923
rect 22928 30880 22980 30889
rect 23296 30880 23348 30932
rect 24400 30923 24452 30932
rect 24400 30889 24409 30923
rect 24409 30889 24443 30923
rect 24443 30889 24452 30923
rect 24400 30880 24452 30889
rect 25412 30880 25464 30932
rect 29000 30923 29052 30932
rect 29000 30889 29009 30923
rect 29009 30889 29043 30923
rect 29043 30889 29052 30923
rect 29000 30880 29052 30889
rect 29644 30880 29696 30932
rect 30012 30880 30064 30932
rect 32312 30880 32364 30932
rect 33416 30880 33468 30932
rect 36176 30880 36228 30932
rect 3976 30787 4028 30796
rect 3976 30753 3985 30787
rect 3985 30753 4019 30787
rect 4019 30753 4028 30787
rect 3976 30744 4028 30753
rect 4068 30744 4120 30796
rect 9312 30676 9364 30728
rect 11336 30787 11388 30796
rect 9496 30608 9548 30660
rect 9312 30540 9364 30592
rect 11336 30753 11345 30787
rect 11345 30753 11379 30787
rect 11379 30753 11388 30787
rect 11336 30744 11388 30753
rect 17776 30812 17828 30864
rect 14740 30787 14792 30796
rect 11152 30719 11204 30728
rect 11152 30685 11161 30719
rect 11161 30685 11195 30719
rect 11195 30685 11204 30719
rect 11152 30676 11204 30685
rect 14740 30753 14749 30787
rect 14749 30753 14783 30787
rect 14783 30753 14792 30787
rect 14740 30744 14792 30753
rect 15108 30744 15160 30796
rect 16304 30744 16356 30796
rect 22560 30812 22612 30864
rect 19984 30744 20036 30796
rect 15384 30719 15436 30728
rect 12992 30651 13044 30660
rect 12992 30617 13001 30651
rect 13001 30617 13035 30651
rect 13035 30617 13044 30651
rect 12992 30608 13044 30617
rect 14556 30651 14608 30660
rect 14556 30617 14565 30651
rect 14565 30617 14599 30651
rect 14599 30617 14608 30651
rect 14556 30608 14608 30617
rect 15384 30685 15393 30719
rect 15393 30685 15427 30719
rect 15427 30685 15436 30719
rect 15384 30676 15436 30685
rect 19524 30719 19576 30728
rect 19524 30685 19533 30719
rect 19533 30685 19567 30719
rect 19567 30685 19576 30719
rect 21916 30744 21968 30796
rect 24492 30787 24544 30796
rect 24492 30753 24501 30787
rect 24501 30753 24535 30787
rect 24535 30753 24544 30787
rect 24492 30744 24544 30753
rect 30840 30744 30892 30796
rect 33140 30744 33192 30796
rect 36728 30744 36780 30796
rect 20904 30719 20956 30728
rect 19524 30676 19576 30685
rect 20904 30685 20913 30719
rect 20913 30685 20947 30719
rect 20947 30685 20956 30719
rect 20904 30676 20956 30685
rect 22192 30676 22244 30728
rect 22744 30719 22796 30728
rect 22744 30685 22753 30719
rect 22753 30685 22787 30719
rect 22787 30685 22796 30719
rect 22744 30676 22796 30685
rect 24216 30676 24268 30728
rect 24584 30676 24636 30728
rect 28448 30719 28500 30728
rect 28448 30685 28457 30719
rect 28457 30685 28491 30719
rect 28491 30685 28500 30719
rect 28448 30676 28500 30685
rect 28632 30719 28684 30728
rect 28632 30685 28641 30719
rect 28641 30685 28675 30719
rect 28675 30685 28684 30719
rect 28632 30676 28684 30685
rect 28816 30719 28868 30728
rect 28816 30685 28825 30719
rect 28825 30685 28859 30719
rect 28859 30685 28868 30719
rect 28816 30676 28868 30685
rect 29920 30719 29972 30728
rect 29920 30685 29929 30719
rect 29929 30685 29963 30719
rect 29963 30685 29972 30719
rect 29920 30676 29972 30685
rect 30104 30676 30156 30728
rect 31392 30676 31444 30728
rect 32404 30676 32456 30728
rect 32496 30719 32548 30728
rect 32496 30685 32505 30719
rect 32505 30685 32539 30719
rect 32539 30685 32548 30719
rect 33508 30719 33560 30728
rect 32496 30676 32548 30685
rect 33508 30685 33517 30719
rect 33517 30685 33551 30719
rect 33551 30685 33560 30719
rect 33508 30676 33560 30685
rect 35440 30719 35492 30728
rect 35440 30685 35449 30719
rect 35449 30685 35483 30719
rect 35483 30685 35492 30719
rect 35440 30676 35492 30685
rect 18052 30608 18104 30660
rect 19340 30608 19392 30660
rect 20260 30608 20312 30660
rect 21548 30651 21600 30660
rect 21548 30617 21557 30651
rect 21557 30617 21591 30651
rect 21591 30617 21600 30651
rect 21548 30608 21600 30617
rect 22836 30608 22888 30660
rect 19248 30540 19300 30592
rect 20076 30540 20128 30592
rect 27988 30583 28040 30592
rect 27988 30549 27997 30583
rect 27997 30549 28031 30583
rect 28031 30549 28040 30583
rect 31852 30608 31904 30660
rect 27988 30540 28040 30549
rect 29644 30540 29696 30592
rect 31116 30583 31168 30592
rect 31116 30549 31125 30583
rect 31125 30549 31159 30583
rect 31159 30549 31168 30583
rect 33416 30583 33468 30592
rect 31116 30540 31168 30549
rect 33416 30549 33425 30583
rect 33425 30549 33459 30583
rect 33459 30549 33468 30583
rect 33416 30540 33468 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 3884 30379 3936 30388
rect 3884 30345 3893 30379
rect 3893 30345 3927 30379
rect 3927 30345 3936 30379
rect 3884 30336 3936 30345
rect 4804 30379 4856 30388
rect 4804 30345 4813 30379
rect 4813 30345 4847 30379
rect 4847 30345 4856 30379
rect 4804 30336 4856 30345
rect 19984 30336 20036 30388
rect 20536 30336 20588 30388
rect 28448 30336 28500 30388
rect 4712 30268 4764 30320
rect 12072 30268 12124 30320
rect 15660 30268 15712 30320
rect 19340 30268 19392 30320
rect 4068 30243 4120 30252
rect 4068 30209 4077 30243
rect 4077 30209 4111 30243
rect 4111 30209 4120 30243
rect 4068 30200 4120 30209
rect 11152 30200 11204 30252
rect 12256 30243 12308 30252
rect 12256 30209 12265 30243
rect 12265 30209 12299 30243
rect 12299 30209 12308 30243
rect 12256 30200 12308 30209
rect 12532 30200 12584 30252
rect 14096 30243 14148 30252
rect 4804 30064 4856 30116
rect 5080 30175 5132 30184
rect 5080 30141 5089 30175
rect 5089 30141 5123 30175
rect 5123 30141 5132 30175
rect 5080 30132 5132 30141
rect 8300 30132 8352 30184
rect 9128 30175 9180 30184
rect 9128 30141 9137 30175
rect 9137 30141 9171 30175
rect 9171 30141 9180 30175
rect 9128 30132 9180 30141
rect 9312 30175 9364 30184
rect 9312 30141 9321 30175
rect 9321 30141 9355 30175
rect 9355 30141 9364 30175
rect 9312 30132 9364 30141
rect 12164 30175 12216 30184
rect 12164 30141 12173 30175
rect 12173 30141 12207 30175
rect 12207 30141 12216 30175
rect 12164 30132 12216 30141
rect 14096 30209 14105 30243
rect 14105 30209 14139 30243
rect 14139 30209 14148 30243
rect 14096 30200 14148 30209
rect 18052 30243 18104 30252
rect 18052 30209 18061 30243
rect 18061 30209 18095 30243
rect 18095 30209 18104 30243
rect 18052 30200 18104 30209
rect 20444 30243 20496 30252
rect 20444 30209 20453 30243
rect 20453 30209 20487 30243
rect 20487 30209 20496 30243
rect 20444 30200 20496 30209
rect 21824 30200 21876 30252
rect 32404 30336 32456 30388
rect 29552 30268 29604 30320
rect 34336 30268 34388 30320
rect 12440 30107 12492 30116
rect 12440 30073 12449 30107
rect 12449 30073 12483 30107
rect 12483 30073 12492 30107
rect 18788 30107 18840 30116
rect 12440 30064 12492 30073
rect 18788 30073 18797 30107
rect 18797 30073 18831 30107
rect 18831 30073 18840 30107
rect 18788 30064 18840 30073
rect 19340 30132 19392 30184
rect 22652 30175 22704 30184
rect 22652 30141 22661 30175
rect 22661 30141 22695 30175
rect 22695 30141 22704 30175
rect 22652 30132 22704 30141
rect 23664 30175 23716 30184
rect 20352 30064 20404 30116
rect 21640 30064 21692 30116
rect 23664 30141 23673 30175
rect 23673 30141 23707 30175
rect 23707 30141 23716 30175
rect 23664 30132 23716 30141
rect 28816 30064 28868 30116
rect 30288 30200 30340 30252
rect 30472 30200 30524 30252
rect 35348 30200 35400 30252
rect 30932 30132 30984 30184
rect 30380 30064 30432 30116
rect 4620 29996 4672 30048
rect 11980 30039 12032 30048
rect 11980 30005 11989 30039
rect 11989 30005 12023 30039
rect 12023 30005 12032 30039
rect 11980 29996 12032 30005
rect 13268 30039 13320 30048
rect 13268 30005 13277 30039
rect 13277 30005 13311 30039
rect 13311 30005 13320 30039
rect 13268 29996 13320 30005
rect 13912 29996 13964 30048
rect 14556 29996 14608 30048
rect 17776 29996 17828 30048
rect 20076 29996 20128 30048
rect 28724 29996 28776 30048
rect 30748 29996 30800 30048
rect 30932 29996 30984 30048
rect 31576 29996 31628 30048
rect 34796 30132 34848 30184
rect 33416 29996 33468 30048
rect 37832 29996 37884 30048
rect 38108 30039 38160 30048
rect 38108 30005 38117 30039
rect 38117 30005 38151 30039
rect 38151 30005 38160 30039
rect 38108 29996 38160 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2780 29792 2832 29844
rect 3792 29792 3844 29844
rect 4620 29792 4672 29844
rect 9312 29792 9364 29844
rect 12072 29792 12124 29844
rect 21640 29835 21692 29844
rect 21640 29801 21649 29835
rect 21649 29801 21683 29835
rect 21683 29801 21692 29835
rect 21640 29792 21692 29801
rect 21824 29835 21876 29844
rect 21824 29801 21833 29835
rect 21833 29801 21867 29835
rect 21867 29801 21876 29835
rect 21824 29792 21876 29801
rect 22744 29835 22796 29844
rect 12164 29724 12216 29776
rect 18144 29724 18196 29776
rect 22744 29801 22753 29835
rect 22753 29801 22787 29835
rect 22787 29801 22796 29835
rect 22744 29792 22796 29801
rect 34796 29792 34848 29844
rect 35348 29792 35400 29844
rect 22652 29724 22704 29776
rect 31392 29724 31444 29776
rect 37188 29724 37240 29776
rect 4804 29656 4856 29708
rect 11980 29656 12032 29708
rect 15660 29699 15712 29708
rect 15660 29665 15669 29699
rect 15669 29665 15703 29699
rect 15703 29665 15712 29699
rect 15660 29656 15712 29665
rect 17776 29699 17828 29708
rect 17776 29665 17785 29699
rect 17785 29665 17819 29699
rect 17819 29665 17828 29699
rect 17776 29656 17828 29665
rect 20352 29656 20404 29708
rect 21548 29699 21600 29708
rect 1400 29631 1452 29640
rect 1400 29597 1409 29631
rect 1409 29597 1443 29631
rect 1443 29597 1452 29631
rect 1400 29588 1452 29597
rect 4068 29631 4120 29640
rect 4068 29597 4077 29631
rect 4077 29597 4111 29631
rect 4111 29597 4120 29631
rect 4068 29588 4120 29597
rect 4712 29588 4764 29640
rect 8116 29520 8168 29572
rect 14096 29588 14148 29640
rect 15844 29588 15896 29640
rect 20444 29588 20496 29640
rect 21548 29665 21557 29699
rect 21557 29665 21591 29699
rect 21591 29665 21600 29699
rect 21548 29656 21600 29665
rect 28724 29656 28776 29708
rect 29920 29656 29972 29708
rect 31852 29699 31904 29708
rect 31852 29665 31861 29699
rect 31861 29665 31895 29699
rect 31895 29665 31904 29699
rect 31852 29656 31904 29665
rect 36728 29699 36780 29708
rect 36728 29665 36737 29699
rect 36737 29665 36771 29699
rect 36771 29665 36780 29699
rect 36728 29656 36780 29665
rect 37832 29699 37884 29708
rect 37832 29665 37841 29699
rect 37841 29665 37875 29699
rect 37875 29665 37884 29699
rect 37832 29656 37884 29665
rect 14004 29452 14056 29504
rect 15292 29452 15344 29504
rect 20904 29588 20956 29640
rect 34520 29588 34572 29640
rect 35900 29588 35952 29640
rect 36544 29631 36596 29640
rect 36544 29597 36553 29631
rect 36553 29597 36587 29631
rect 36587 29597 36596 29631
rect 36544 29588 36596 29597
rect 37740 29631 37792 29640
rect 37740 29597 37749 29631
rect 37749 29597 37783 29631
rect 37783 29597 37792 29631
rect 37740 29588 37792 29597
rect 21364 29563 21416 29572
rect 21364 29529 21373 29563
rect 21373 29529 21407 29563
rect 21407 29529 21416 29563
rect 21364 29520 21416 29529
rect 28816 29563 28868 29572
rect 28816 29529 28825 29563
rect 28825 29529 28859 29563
rect 28859 29529 28868 29563
rect 28816 29520 28868 29529
rect 30748 29563 30800 29572
rect 30748 29529 30757 29563
rect 30757 29529 30791 29563
rect 30791 29529 30800 29563
rect 30748 29520 30800 29529
rect 29000 29452 29052 29504
rect 29736 29495 29788 29504
rect 29736 29461 29745 29495
rect 29745 29461 29779 29495
rect 29779 29461 29788 29495
rect 29736 29452 29788 29461
rect 36176 29495 36228 29504
rect 36176 29461 36185 29495
rect 36185 29461 36219 29495
rect 36219 29461 36228 29495
rect 36176 29452 36228 29461
rect 37372 29495 37424 29504
rect 37372 29461 37381 29495
rect 37381 29461 37415 29495
rect 37415 29461 37424 29495
rect 37372 29452 37424 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 9128 29248 9180 29300
rect 18144 29291 18196 29300
rect 18144 29257 18153 29291
rect 18153 29257 18187 29291
rect 18187 29257 18196 29291
rect 18144 29248 18196 29257
rect 20260 29291 20312 29300
rect 20260 29257 20269 29291
rect 20269 29257 20303 29291
rect 20303 29257 20312 29291
rect 20260 29248 20312 29257
rect 30472 29291 30524 29300
rect 13268 29180 13320 29232
rect 3700 29087 3752 29096
rect 3700 29053 3709 29087
rect 3709 29053 3743 29087
rect 3743 29053 3752 29087
rect 3700 29044 3752 29053
rect 3884 29044 3936 29096
rect 9772 29044 9824 29096
rect 12992 29087 13044 29096
rect 12992 29053 13001 29087
rect 13001 29053 13035 29087
rect 13035 29053 13044 29087
rect 12992 29044 13044 29053
rect 13820 29087 13872 29096
rect 13820 29053 13829 29087
rect 13829 29053 13863 29087
rect 13863 29053 13872 29087
rect 13820 29044 13872 29053
rect 15108 29155 15160 29164
rect 15108 29121 15117 29155
rect 15117 29121 15151 29155
rect 15151 29121 15160 29155
rect 15108 29112 15160 29121
rect 15292 29155 15344 29164
rect 15292 29121 15301 29155
rect 15301 29121 15335 29155
rect 15335 29121 15344 29155
rect 24492 29180 24544 29232
rect 15292 29112 15344 29121
rect 17224 29155 17276 29164
rect 17224 29121 17233 29155
rect 17233 29121 17267 29155
rect 17267 29121 17276 29155
rect 17224 29112 17276 29121
rect 16672 29044 16724 29096
rect 18880 29044 18932 29096
rect 19340 29112 19392 29164
rect 20720 29112 20772 29164
rect 19432 29044 19484 29096
rect 24124 29155 24176 29164
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 15936 29019 15988 29028
rect 15936 28985 15945 29019
rect 15945 28985 15979 29019
rect 15979 28985 15988 29019
rect 15936 28976 15988 28985
rect 23296 28976 23348 29028
rect 24308 29019 24360 29028
rect 24308 28985 24317 29019
rect 24317 28985 24351 29019
rect 24351 28985 24360 29019
rect 24308 28976 24360 28985
rect 28908 29044 28960 29096
rect 29736 29180 29788 29232
rect 30472 29257 30481 29291
rect 30481 29257 30515 29291
rect 30515 29257 30524 29291
rect 30472 29248 30524 29257
rect 31116 29180 31168 29232
rect 31392 29180 31444 29232
rect 30104 29155 30156 29164
rect 30104 29121 30113 29155
rect 30113 29121 30147 29155
rect 30147 29121 30156 29155
rect 30104 29112 30156 29121
rect 30288 29155 30340 29164
rect 30288 29121 30297 29155
rect 30297 29121 30331 29155
rect 30331 29121 30340 29155
rect 30288 29112 30340 29121
rect 31300 28976 31352 29028
rect 8668 28951 8720 28960
rect 8668 28917 8677 28951
rect 8677 28917 8711 28951
rect 8711 28917 8720 28951
rect 8668 28908 8720 28917
rect 9128 28908 9180 28960
rect 14832 28951 14884 28960
rect 14832 28917 14841 28951
rect 14841 28917 14875 28951
rect 14875 28917 14884 28951
rect 14832 28908 14884 28917
rect 15844 28908 15896 28960
rect 20720 28951 20772 28960
rect 20720 28917 20729 28951
rect 20729 28917 20763 28951
rect 20763 28917 20772 28951
rect 20720 28908 20772 28917
rect 24216 28908 24268 28960
rect 32036 28976 32088 29028
rect 32496 28908 32548 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 3700 28704 3752 28756
rect 4620 28704 4672 28756
rect 15844 28747 15896 28756
rect 15844 28713 15853 28747
rect 15853 28713 15887 28747
rect 15887 28713 15896 28747
rect 15844 28704 15896 28713
rect 24400 28747 24452 28756
rect 24400 28713 24409 28747
rect 24409 28713 24443 28747
rect 24443 28713 24452 28747
rect 24400 28704 24452 28713
rect 30104 28704 30156 28756
rect 31392 28704 31444 28756
rect 33600 28747 33652 28756
rect 33600 28713 33609 28747
rect 33609 28713 33643 28747
rect 33643 28713 33652 28747
rect 33600 28704 33652 28713
rect 1400 28543 1452 28552
rect 1400 28509 1409 28543
rect 1409 28509 1443 28543
rect 1443 28509 1452 28543
rect 1400 28500 1452 28509
rect 2780 28500 2832 28552
rect 4804 28568 4856 28620
rect 8668 28568 8720 28620
rect 9772 28611 9824 28620
rect 9772 28577 9781 28611
rect 9781 28577 9815 28611
rect 9815 28577 9824 28611
rect 9772 28568 9824 28577
rect 12256 28568 12308 28620
rect 13820 28568 13872 28620
rect 14832 28568 14884 28620
rect 16580 28568 16632 28620
rect 24032 28568 24084 28620
rect 29828 28568 29880 28620
rect 4160 28543 4212 28552
rect 4160 28509 4169 28543
rect 4169 28509 4203 28543
rect 4203 28509 4212 28543
rect 4160 28500 4212 28509
rect 4712 28500 4764 28552
rect 5264 28500 5316 28552
rect 8116 28500 8168 28552
rect 13084 28500 13136 28552
rect 15936 28500 15988 28552
rect 2596 28364 2648 28416
rect 4988 28407 5040 28416
rect 4988 28373 4997 28407
rect 4997 28373 5031 28407
rect 5031 28373 5040 28407
rect 9220 28432 9272 28484
rect 17040 28432 17092 28484
rect 24216 28500 24268 28552
rect 25504 28543 25556 28552
rect 25504 28509 25513 28543
rect 25513 28509 25547 28543
rect 25547 28509 25556 28543
rect 25504 28500 25556 28509
rect 29644 28500 29696 28552
rect 29920 28543 29972 28552
rect 29920 28509 29929 28543
rect 29929 28509 29963 28543
rect 29963 28509 29972 28543
rect 29920 28500 29972 28509
rect 35900 28500 35952 28552
rect 36360 28500 36412 28552
rect 23940 28432 23992 28484
rect 33784 28432 33836 28484
rect 4988 28364 5040 28373
rect 16856 28364 16908 28416
rect 22744 28364 22796 28416
rect 24860 28407 24912 28416
rect 24860 28373 24869 28407
rect 24869 28373 24903 28407
rect 24903 28373 24912 28407
rect 24860 28364 24912 28373
rect 29644 28364 29696 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4712 28160 4764 28212
rect 1400 28135 1452 28144
rect 1400 28101 1409 28135
rect 1409 28101 1443 28135
rect 1443 28101 1452 28135
rect 1400 28092 1452 28101
rect 2780 28067 2832 28076
rect 2780 28033 2789 28067
rect 2789 28033 2823 28067
rect 2823 28033 2832 28067
rect 2780 28024 2832 28033
rect 5264 28067 5316 28076
rect 5264 28033 5273 28067
rect 5273 28033 5307 28067
rect 5307 28033 5316 28067
rect 5264 28024 5316 28033
rect 9128 28067 9180 28076
rect 9128 28033 9137 28067
rect 9137 28033 9171 28067
rect 9171 28033 9180 28067
rect 9128 28024 9180 28033
rect 14924 28067 14976 28076
rect 14924 28033 14933 28067
rect 14933 28033 14967 28067
rect 14967 28033 14976 28067
rect 14924 28024 14976 28033
rect 2964 27999 3016 28008
rect 2964 27965 2973 27999
rect 2973 27965 3007 27999
rect 3007 27965 3016 27999
rect 2964 27956 3016 27965
rect 3240 27999 3292 28008
rect 3240 27965 3249 27999
rect 3249 27965 3283 27999
rect 3283 27965 3292 27999
rect 9312 27999 9364 28008
rect 3240 27956 3292 27965
rect 9312 27965 9321 27999
rect 9321 27965 9355 27999
rect 9355 27965 9364 27999
rect 9312 27956 9364 27965
rect 12992 27956 13044 28008
rect 16580 28160 16632 28212
rect 29644 28203 29696 28212
rect 29644 28169 29653 28203
rect 29653 28169 29687 28203
rect 29687 28169 29696 28203
rect 29644 28160 29696 28169
rect 30012 28203 30064 28212
rect 30012 28169 30021 28203
rect 30021 28169 30055 28203
rect 30055 28169 30064 28203
rect 30012 28160 30064 28169
rect 35440 28160 35492 28212
rect 17040 28092 17092 28144
rect 23664 28135 23716 28144
rect 23664 28101 23673 28135
rect 23673 28101 23707 28135
rect 23707 28101 23716 28135
rect 23664 28092 23716 28101
rect 32496 28135 32548 28144
rect 32496 28101 32505 28135
rect 32505 28101 32539 28135
rect 32539 28101 32548 28135
rect 32496 28092 32548 28101
rect 15936 28024 15988 28076
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 25504 28067 25556 28076
rect 25504 28033 25513 28067
rect 25513 28033 25547 28067
rect 25547 28033 25556 28067
rect 25504 28024 25556 28033
rect 28816 28024 28868 28076
rect 32220 28024 32272 28076
rect 33324 28024 33376 28076
rect 18880 27956 18932 28008
rect 21640 27956 21692 28008
rect 25320 27999 25372 28008
rect 25320 27965 25329 27999
rect 25329 27965 25363 27999
rect 25363 27965 25372 27999
rect 25320 27956 25372 27965
rect 26240 27956 26292 28008
rect 29736 27956 29788 28008
rect 30840 27956 30892 28008
rect 33600 27956 33652 28008
rect 13084 27820 13136 27872
rect 14280 27863 14332 27872
rect 14280 27829 14289 27863
rect 14289 27829 14323 27863
rect 14323 27829 14332 27863
rect 14280 27820 14332 27829
rect 14464 27820 14516 27872
rect 15384 27863 15436 27872
rect 15384 27829 15393 27863
rect 15393 27829 15427 27863
rect 15427 27829 15436 27863
rect 15384 27820 15436 27829
rect 15844 27888 15896 27940
rect 16488 27888 16540 27940
rect 15660 27820 15712 27872
rect 20720 27863 20772 27872
rect 20720 27829 20729 27863
rect 20729 27829 20763 27863
rect 20763 27829 20772 27863
rect 20720 27820 20772 27829
rect 26148 27863 26200 27872
rect 26148 27829 26157 27863
rect 26157 27829 26191 27863
rect 26191 27829 26200 27863
rect 26148 27820 26200 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2964 27616 3016 27668
rect 4620 27616 4672 27668
rect 5080 27616 5132 27668
rect 16488 27616 16540 27668
rect 29736 27616 29788 27668
rect 9312 27548 9364 27600
rect 25320 27548 25372 27600
rect 26148 27548 26200 27600
rect 4620 27480 4672 27532
rect 4804 27480 4856 27532
rect 14280 27480 14332 27532
rect 15660 27480 15712 27532
rect 15752 27523 15804 27532
rect 15752 27489 15761 27523
rect 15761 27489 15795 27523
rect 15795 27489 15804 27523
rect 15752 27480 15804 27489
rect 16580 27480 16632 27532
rect 17684 27480 17736 27532
rect 24032 27480 24084 27532
rect 24308 27480 24360 27532
rect 34520 27548 34572 27600
rect 28908 27480 28960 27532
rect 33600 27480 33652 27532
rect 4712 27412 4764 27464
rect 9036 27455 9088 27464
rect 9036 27421 9045 27455
rect 9045 27421 9079 27455
rect 9079 27421 9088 27455
rect 9036 27412 9088 27421
rect 9220 27412 9272 27464
rect 9772 27412 9824 27464
rect 11428 27412 11480 27464
rect 15936 27412 15988 27464
rect 4160 27344 4212 27396
rect 17040 27344 17092 27396
rect 18512 27455 18564 27464
rect 18512 27421 18521 27455
rect 18521 27421 18555 27455
rect 18555 27421 18564 27455
rect 18512 27412 18564 27421
rect 19340 27412 19392 27464
rect 20628 27412 20680 27464
rect 21364 27412 21416 27464
rect 24860 27412 24912 27464
rect 26700 27455 26752 27464
rect 26700 27421 26709 27455
rect 26709 27421 26743 27455
rect 26743 27421 26752 27455
rect 26700 27412 26752 27421
rect 33692 27455 33744 27464
rect 33692 27421 33701 27455
rect 33701 27421 33735 27455
rect 33735 27421 33744 27455
rect 33692 27412 33744 27421
rect 35992 27480 36044 27532
rect 37004 27523 37056 27532
rect 37004 27489 37013 27523
rect 37013 27489 37047 27523
rect 37047 27489 37056 27523
rect 37004 27480 37056 27489
rect 19432 27344 19484 27396
rect 20260 27344 20312 27396
rect 24676 27344 24728 27396
rect 25044 27344 25096 27396
rect 36176 27412 36228 27464
rect 37648 27412 37700 27464
rect 36084 27344 36136 27396
rect 18696 27276 18748 27328
rect 31944 27276 31996 27328
rect 33232 27276 33284 27328
rect 35624 27276 35676 27328
rect 36820 27319 36872 27328
rect 36820 27285 36829 27319
rect 36829 27285 36863 27319
rect 36863 27285 36872 27319
rect 36820 27276 36872 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 9772 27115 9824 27124
rect 9772 27081 9781 27115
rect 9781 27081 9815 27115
rect 9815 27081 9824 27115
rect 9772 27072 9824 27081
rect 24124 27072 24176 27124
rect 31392 27072 31444 27124
rect 31668 27072 31720 27124
rect 9496 27004 9548 27056
rect 14464 27047 14516 27056
rect 14464 27013 14473 27047
rect 14473 27013 14507 27047
rect 14507 27013 14516 27047
rect 14464 27004 14516 27013
rect 18696 27047 18748 27056
rect 18696 27013 18705 27047
rect 18705 27013 18739 27047
rect 18739 27013 18748 27047
rect 18696 27004 18748 27013
rect 23940 27047 23992 27056
rect 23940 27013 23949 27047
rect 23949 27013 23983 27047
rect 23983 27013 23992 27047
rect 23940 27004 23992 27013
rect 31944 27004 31996 27056
rect 1400 26979 1452 26988
rect 1400 26945 1409 26979
rect 1409 26945 1443 26979
rect 1443 26945 1452 26979
rect 1400 26936 1452 26945
rect 9588 26979 9640 26988
rect 9588 26945 9597 26979
rect 9597 26945 9631 26979
rect 9631 26945 9640 26979
rect 9588 26936 9640 26945
rect 10416 26979 10468 26988
rect 10416 26945 10425 26979
rect 10425 26945 10459 26979
rect 10459 26945 10468 26979
rect 10416 26936 10468 26945
rect 18052 26936 18104 26988
rect 18512 26979 18564 26988
rect 18512 26945 18521 26979
rect 18521 26945 18555 26979
rect 18555 26945 18564 26979
rect 18512 26936 18564 26945
rect 24216 26979 24268 26988
rect 24216 26945 24225 26979
rect 24225 26945 24259 26979
rect 24259 26945 24268 26979
rect 24216 26936 24268 26945
rect 30012 26936 30064 26988
rect 32220 26979 32272 26988
rect 32220 26945 32229 26979
rect 32229 26945 32263 26979
rect 32263 26945 32272 26979
rect 32220 26936 32272 26945
rect 32404 26979 32456 26988
rect 32404 26945 32413 26979
rect 32413 26945 32447 26979
rect 32447 26945 32456 26979
rect 32404 26936 32456 26945
rect 33692 27072 33744 27124
rect 34060 27115 34112 27124
rect 34060 27081 34069 27115
rect 34069 27081 34103 27115
rect 34103 27081 34112 27115
rect 34060 27072 34112 27081
rect 36820 27072 36872 27124
rect 37188 27004 37240 27056
rect 9220 26868 9272 26920
rect 9404 26911 9456 26920
rect 9404 26877 9413 26911
rect 9413 26877 9447 26911
rect 9447 26877 9456 26911
rect 9404 26868 9456 26877
rect 14280 26911 14332 26920
rect 14280 26877 14289 26911
rect 14289 26877 14323 26911
rect 14323 26877 14332 26911
rect 14280 26868 14332 26877
rect 3976 26800 4028 26852
rect 5540 26800 5592 26852
rect 11888 26800 11940 26852
rect 15752 26868 15804 26920
rect 17684 26868 17736 26920
rect 19432 26911 19484 26920
rect 19432 26877 19441 26911
rect 19441 26877 19475 26911
rect 19475 26877 19484 26911
rect 19432 26868 19484 26877
rect 24032 26911 24084 26920
rect 24032 26877 24041 26911
rect 24041 26877 24075 26911
rect 24075 26877 24084 26911
rect 24032 26868 24084 26877
rect 24492 26868 24544 26920
rect 27988 26911 28040 26920
rect 27988 26877 27997 26911
rect 27997 26877 28031 26911
rect 28031 26877 28040 26911
rect 27988 26868 28040 26877
rect 28080 26868 28132 26920
rect 31392 26800 31444 26852
rect 34060 26800 34112 26852
rect 1584 26775 1636 26784
rect 1584 26741 1593 26775
rect 1593 26741 1627 26775
rect 1627 26741 1636 26775
rect 1584 26732 1636 26741
rect 4712 26775 4764 26784
rect 4712 26741 4721 26775
rect 4721 26741 4755 26775
rect 4755 26741 4764 26775
rect 4712 26732 4764 26741
rect 5172 26775 5224 26784
rect 5172 26741 5181 26775
rect 5181 26741 5215 26775
rect 5215 26741 5224 26775
rect 5172 26732 5224 26741
rect 9404 26775 9456 26784
rect 9404 26741 9413 26775
rect 9413 26741 9447 26775
rect 9447 26741 9456 26775
rect 9404 26732 9456 26741
rect 11612 26732 11664 26784
rect 24400 26732 24452 26784
rect 33508 26732 33560 26784
rect 36452 26936 36504 26988
rect 37096 26936 37148 26988
rect 35992 26868 36044 26920
rect 36176 26868 36228 26920
rect 37188 26800 37240 26852
rect 35900 26732 35952 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 4620 26528 4672 26580
rect 5540 26460 5592 26512
rect 11888 26528 11940 26580
rect 14280 26528 14332 26580
rect 14924 26528 14976 26580
rect 16488 26571 16540 26580
rect 16488 26537 16497 26571
rect 16497 26537 16531 26571
rect 16531 26537 16540 26571
rect 16488 26528 16540 26537
rect 18052 26571 18104 26580
rect 18052 26537 18061 26571
rect 18061 26537 18095 26571
rect 18095 26537 18104 26571
rect 18052 26528 18104 26537
rect 18420 26528 18472 26580
rect 32404 26528 32456 26580
rect 36452 26571 36504 26580
rect 36452 26537 36461 26571
rect 36461 26537 36495 26571
rect 36495 26537 36504 26571
rect 36452 26528 36504 26537
rect 5172 26435 5224 26444
rect 5172 26401 5181 26435
rect 5181 26401 5215 26435
rect 5215 26401 5224 26435
rect 5172 26392 5224 26401
rect 11428 26435 11480 26444
rect 5356 26299 5408 26308
rect 5356 26265 5365 26299
rect 5365 26265 5399 26299
rect 5399 26265 5408 26299
rect 5356 26256 5408 26265
rect 5632 26256 5684 26308
rect 11428 26401 11437 26435
rect 11437 26401 11471 26435
rect 11471 26401 11480 26435
rect 11428 26392 11480 26401
rect 11612 26435 11664 26444
rect 11612 26401 11621 26435
rect 11621 26401 11655 26435
rect 11655 26401 11664 26435
rect 11612 26392 11664 26401
rect 29552 26460 29604 26512
rect 30288 26460 30340 26512
rect 31852 26460 31904 26512
rect 15384 26392 15436 26444
rect 14096 26324 14148 26376
rect 15936 26324 15988 26376
rect 16396 26367 16448 26376
rect 16396 26333 16405 26367
rect 16405 26333 16439 26367
rect 16439 26333 16448 26367
rect 16396 26324 16448 26333
rect 9312 26299 9364 26308
rect 5448 26188 5500 26240
rect 9312 26265 9321 26299
rect 9321 26265 9355 26299
rect 9355 26265 9364 26299
rect 9312 26256 9364 26265
rect 19432 26392 19484 26444
rect 30932 26392 30984 26444
rect 31392 26435 31444 26444
rect 31392 26401 31401 26435
rect 31401 26401 31435 26435
rect 31435 26401 31444 26435
rect 31392 26392 31444 26401
rect 32220 26392 32272 26444
rect 33140 26460 33192 26512
rect 38016 26503 38068 26512
rect 38016 26469 38025 26503
rect 38025 26469 38059 26503
rect 38059 26469 38068 26503
rect 38016 26460 38068 26469
rect 33324 26392 33376 26444
rect 33508 26435 33560 26444
rect 33508 26401 33517 26435
rect 33517 26401 33551 26435
rect 33551 26401 33560 26435
rect 33508 26392 33560 26401
rect 33784 26392 33836 26444
rect 35992 26392 36044 26444
rect 36636 26392 36688 26444
rect 37096 26435 37148 26444
rect 37096 26401 37105 26435
rect 37105 26401 37139 26435
rect 37139 26401 37148 26435
rect 37096 26392 37148 26401
rect 16672 26324 16724 26376
rect 27712 26367 27764 26376
rect 27712 26333 27721 26367
rect 27721 26333 27755 26367
rect 27755 26333 27764 26367
rect 27712 26324 27764 26333
rect 29552 26367 29604 26376
rect 29552 26333 29561 26367
rect 29561 26333 29595 26367
rect 29595 26333 29604 26367
rect 29552 26324 29604 26333
rect 32036 26367 32088 26376
rect 32036 26333 32045 26367
rect 32045 26333 32079 26367
rect 32079 26333 32088 26367
rect 32036 26324 32088 26333
rect 19432 26299 19484 26308
rect 19432 26265 19441 26299
rect 19441 26265 19475 26299
rect 19475 26265 19484 26299
rect 19432 26256 19484 26265
rect 25688 26256 25740 26308
rect 26884 26256 26936 26308
rect 30012 26256 30064 26308
rect 32220 26299 32272 26308
rect 32220 26265 32229 26299
rect 32229 26265 32263 26299
rect 32263 26265 32272 26299
rect 32220 26256 32272 26265
rect 35624 26324 35676 26376
rect 37372 26324 37424 26376
rect 37648 26324 37700 26376
rect 32680 26256 32732 26308
rect 33416 26299 33468 26308
rect 33416 26265 33425 26299
rect 33425 26265 33459 26299
rect 33459 26265 33468 26299
rect 33416 26256 33468 26265
rect 35900 26188 35952 26240
rect 36084 26188 36136 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 2964 25984 3016 26036
rect 5356 26027 5408 26036
rect 5356 25993 5365 26027
rect 5365 25993 5399 26027
rect 5399 25993 5408 26027
rect 5356 25984 5408 25993
rect 9036 25984 9088 26036
rect 9404 25984 9456 26036
rect 9772 25984 9824 26036
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 1584 25848 1636 25900
rect 2872 25848 2924 25900
rect 4160 25848 4212 25900
rect 4804 25848 4856 25900
rect 5172 25891 5224 25900
rect 5172 25857 5181 25891
rect 5181 25857 5215 25891
rect 5215 25857 5224 25891
rect 5172 25848 5224 25857
rect 9588 25916 9640 25968
rect 10048 25916 10100 25968
rect 9404 25891 9456 25900
rect 9404 25857 9413 25891
rect 9413 25857 9447 25891
rect 9447 25857 9456 25891
rect 9404 25848 9456 25857
rect 9956 25848 10008 25900
rect 12532 25916 12584 25968
rect 14004 25984 14056 26036
rect 36176 25984 36228 26036
rect 36360 26027 36412 26036
rect 36360 25993 36369 26027
rect 36369 25993 36403 26027
rect 36403 25993 36412 26027
rect 36360 25984 36412 25993
rect 14096 25959 14148 25968
rect 14096 25925 14105 25959
rect 14105 25925 14139 25959
rect 14139 25925 14148 25959
rect 14096 25916 14148 25925
rect 30932 25959 30984 25968
rect 30932 25925 30941 25959
rect 30941 25925 30975 25959
rect 30975 25925 30984 25959
rect 30932 25916 30984 25925
rect 32036 25916 32088 25968
rect 33416 25916 33468 25968
rect 13268 25848 13320 25900
rect 24492 25848 24544 25900
rect 28080 25848 28132 25900
rect 32128 25848 32180 25900
rect 32680 25891 32732 25900
rect 32680 25857 32689 25891
rect 32689 25857 32723 25891
rect 32723 25857 32732 25891
rect 32680 25848 32732 25857
rect 33232 25848 33284 25900
rect 4620 25780 4672 25832
rect 4988 25780 5040 25832
rect 5356 25780 5408 25832
rect 9220 25823 9272 25832
rect 9220 25789 9229 25823
rect 9229 25789 9263 25823
rect 9263 25789 9272 25823
rect 9220 25780 9272 25789
rect 10232 25780 10284 25832
rect 15292 25823 15344 25832
rect 15292 25789 15301 25823
rect 15301 25789 15335 25823
rect 15335 25789 15344 25823
rect 15292 25780 15344 25789
rect 25872 25780 25924 25832
rect 29276 25823 29328 25832
rect 29276 25789 29285 25823
rect 29285 25789 29319 25823
rect 29319 25789 29328 25823
rect 29276 25780 29328 25789
rect 33416 25780 33468 25832
rect 36636 25823 36688 25832
rect 36636 25789 36645 25823
rect 36645 25789 36679 25823
rect 36679 25789 36688 25823
rect 36636 25780 36688 25789
rect 2596 25687 2648 25696
rect 2596 25653 2605 25687
rect 2605 25653 2639 25687
rect 2639 25653 2648 25687
rect 2596 25644 2648 25653
rect 5080 25712 5132 25764
rect 9312 25712 9364 25764
rect 22468 25755 22520 25764
rect 4988 25644 5040 25696
rect 9772 25644 9824 25696
rect 10324 25644 10376 25696
rect 22468 25721 22477 25755
rect 22477 25721 22511 25755
rect 22511 25721 22520 25755
rect 22468 25712 22520 25721
rect 31944 25712 31996 25764
rect 32128 25712 32180 25764
rect 10968 25644 11020 25696
rect 11704 25644 11756 25696
rect 23020 25644 23072 25696
rect 25412 25644 25464 25696
rect 26056 25644 26108 25696
rect 32956 25687 33008 25696
rect 32956 25653 32965 25687
rect 32965 25653 32999 25687
rect 32999 25653 33008 25687
rect 32956 25644 33008 25653
rect 35900 25644 35952 25696
rect 36268 25644 36320 25696
rect 37648 25687 37700 25696
rect 37648 25653 37657 25687
rect 37657 25653 37691 25687
rect 37691 25653 37700 25687
rect 37648 25644 37700 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1400 25415 1452 25424
rect 1400 25381 1409 25415
rect 1409 25381 1443 25415
rect 1443 25381 1452 25415
rect 1400 25372 1452 25381
rect 5172 25440 5224 25492
rect 10416 25440 10468 25492
rect 11704 25483 11756 25492
rect 11704 25449 11713 25483
rect 11713 25449 11747 25483
rect 11747 25449 11756 25483
rect 11704 25440 11756 25449
rect 19432 25483 19484 25492
rect 19432 25449 19441 25483
rect 19441 25449 19475 25483
rect 19475 25449 19484 25483
rect 19432 25440 19484 25449
rect 21824 25483 21876 25492
rect 21824 25449 21833 25483
rect 21833 25449 21867 25483
rect 21867 25449 21876 25483
rect 21824 25440 21876 25449
rect 25872 25483 25924 25492
rect 5080 25372 5132 25424
rect 10232 25372 10284 25424
rect 25872 25449 25881 25483
rect 25881 25449 25915 25483
rect 25915 25449 25924 25483
rect 25872 25440 25924 25449
rect 4620 25304 4672 25356
rect 4712 25304 4764 25356
rect 4988 25347 5040 25356
rect 4988 25313 4997 25347
rect 4997 25313 5031 25347
rect 5031 25313 5040 25347
rect 4988 25304 5040 25313
rect 5540 25347 5592 25356
rect 5540 25313 5549 25347
rect 5549 25313 5583 25347
rect 5583 25313 5592 25347
rect 5540 25304 5592 25313
rect 9772 25347 9824 25356
rect 9772 25313 9781 25347
rect 9781 25313 9815 25347
rect 9815 25313 9824 25347
rect 9772 25304 9824 25313
rect 10048 25304 10100 25356
rect 10968 25304 11020 25356
rect 26148 25372 26200 25424
rect 26700 25440 26752 25492
rect 32220 25440 32272 25492
rect 2596 25279 2648 25288
rect 2596 25245 2605 25279
rect 2605 25245 2639 25279
rect 2639 25245 2648 25279
rect 2596 25236 2648 25245
rect 3240 25279 3292 25288
rect 3240 25245 3249 25279
rect 3249 25245 3283 25279
rect 3283 25245 3292 25279
rect 3240 25236 3292 25245
rect 4160 25279 4212 25288
rect 4160 25245 4169 25279
rect 4169 25245 4203 25279
rect 4203 25245 4212 25279
rect 21640 25347 21692 25356
rect 21640 25313 21649 25347
rect 21649 25313 21683 25347
rect 21683 25313 21692 25347
rect 21640 25304 21692 25313
rect 24952 25304 25004 25356
rect 26056 25304 26108 25356
rect 30012 25304 30064 25356
rect 30840 25304 30892 25356
rect 4160 25236 4212 25245
rect 4712 25168 4764 25220
rect 19248 25279 19300 25288
rect 19248 25245 19257 25279
rect 19257 25245 19291 25279
rect 19291 25245 19300 25279
rect 19248 25236 19300 25245
rect 21364 25236 21416 25288
rect 9128 25211 9180 25220
rect 9128 25177 9137 25211
rect 9137 25177 9171 25211
rect 9171 25177 9180 25211
rect 9128 25168 9180 25177
rect 9956 25168 10008 25220
rect 21916 25236 21968 25288
rect 25688 25279 25740 25288
rect 25688 25245 25697 25279
rect 25697 25245 25731 25279
rect 25731 25245 25740 25279
rect 25688 25236 25740 25245
rect 26976 25236 27028 25288
rect 30380 25279 30432 25288
rect 30380 25245 30389 25279
rect 30389 25245 30423 25279
rect 30423 25245 30432 25279
rect 30380 25236 30432 25245
rect 30932 25236 30984 25288
rect 21732 25168 21784 25220
rect 22836 25168 22888 25220
rect 25412 25211 25464 25220
rect 25412 25177 25421 25211
rect 25421 25177 25455 25211
rect 25455 25177 25464 25211
rect 25412 25168 25464 25177
rect 2780 25100 2832 25152
rect 4804 25100 4856 25152
rect 22008 25143 22060 25152
rect 22008 25109 22017 25143
rect 22017 25109 22051 25143
rect 22051 25109 22060 25143
rect 22008 25100 22060 25109
rect 24952 25143 25004 25152
rect 24952 25109 24961 25143
rect 24961 25109 24995 25143
rect 24995 25109 25004 25143
rect 24952 25100 25004 25109
rect 25780 25100 25832 25152
rect 26056 25100 26108 25152
rect 31116 25168 31168 25220
rect 29552 25100 29604 25152
rect 32128 25236 32180 25288
rect 32312 25236 32364 25288
rect 32680 25236 32732 25288
rect 33140 25304 33192 25356
rect 33232 25279 33284 25288
rect 33232 25245 33241 25279
rect 33241 25245 33275 25279
rect 33275 25245 33284 25279
rect 33232 25236 33284 25245
rect 31852 25100 31904 25152
rect 33508 25100 33560 25152
rect 36268 25100 36320 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9128 24896 9180 24948
rect 2780 24871 2832 24880
rect 2780 24837 2789 24871
rect 2789 24837 2823 24871
rect 2823 24837 2832 24871
rect 2780 24828 2832 24837
rect 9772 24828 9824 24880
rect 2596 24803 2648 24812
rect 2596 24769 2605 24803
rect 2605 24769 2639 24803
rect 2639 24769 2648 24803
rect 2596 24760 2648 24769
rect 5080 24760 5132 24812
rect 10048 24803 10100 24812
rect 3056 24735 3108 24744
rect 3056 24701 3065 24735
rect 3065 24701 3099 24735
rect 3099 24701 3108 24735
rect 3056 24692 3108 24701
rect 10048 24769 10057 24803
rect 10057 24769 10091 24803
rect 10091 24769 10100 24803
rect 10048 24760 10100 24769
rect 10140 24760 10192 24812
rect 10232 24735 10284 24744
rect 10232 24701 10241 24735
rect 10241 24701 10275 24735
rect 10275 24701 10284 24735
rect 10232 24692 10284 24701
rect 21732 24828 21784 24880
rect 21916 24828 21968 24880
rect 25412 24871 25464 24880
rect 25412 24837 25421 24871
rect 25421 24837 25455 24871
rect 25455 24837 25464 24871
rect 25412 24828 25464 24837
rect 16672 24760 16724 24812
rect 20168 24760 20220 24812
rect 23020 24803 23072 24812
rect 23020 24769 23029 24803
rect 23029 24769 23063 24803
rect 23063 24769 23072 24803
rect 23020 24760 23072 24769
rect 15292 24692 15344 24744
rect 15660 24735 15712 24744
rect 15660 24701 15669 24735
rect 15669 24701 15703 24735
rect 15703 24701 15712 24735
rect 15660 24692 15712 24701
rect 15844 24735 15896 24744
rect 15844 24701 15853 24735
rect 15853 24701 15887 24735
rect 15887 24701 15896 24735
rect 15844 24692 15896 24701
rect 20352 24735 20404 24744
rect 20352 24701 20361 24735
rect 20361 24701 20395 24735
rect 20395 24701 20404 24735
rect 20352 24692 20404 24701
rect 21640 24692 21692 24744
rect 22928 24692 22980 24744
rect 23480 24735 23532 24744
rect 23480 24701 23489 24735
rect 23489 24701 23523 24735
rect 23523 24701 23532 24735
rect 23480 24692 23532 24701
rect 24952 24692 25004 24744
rect 25688 24803 25740 24812
rect 25688 24769 25697 24803
rect 25697 24769 25731 24803
rect 25731 24769 25740 24803
rect 25688 24760 25740 24769
rect 26056 24760 26108 24812
rect 29920 24828 29972 24880
rect 30656 24803 30708 24812
rect 30656 24769 30665 24803
rect 30665 24769 30699 24803
rect 30699 24769 30708 24803
rect 30656 24760 30708 24769
rect 30932 24760 30984 24812
rect 33600 24760 33652 24812
rect 25596 24692 25648 24744
rect 26148 24692 26200 24744
rect 3424 24556 3476 24608
rect 4896 24556 4948 24608
rect 5816 24556 5868 24608
rect 10324 24599 10376 24608
rect 10324 24565 10333 24599
rect 10333 24565 10367 24599
rect 10367 24565 10376 24599
rect 10324 24556 10376 24565
rect 21824 24599 21876 24608
rect 21824 24565 21833 24599
rect 21833 24565 21867 24599
rect 21867 24565 21876 24599
rect 21824 24556 21876 24565
rect 26608 24624 26660 24676
rect 23664 24556 23716 24608
rect 25412 24599 25464 24608
rect 25412 24565 25421 24599
rect 25421 24565 25455 24599
rect 25455 24565 25464 24599
rect 25412 24556 25464 24565
rect 26240 24556 26292 24608
rect 27068 24735 27120 24744
rect 27068 24701 27077 24735
rect 27077 24701 27111 24735
rect 27111 24701 27120 24735
rect 27068 24692 27120 24701
rect 29000 24692 29052 24744
rect 29644 24735 29696 24744
rect 29644 24701 29653 24735
rect 29653 24701 29687 24735
rect 29687 24701 29696 24735
rect 29644 24692 29696 24701
rect 29920 24735 29972 24744
rect 29920 24701 29929 24735
rect 29929 24701 29963 24735
rect 29963 24701 29972 24735
rect 29920 24692 29972 24701
rect 27712 24624 27764 24676
rect 31668 24624 31720 24676
rect 33232 24624 33284 24676
rect 30564 24556 30616 24608
rect 30840 24556 30892 24608
rect 31116 24556 31168 24608
rect 31852 24556 31904 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2872 24352 2924 24404
rect 3240 24352 3292 24404
rect 5080 24352 5132 24404
rect 15844 24352 15896 24404
rect 17132 24395 17184 24404
rect 3056 24284 3108 24336
rect 9772 24284 9824 24336
rect 4620 24216 4672 24268
rect 4896 24216 4948 24268
rect 15660 24216 15712 24268
rect 17132 24361 17141 24395
rect 17141 24361 17175 24395
rect 17175 24361 17184 24395
rect 17132 24352 17184 24361
rect 18144 24395 18196 24404
rect 18144 24361 18153 24395
rect 18153 24361 18187 24395
rect 18187 24361 18196 24395
rect 18144 24352 18196 24361
rect 19248 24352 19300 24404
rect 22928 24395 22980 24404
rect 22928 24361 22937 24395
rect 22937 24361 22971 24395
rect 22971 24361 22980 24395
rect 22928 24352 22980 24361
rect 25412 24352 25464 24404
rect 26976 24352 27028 24404
rect 30656 24352 30708 24404
rect 36636 24352 36688 24404
rect 23480 24284 23532 24336
rect 16396 24216 16448 24268
rect 16948 24259 17000 24268
rect 16948 24225 16957 24259
rect 16957 24225 16991 24259
rect 16991 24225 17000 24259
rect 16948 24216 17000 24225
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 4804 24148 4856 24200
rect 5448 24148 5500 24200
rect 6644 24148 6696 24200
rect 16856 24191 16908 24200
rect 16856 24157 16865 24191
rect 16865 24157 16899 24191
rect 16899 24157 16908 24191
rect 16856 24148 16908 24157
rect 18512 24148 18564 24200
rect 4712 24080 4764 24132
rect 4620 24012 4672 24064
rect 16672 24080 16724 24132
rect 17316 24080 17368 24132
rect 21640 24216 21692 24268
rect 23112 24216 23164 24268
rect 25688 24216 25740 24268
rect 19984 24148 20036 24200
rect 20352 24148 20404 24200
rect 21824 24148 21876 24200
rect 22008 24148 22060 24200
rect 23664 24191 23716 24200
rect 23664 24157 23673 24191
rect 23673 24157 23707 24191
rect 23707 24157 23716 24191
rect 23664 24148 23716 24157
rect 24308 24148 24360 24200
rect 29920 24216 29972 24268
rect 32312 24259 32364 24268
rect 32312 24225 32321 24259
rect 32321 24225 32355 24259
rect 32355 24225 32364 24259
rect 32312 24216 32364 24225
rect 33600 24216 33652 24268
rect 26608 24191 26660 24200
rect 22468 24080 22520 24132
rect 25228 24080 25280 24132
rect 26608 24157 26617 24191
rect 26617 24157 26651 24191
rect 26651 24157 26660 24191
rect 26608 24148 26660 24157
rect 27068 24148 27120 24200
rect 32680 24148 32732 24200
rect 33508 24191 33560 24200
rect 33508 24157 33517 24191
rect 33517 24157 33551 24191
rect 33551 24157 33560 24191
rect 33508 24148 33560 24157
rect 26240 24080 26292 24132
rect 26976 24080 27028 24132
rect 19248 24055 19300 24064
rect 19248 24021 19257 24055
rect 19257 24021 19291 24055
rect 19291 24021 19300 24055
rect 19248 24012 19300 24021
rect 29828 24012 29880 24064
rect 34336 24012 34388 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 16856 23808 16908 23860
rect 17224 23808 17276 23860
rect 4988 23672 5040 23724
rect 5264 23672 5316 23724
rect 5448 23672 5500 23724
rect 6736 23672 6788 23724
rect 16856 23715 16908 23724
rect 16856 23681 16872 23715
rect 16872 23681 16906 23715
rect 16906 23681 16908 23715
rect 16856 23672 16908 23681
rect 16948 23647 17000 23656
rect 16948 23613 16957 23647
rect 16957 23613 16991 23647
rect 16991 23613 17000 23647
rect 16948 23604 17000 23613
rect 17040 23604 17092 23656
rect 17316 23672 17368 23724
rect 18236 23740 18288 23792
rect 19248 23740 19300 23792
rect 23664 23808 23716 23860
rect 25228 23808 25280 23860
rect 26056 23808 26108 23860
rect 29828 23783 29880 23792
rect 18052 23604 18104 23656
rect 7748 23536 7800 23588
rect 18972 23672 19024 23724
rect 20168 23672 20220 23724
rect 20352 23715 20404 23724
rect 20352 23681 20361 23715
rect 20361 23681 20395 23715
rect 20395 23681 20404 23715
rect 20352 23672 20404 23681
rect 29828 23749 29837 23783
rect 29837 23749 29871 23783
rect 29871 23749 29880 23783
rect 29828 23740 29880 23749
rect 22928 23672 22980 23724
rect 23388 23715 23440 23724
rect 23388 23681 23397 23715
rect 23397 23681 23431 23715
rect 23431 23681 23440 23715
rect 23388 23672 23440 23681
rect 4712 23468 4764 23520
rect 12900 23468 12952 23520
rect 15292 23511 15344 23520
rect 15292 23477 15301 23511
rect 15301 23477 15335 23511
rect 15335 23477 15344 23511
rect 15292 23468 15344 23477
rect 16028 23468 16080 23520
rect 17132 23511 17184 23520
rect 17132 23477 17141 23511
rect 17141 23477 17175 23511
rect 17175 23477 17184 23511
rect 17132 23468 17184 23477
rect 19156 23604 19208 23656
rect 19248 23604 19300 23656
rect 22468 23604 22520 23656
rect 26240 23672 26292 23724
rect 30656 23672 30708 23724
rect 34336 23715 34388 23724
rect 34336 23681 34345 23715
rect 34345 23681 34379 23715
rect 34379 23681 34388 23715
rect 34336 23672 34388 23681
rect 18512 23536 18564 23588
rect 18972 23536 19024 23588
rect 24860 23647 24912 23656
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 28172 23647 28224 23656
rect 28172 23613 28181 23647
rect 28181 23613 28215 23647
rect 28215 23613 28224 23647
rect 28172 23604 28224 23613
rect 19156 23468 19208 23520
rect 23112 23511 23164 23520
rect 23112 23477 23121 23511
rect 23121 23477 23155 23511
rect 23155 23477 23164 23511
rect 23112 23468 23164 23477
rect 27068 23511 27120 23520
rect 27068 23477 27077 23511
rect 27077 23477 27111 23511
rect 27111 23477 27120 23511
rect 27068 23468 27120 23477
rect 30472 23511 30524 23520
rect 30472 23477 30481 23511
rect 30481 23477 30515 23511
rect 30515 23477 30524 23511
rect 30472 23468 30524 23477
rect 32680 23511 32732 23520
rect 32680 23477 32689 23511
rect 32689 23477 32723 23511
rect 32723 23477 32732 23511
rect 32680 23468 32732 23477
rect 34520 23511 34572 23520
rect 34520 23477 34529 23511
rect 34529 23477 34563 23511
rect 34563 23477 34572 23511
rect 34520 23468 34572 23477
rect 34796 23468 34848 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4804 23264 4856 23316
rect 6644 23307 6696 23316
rect 6644 23273 6653 23307
rect 6653 23273 6687 23307
rect 6687 23273 6696 23307
rect 6644 23264 6696 23273
rect 12532 23307 12584 23316
rect 12532 23273 12541 23307
rect 12541 23273 12575 23307
rect 12575 23273 12584 23307
rect 12532 23264 12584 23273
rect 13268 23307 13320 23316
rect 13268 23273 13277 23307
rect 13277 23273 13311 23307
rect 13311 23273 13320 23307
rect 13268 23264 13320 23273
rect 18144 23264 18196 23316
rect 19248 23264 19300 23316
rect 20352 23307 20404 23316
rect 20352 23273 20361 23307
rect 20361 23273 20395 23307
rect 20395 23273 20404 23307
rect 20352 23264 20404 23273
rect 36084 23264 36136 23316
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2780 23060 2832 23112
rect 19984 23196 20036 23248
rect 4620 23128 4672 23180
rect 9220 23128 9272 23180
rect 15292 23128 15344 23180
rect 17684 23171 17736 23180
rect 17684 23137 17693 23171
rect 17693 23137 17727 23171
rect 17727 23137 17736 23171
rect 17684 23128 17736 23137
rect 24492 23128 24544 23180
rect 24860 23128 24912 23180
rect 29736 23128 29788 23180
rect 30932 23128 30984 23180
rect 4160 23103 4212 23112
rect 4160 23069 4169 23103
rect 4169 23069 4203 23103
rect 4203 23069 4212 23103
rect 4160 23060 4212 23069
rect 4988 23060 5040 23112
rect 10876 23103 10928 23112
rect 10876 23069 10885 23103
rect 10885 23069 10919 23103
rect 10919 23069 10928 23103
rect 10876 23060 10928 23069
rect 11336 23103 11388 23112
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 12900 23060 12952 23112
rect 14004 23060 14056 23112
rect 18236 23103 18288 23112
rect 4712 22992 4764 23044
rect 7840 23035 7892 23044
rect 7840 23001 7849 23035
rect 7849 23001 7883 23035
rect 7883 23001 7892 23035
rect 7840 22992 7892 23001
rect 15292 22992 15344 23044
rect 16672 23035 16724 23044
rect 16672 23001 16681 23035
rect 16681 23001 16715 23035
rect 16715 23001 16724 23035
rect 16672 22992 16724 23001
rect 18236 23069 18245 23103
rect 18245 23069 18279 23103
rect 18279 23069 18288 23103
rect 18236 23060 18288 23069
rect 18512 23103 18564 23112
rect 18512 23069 18521 23103
rect 18521 23069 18555 23103
rect 18555 23069 18564 23103
rect 18512 23060 18564 23069
rect 20168 23060 20220 23112
rect 29920 23103 29972 23112
rect 29920 23069 29929 23103
rect 29929 23069 29963 23103
rect 29963 23069 29972 23103
rect 29920 23060 29972 23069
rect 30840 23103 30892 23112
rect 30840 23069 30849 23103
rect 30849 23069 30883 23103
rect 30883 23069 30892 23103
rect 30840 23060 30892 23069
rect 33876 23060 33928 23112
rect 34796 23103 34848 23112
rect 34796 23069 34805 23103
rect 34805 23069 34839 23103
rect 34839 23069 34848 23103
rect 34796 23060 34848 23069
rect 18972 22992 19024 23044
rect 25964 22992 26016 23044
rect 1584 22967 1636 22976
rect 1584 22933 1593 22967
rect 1593 22933 1627 22967
rect 1627 22933 1636 22967
rect 1584 22924 1636 22933
rect 2964 22924 3016 22976
rect 16856 22924 16908 22976
rect 19432 22924 19484 22976
rect 20812 22924 20864 22976
rect 22928 22967 22980 22976
rect 22928 22933 22937 22967
rect 22937 22933 22971 22967
rect 22971 22933 22980 22967
rect 22928 22924 22980 22933
rect 25228 22967 25280 22976
rect 25228 22933 25237 22967
rect 25237 22933 25271 22967
rect 25271 22933 25280 22967
rect 25228 22924 25280 22933
rect 30104 22967 30156 22976
rect 30104 22933 30113 22967
rect 30113 22933 30147 22967
rect 30147 22933 30156 22967
rect 30104 22924 30156 22933
rect 31484 22967 31536 22976
rect 31484 22933 31493 22967
rect 31493 22933 31527 22967
rect 31527 22933 31536 22967
rect 31484 22924 31536 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4160 22720 4212 22772
rect 7840 22720 7892 22772
rect 8208 22720 8260 22772
rect 25228 22720 25280 22772
rect 29920 22763 29972 22772
rect 29920 22729 29929 22763
rect 29929 22729 29963 22763
rect 29963 22729 29972 22763
rect 29920 22720 29972 22729
rect 30564 22720 30616 22772
rect 33692 22720 33744 22772
rect 33876 22763 33928 22772
rect 33876 22729 33885 22763
rect 33885 22729 33919 22763
rect 33919 22729 33928 22763
rect 33876 22720 33928 22729
rect 1400 22695 1452 22704
rect 1400 22661 1409 22695
rect 1409 22661 1443 22695
rect 1443 22661 1452 22695
rect 1400 22652 1452 22661
rect 2964 22695 3016 22704
rect 2964 22661 2973 22695
rect 2973 22661 3007 22695
rect 3007 22661 3016 22695
rect 2964 22652 3016 22661
rect 7656 22695 7708 22704
rect 7656 22661 7665 22695
rect 7665 22661 7699 22695
rect 7699 22661 7708 22695
rect 7656 22652 7708 22661
rect 2780 22627 2832 22636
rect 2780 22593 2789 22627
rect 2789 22593 2823 22627
rect 2823 22593 2832 22627
rect 2780 22584 2832 22593
rect 5264 22627 5316 22636
rect 5264 22593 5273 22627
rect 5273 22593 5307 22627
rect 5307 22593 5316 22627
rect 5264 22584 5316 22593
rect 6644 22584 6696 22636
rect 9404 22584 9456 22636
rect 12348 22584 12400 22636
rect 3240 22559 3292 22568
rect 3240 22525 3249 22559
rect 3249 22525 3283 22559
rect 3283 22525 3292 22559
rect 9864 22559 9916 22568
rect 3240 22516 3292 22525
rect 9864 22525 9873 22559
rect 9873 22525 9907 22559
rect 9907 22525 9916 22559
rect 9864 22516 9916 22525
rect 12532 22516 12584 22568
rect 11520 22448 11572 22500
rect 5080 22423 5132 22432
rect 5080 22389 5089 22423
rect 5089 22389 5123 22423
rect 5123 22389 5132 22423
rect 5080 22380 5132 22389
rect 5816 22423 5868 22432
rect 5816 22389 5825 22423
rect 5825 22389 5859 22423
rect 5859 22389 5868 22423
rect 5816 22380 5868 22389
rect 7104 22423 7156 22432
rect 7104 22389 7113 22423
rect 7113 22389 7147 22423
rect 7147 22389 7156 22423
rect 7104 22380 7156 22389
rect 11704 22423 11756 22432
rect 11704 22389 11713 22423
rect 11713 22389 11747 22423
rect 11747 22389 11756 22423
rect 11704 22380 11756 22389
rect 18236 22652 18288 22704
rect 16028 22627 16080 22636
rect 16028 22593 16037 22627
rect 16037 22593 16071 22627
rect 16071 22593 16080 22627
rect 16028 22584 16080 22593
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 18512 22584 18564 22636
rect 19432 22584 19484 22636
rect 20812 22627 20864 22636
rect 20812 22593 20821 22627
rect 20821 22593 20855 22627
rect 20855 22593 20864 22627
rect 20812 22584 20864 22593
rect 22468 22584 22520 22636
rect 22928 22584 22980 22636
rect 23388 22652 23440 22704
rect 18052 22559 18104 22568
rect 18052 22525 18061 22559
rect 18061 22525 18095 22559
rect 18095 22525 18104 22559
rect 18052 22516 18104 22525
rect 18236 22516 18288 22568
rect 18972 22559 19024 22568
rect 18972 22525 18981 22559
rect 18981 22525 19015 22559
rect 19015 22525 19024 22559
rect 18972 22516 19024 22525
rect 16672 22491 16724 22500
rect 16672 22457 16681 22491
rect 16681 22457 16715 22491
rect 16715 22457 16724 22491
rect 16672 22448 16724 22457
rect 14004 22380 14056 22432
rect 14924 22380 14976 22432
rect 15200 22380 15252 22432
rect 17684 22423 17736 22432
rect 17684 22389 17693 22423
rect 17693 22389 17727 22423
rect 17727 22389 17736 22423
rect 17684 22380 17736 22389
rect 18144 22423 18196 22432
rect 18144 22389 18153 22423
rect 18153 22389 18187 22423
rect 18187 22389 18196 22423
rect 18144 22380 18196 22389
rect 18604 22423 18656 22432
rect 18604 22389 18613 22423
rect 18613 22389 18647 22423
rect 18647 22389 18656 22423
rect 18604 22380 18656 22389
rect 27436 22627 27488 22636
rect 27436 22593 27445 22627
rect 27445 22593 27479 22627
rect 27479 22593 27488 22627
rect 27436 22584 27488 22593
rect 30932 22652 30984 22704
rect 34520 22652 34572 22704
rect 29736 22627 29788 22636
rect 29736 22593 29745 22627
rect 29745 22593 29779 22627
rect 29779 22593 29788 22627
rect 29736 22584 29788 22593
rect 30012 22584 30064 22636
rect 30288 22584 30340 22636
rect 32956 22584 33008 22636
rect 30472 22559 30524 22568
rect 30472 22525 30481 22559
rect 30481 22525 30515 22559
rect 30515 22525 30524 22559
rect 30472 22516 30524 22525
rect 34612 22584 34664 22636
rect 19432 22380 19484 22432
rect 20352 22380 20404 22432
rect 23112 22423 23164 22432
rect 23112 22389 23121 22423
rect 23121 22389 23155 22423
rect 23155 22389 23164 22423
rect 23112 22380 23164 22389
rect 30748 22448 30800 22500
rect 33784 22448 33836 22500
rect 34796 22516 34848 22568
rect 23480 22380 23532 22432
rect 27528 22380 27580 22432
rect 28172 22380 28224 22432
rect 30012 22380 30064 22432
rect 34520 22380 34572 22432
rect 36268 22423 36320 22432
rect 36268 22389 36277 22423
rect 36277 22389 36311 22423
rect 36311 22389 36320 22423
rect 36268 22380 36320 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 5264 22176 5316 22228
rect 6644 22176 6696 22228
rect 7380 22176 7432 22228
rect 9404 22176 9456 22228
rect 29736 22176 29788 22228
rect 4804 22108 4856 22160
rect 4620 22040 4672 22092
rect 8392 22040 8444 22092
rect 12532 22108 12584 22160
rect 15292 22108 15344 22160
rect 11336 22040 11388 22092
rect 11428 22040 11480 22092
rect 12624 22083 12676 22092
rect 12624 22049 12633 22083
rect 12633 22049 12667 22083
rect 12667 22049 12676 22083
rect 12624 22040 12676 22049
rect 14924 22083 14976 22092
rect 14924 22049 14933 22083
rect 14933 22049 14967 22083
rect 14967 22049 14976 22083
rect 14924 22040 14976 22049
rect 15200 22040 15252 22092
rect 18052 22040 18104 22092
rect 18420 22040 18472 22092
rect 20352 22083 20404 22092
rect 20352 22049 20361 22083
rect 20361 22049 20395 22083
rect 20395 22049 20404 22083
rect 20352 22040 20404 22049
rect 20444 22040 20496 22092
rect 27620 22083 27672 22092
rect 27620 22049 27629 22083
rect 27629 22049 27663 22083
rect 27663 22049 27672 22083
rect 27620 22040 27672 22049
rect 31024 22040 31076 22092
rect 34520 22040 34572 22092
rect 2688 22015 2740 22024
rect 2688 21981 2697 22015
rect 2697 21981 2731 22015
rect 2731 21981 2740 22015
rect 2688 21972 2740 21981
rect 4252 22015 4304 22024
rect 4252 21981 4261 22015
rect 4261 21981 4295 22015
rect 4295 21981 4304 22015
rect 4252 21972 4304 21981
rect 4988 22015 5040 22024
rect 4988 21981 4997 22015
rect 4997 21981 5031 22015
rect 5031 21981 5040 22015
rect 4988 21972 5040 21981
rect 5816 21972 5868 22024
rect 7104 21972 7156 22024
rect 7656 22015 7708 22024
rect 7656 21981 7665 22015
rect 7665 21981 7699 22015
rect 7699 21981 7708 22015
rect 7656 21972 7708 21981
rect 4712 21904 4764 21956
rect 9588 21972 9640 22024
rect 11336 21947 11388 21956
rect 4620 21836 4672 21888
rect 7380 21836 7432 21888
rect 7840 21879 7892 21888
rect 7840 21845 7849 21879
rect 7849 21845 7883 21879
rect 7883 21845 7892 21879
rect 7840 21836 7892 21845
rect 9772 21836 9824 21888
rect 9864 21836 9916 21888
rect 10600 21879 10652 21888
rect 10600 21845 10609 21879
rect 10609 21845 10643 21879
rect 10643 21845 10652 21879
rect 10600 21836 10652 21845
rect 11336 21913 11345 21947
rect 11345 21913 11379 21947
rect 11379 21913 11388 21947
rect 11336 21904 11388 21913
rect 11428 21904 11480 21956
rect 18052 21904 18104 21956
rect 13544 21879 13596 21888
rect 13544 21845 13553 21879
rect 13553 21845 13587 21879
rect 13587 21845 13596 21879
rect 13544 21836 13596 21845
rect 13820 21836 13872 21888
rect 15108 21836 15160 21888
rect 18236 21879 18288 21888
rect 18236 21845 18245 21879
rect 18245 21845 18279 21879
rect 18279 21845 18288 21879
rect 18236 21836 18288 21845
rect 23572 22015 23624 22024
rect 23572 21981 23581 22015
rect 23581 21981 23615 22015
rect 23615 21981 23624 22015
rect 23572 21972 23624 21981
rect 30932 21972 30984 22024
rect 32128 21972 32180 22024
rect 33692 21972 33744 22024
rect 35808 21972 35860 22024
rect 24952 21904 25004 21956
rect 25964 21947 26016 21956
rect 25964 21913 25973 21947
rect 25973 21913 26007 21947
rect 26007 21913 26016 21947
rect 25964 21904 26016 21913
rect 31484 21904 31536 21956
rect 33968 21947 34020 21956
rect 33968 21913 33977 21947
rect 33977 21913 34011 21947
rect 34011 21913 34020 21947
rect 33968 21904 34020 21913
rect 22468 21879 22520 21888
rect 22468 21845 22477 21879
rect 22477 21845 22511 21879
rect 22511 21845 22520 21879
rect 22468 21836 22520 21845
rect 29644 21836 29696 21888
rect 31760 21836 31812 21888
rect 31944 21836 31996 21888
rect 32312 21836 32364 21888
rect 36636 21836 36688 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4160 21632 4212 21684
rect 5080 21564 5132 21616
rect 5172 21564 5224 21616
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 2688 21539 2740 21548
rect 2688 21505 2697 21539
rect 2697 21505 2731 21539
rect 2731 21505 2740 21539
rect 2688 21496 2740 21505
rect 4528 21539 4580 21548
rect 4528 21505 4537 21539
rect 4537 21505 4571 21539
rect 4571 21505 4580 21539
rect 4528 21496 4580 21505
rect 5448 21539 5500 21548
rect 5448 21505 5457 21539
rect 5457 21505 5491 21539
rect 5491 21505 5500 21539
rect 5448 21496 5500 21505
rect 9772 21632 9824 21684
rect 9956 21632 10008 21684
rect 10232 21632 10284 21684
rect 10692 21675 10744 21684
rect 10692 21641 10701 21675
rect 10701 21641 10735 21675
rect 10735 21641 10744 21675
rect 10692 21632 10744 21641
rect 13544 21632 13596 21684
rect 22468 21632 22520 21684
rect 30932 21632 30984 21684
rect 31944 21632 31996 21684
rect 32128 21675 32180 21684
rect 32128 21641 32137 21675
rect 32137 21641 32171 21675
rect 32171 21641 32180 21675
rect 32128 21632 32180 21641
rect 35808 21632 35860 21684
rect 38016 21675 38068 21684
rect 38016 21641 38025 21675
rect 38025 21641 38059 21675
rect 38059 21641 38068 21675
rect 38016 21632 38068 21641
rect 11704 21607 11756 21616
rect 11704 21573 11713 21607
rect 11713 21573 11747 21607
rect 11747 21573 11756 21607
rect 11704 21564 11756 21573
rect 12440 21564 12492 21616
rect 18236 21564 18288 21616
rect 19432 21564 19484 21616
rect 23572 21564 23624 21616
rect 4988 21428 5040 21480
rect 5356 21428 5408 21480
rect 9588 21496 9640 21548
rect 10876 21539 10928 21548
rect 10876 21505 10885 21539
rect 10885 21505 10919 21539
rect 10919 21505 10928 21539
rect 10876 21496 10928 21505
rect 11520 21539 11572 21548
rect 11520 21505 11529 21539
rect 11529 21505 11563 21539
rect 11563 21505 11572 21539
rect 11520 21496 11572 21505
rect 13820 21539 13872 21548
rect 13820 21505 13829 21539
rect 13829 21505 13863 21539
rect 13863 21505 13872 21539
rect 13820 21496 13872 21505
rect 14004 21496 14056 21548
rect 17684 21496 17736 21548
rect 30104 21564 30156 21616
rect 25964 21539 26016 21548
rect 25964 21505 25973 21539
rect 25973 21505 26007 21539
rect 26007 21505 26016 21539
rect 25964 21496 26016 21505
rect 7380 21428 7432 21480
rect 9956 21428 10008 21480
rect 12532 21471 12584 21480
rect 12532 21437 12541 21471
rect 12541 21437 12575 21471
rect 12575 21437 12584 21471
rect 12532 21428 12584 21437
rect 17408 21471 17460 21480
rect 17408 21437 17417 21471
rect 17417 21437 17451 21471
rect 17451 21437 17460 21471
rect 17408 21428 17460 21437
rect 19708 21428 19760 21480
rect 12440 21360 12492 21412
rect 12624 21360 12676 21412
rect 20444 21428 20496 21480
rect 23664 21471 23716 21480
rect 23664 21437 23673 21471
rect 23673 21437 23707 21471
rect 23707 21437 23716 21471
rect 23664 21428 23716 21437
rect 25044 21471 25096 21480
rect 25044 21437 25053 21471
rect 25053 21437 25087 21471
rect 25087 21437 25096 21471
rect 25044 21428 25096 21437
rect 2504 21292 2556 21344
rect 5264 21335 5316 21344
rect 5264 21301 5273 21335
rect 5273 21301 5307 21335
rect 5307 21301 5316 21335
rect 5264 21292 5316 21301
rect 5356 21292 5408 21344
rect 7656 21292 7708 21344
rect 7932 21335 7984 21344
rect 7932 21301 7941 21335
rect 7941 21301 7975 21335
rect 7975 21301 7984 21335
rect 7932 21292 7984 21301
rect 13912 21292 13964 21344
rect 22744 21292 22796 21344
rect 26332 21292 26384 21344
rect 37832 21539 37884 21548
rect 37832 21505 37841 21539
rect 37841 21505 37875 21539
rect 37875 21505 37884 21539
rect 37832 21496 37884 21505
rect 31760 21292 31812 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 4804 21088 4856 21140
rect 5356 21088 5408 21140
rect 7840 21088 7892 21140
rect 11888 21131 11940 21140
rect 5172 21020 5224 21072
rect 5264 20995 5316 21004
rect 5264 20961 5273 20995
rect 5273 20961 5307 20995
rect 5307 20961 5316 20995
rect 5264 20952 5316 20961
rect 5540 20995 5592 21004
rect 5540 20961 5549 20995
rect 5549 20961 5583 20995
rect 5583 20961 5592 20995
rect 5540 20952 5592 20961
rect 11888 21097 11897 21131
rect 11897 21097 11931 21131
rect 11931 21097 11940 21131
rect 11888 21088 11940 21097
rect 12348 21131 12400 21140
rect 12348 21097 12357 21131
rect 12357 21097 12391 21131
rect 12391 21097 12400 21131
rect 12348 21088 12400 21097
rect 19708 21131 19760 21140
rect 19708 21097 19717 21131
rect 19717 21097 19751 21131
rect 19751 21097 19760 21131
rect 19708 21088 19760 21097
rect 24400 21131 24452 21140
rect 24400 21097 24409 21131
rect 24409 21097 24443 21131
rect 24443 21097 24452 21131
rect 24400 21088 24452 21097
rect 25044 21088 25096 21140
rect 26332 21088 26384 21140
rect 29552 21088 29604 21140
rect 29920 21131 29972 21140
rect 29920 21097 29929 21131
rect 29929 21097 29963 21131
rect 29963 21097 29972 21131
rect 29920 21088 29972 21097
rect 30840 21088 30892 21140
rect 9956 21020 10008 21072
rect 24308 21020 24360 21072
rect 9404 20952 9456 21004
rect 10692 20952 10744 21004
rect 18604 20952 18656 21004
rect 24492 20995 24544 21004
rect 24492 20961 24501 20995
rect 24501 20961 24535 20995
rect 24535 20961 24544 20995
rect 24492 20952 24544 20961
rect 29644 20952 29696 21004
rect 31024 20995 31076 21004
rect 31024 20961 31033 20995
rect 31033 20961 31067 20995
rect 31067 20961 31076 20995
rect 31024 20952 31076 20961
rect 4160 20884 4212 20936
rect 4620 20927 4672 20936
rect 4620 20893 4629 20927
rect 4629 20893 4663 20927
rect 4663 20893 4672 20927
rect 4620 20884 4672 20893
rect 5080 20927 5132 20936
rect 5080 20893 5089 20927
rect 5089 20893 5123 20927
rect 5123 20893 5132 20927
rect 5080 20884 5132 20893
rect 12716 20884 12768 20936
rect 12900 20927 12952 20936
rect 12900 20893 12909 20927
rect 12909 20893 12943 20927
rect 12943 20893 12952 20927
rect 12900 20884 12952 20893
rect 13268 20884 13320 20936
rect 16304 20927 16356 20936
rect 16304 20893 16313 20927
rect 16313 20893 16347 20927
rect 16347 20893 16356 20927
rect 16304 20884 16356 20893
rect 16948 20884 17000 20936
rect 22468 20884 22520 20936
rect 23940 20884 23992 20936
rect 24584 20884 24636 20936
rect 5264 20816 5316 20868
rect 9772 20816 9824 20868
rect 4160 20791 4212 20800
rect 4160 20757 4169 20791
rect 4169 20757 4203 20791
rect 4203 20757 4212 20791
rect 4160 20748 4212 20757
rect 11796 20748 11848 20800
rect 13084 20791 13136 20800
rect 13084 20757 13093 20791
rect 13093 20757 13127 20791
rect 13127 20757 13136 20791
rect 13084 20748 13136 20757
rect 31760 20884 31812 20936
rect 32588 20884 32640 20936
rect 27528 20816 27580 20868
rect 30932 20859 30984 20868
rect 30932 20825 30941 20859
rect 30941 20825 30975 20859
rect 30975 20825 30984 20859
rect 30932 20816 30984 20825
rect 25320 20748 25372 20800
rect 25964 20791 26016 20800
rect 25964 20757 25973 20791
rect 25973 20757 26007 20791
rect 26007 20757 26016 20791
rect 25964 20748 26016 20757
rect 29920 20748 29972 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5448 20587 5500 20596
rect 5448 20553 5457 20587
rect 5457 20553 5491 20587
rect 5491 20553 5500 20587
rect 5448 20544 5500 20553
rect 11336 20544 11388 20596
rect 12716 20587 12768 20596
rect 12716 20553 12725 20587
rect 12725 20553 12759 20587
rect 12759 20553 12768 20587
rect 12716 20544 12768 20553
rect 4068 20476 4120 20528
rect 5540 20476 5592 20528
rect 7656 20519 7708 20528
rect 7656 20485 7665 20519
rect 7665 20485 7699 20519
rect 7699 20485 7708 20519
rect 7656 20476 7708 20485
rect 1400 20451 1452 20460
rect 1400 20417 1409 20451
rect 1409 20417 1443 20451
rect 1443 20417 1452 20451
rect 1400 20408 1452 20417
rect 4160 20408 4212 20460
rect 4620 20408 4672 20460
rect 5172 20451 5224 20460
rect 5172 20417 5181 20451
rect 5181 20417 5215 20451
rect 5215 20417 5224 20451
rect 5172 20408 5224 20417
rect 5264 20451 5316 20460
rect 5264 20417 5273 20451
rect 5273 20417 5307 20451
rect 5307 20417 5316 20451
rect 11796 20451 11848 20460
rect 5264 20408 5316 20417
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 13084 20408 13136 20460
rect 17408 20476 17460 20528
rect 16304 20408 16356 20460
rect 7932 20340 7984 20392
rect 5540 20272 5592 20324
rect 14924 20340 14976 20392
rect 23940 20476 23992 20528
rect 24584 20408 24636 20460
rect 27528 20544 27580 20596
rect 23296 20340 23348 20392
rect 24308 20383 24360 20392
rect 2320 20204 2372 20256
rect 2596 20204 2648 20256
rect 5356 20204 5408 20256
rect 9680 20272 9732 20324
rect 19616 20272 19668 20324
rect 12624 20204 12676 20256
rect 13268 20204 13320 20256
rect 19340 20204 19392 20256
rect 19984 20204 20036 20256
rect 22100 20204 22152 20256
rect 23480 20204 23532 20256
rect 24308 20349 24317 20383
rect 24317 20349 24351 20383
rect 24351 20349 24360 20383
rect 24308 20340 24360 20349
rect 24400 20247 24452 20256
rect 24400 20213 24409 20247
rect 24409 20213 24443 20247
rect 24443 20213 24452 20247
rect 24400 20204 24452 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 5080 20000 5132 20052
rect 7840 20000 7892 20052
rect 24400 20043 24452 20052
rect 24400 20009 24409 20043
rect 24409 20009 24443 20043
rect 24443 20009 24452 20043
rect 24400 20000 24452 20009
rect 35992 20043 36044 20052
rect 35992 20009 36001 20043
rect 36001 20009 36035 20043
rect 36035 20009 36044 20043
rect 35992 20000 36044 20009
rect 37004 20000 37056 20052
rect 13912 19932 13964 19984
rect 20904 19932 20956 19984
rect 27436 19932 27488 19984
rect 12624 19864 12676 19916
rect 14924 19907 14976 19916
rect 14924 19873 14933 19907
rect 14933 19873 14967 19907
rect 14967 19873 14976 19907
rect 14924 19864 14976 19873
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 17960 19907 18012 19916
rect 17960 19873 17969 19907
rect 17969 19873 18003 19907
rect 18003 19873 18012 19907
rect 17960 19864 18012 19873
rect 24308 19864 24360 19916
rect 36820 19864 36872 19916
rect 2412 19839 2464 19848
rect 2412 19805 2421 19839
rect 2421 19805 2455 19839
rect 2455 19805 2464 19839
rect 2412 19796 2464 19805
rect 7288 19839 7340 19848
rect 7288 19805 7297 19839
rect 7297 19805 7331 19839
rect 7331 19805 7340 19839
rect 7288 19796 7340 19805
rect 14464 19839 14516 19848
rect 11888 19728 11940 19780
rect 12348 19728 12400 19780
rect 14464 19805 14473 19839
rect 14473 19805 14507 19839
rect 14507 19805 14516 19839
rect 14464 19796 14516 19805
rect 16764 19839 16816 19848
rect 16764 19805 16773 19839
rect 16773 19805 16807 19839
rect 16807 19805 16816 19839
rect 16764 19796 16816 19805
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19616 19796 19668 19805
rect 22376 19796 22428 19848
rect 22744 19839 22796 19848
rect 22744 19805 22753 19839
rect 22753 19805 22787 19839
rect 22787 19805 22796 19839
rect 22744 19796 22796 19805
rect 23296 19796 23348 19848
rect 23940 19796 23992 19848
rect 24584 19796 24636 19848
rect 14648 19771 14700 19780
rect 14648 19737 14657 19771
rect 14657 19737 14691 19771
rect 14691 19737 14700 19771
rect 14648 19728 14700 19737
rect 20904 19703 20956 19712
rect 20904 19669 20913 19703
rect 20913 19669 20947 19703
rect 20947 19669 20956 19703
rect 20904 19660 20956 19669
rect 24584 19660 24636 19712
rect 28908 19796 28960 19848
rect 35992 19728 36044 19780
rect 36452 19703 36504 19712
rect 36452 19669 36461 19703
rect 36461 19669 36495 19703
rect 36495 19669 36504 19703
rect 36452 19660 36504 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 5172 19456 5224 19508
rect 8392 19499 8444 19508
rect 8392 19465 8401 19499
rect 8401 19465 8435 19499
rect 8435 19465 8444 19499
rect 8392 19456 8444 19465
rect 2596 19431 2648 19440
rect 2596 19397 2605 19431
rect 2605 19397 2639 19431
rect 2639 19397 2648 19431
rect 2596 19388 2648 19397
rect 6736 19388 6788 19440
rect 2412 19363 2464 19372
rect 2412 19329 2421 19363
rect 2421 19329 2455 19363
rect 2455 19329 2464 19363
rect 2412 19320 2464 19329
rect 5540 19363 5592 19372
rect 5540 19329 5549 19363
rect 5549 19329 5583 19363
rect 5583 19329 5592 19363
rect 5540 19320 5592 19329
rect 9864 19320 9916 19372
rect 18880 19388 18932 19440
rect 12808 19363 12860 19372
rect 12808 19329 12817 19363
rect 12817 19329 12851 19363
rect 12851 19329 12860 19363
rect 12808 19320 12860 19329
rect 14464 19363 14516 19372
rect 14464 19329 14473 19363
rect 14473 19329 14507 19363
rect 14507 19329 14516 19363
rect 14464 19320 14516 19329
rect 16764 19320 16816 19372
rect 2872 19295 2924 19304
rect 2872 19261 2881 19295
rect 2881 19261 2915 19295
rect 2915 19261 2924 19295
rect 2872 19252 2924 19261
rect 7380 19252 7432 19304
rect 10876 19184 10928 19236
rect 19892 19363 19944 19372
rect 19892 19329 19901 19363
rect 19901 19329 19935 19363
rect 19935 19329 19944 19363
rect 19892 19320 19944 19329
rect 23296 19431 23348 19440
rect 23296 19397 23305 19431
rect 23305 19397 23339 19431
rect 23339 19397 23348 19431
rect 23296 19388 23348 19397
rect 26424 19456 26476 19508
rect 29920 19456 29972 19508
rect 27068 19388 27120 19440
rect 27988 19388 28040 19440
rect 28908 19431 28960 19440
rect 28908 19397 28917 19431
rect 28917 19397 28951 19431
rect 28951 19397 28960 19431
rect 28908 19388 28960 19397
rect 22468 19363 22520 19372
rect 22468 19329 22477 19363
rect 22477 19329 22511 19363
rect 22511 19329 22520 19363
rect 22468 19320 22520 19329
rect 22652 19320 22704 19372
rect 23388 19320 23440 19372
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 24308 19363 24360 19372
rect 24308 19329 24317 19363
rect 24317 19329 24351 19363
rect 24351 19329 24360 19363
rect 24308 19320 24360 19329
rect 24584 19320 24636 19372
rect 32312 19363 32364 19372
rect 32312 19329 32321 19363
rect 32321 19329 32355 19363
rect 32355 19329 32364 19363
rect 32312 19320 32364 19329
rect 32496 19363 32548 19372
rect 32496 19329 32505 19363
rect 32505 19329 32539 19363
rect 32539 19329 32548 19363
rect 32496 19320 32548 19329
rect 35440 19320 35492 19372
rect 29828 19252 29880 19304
rect 20628 19184 20680 19236
rect 31668 19252 31720 19304
rect 31208 19184 31260 19236
rect 34520 19252 34572 19304
rect 7012 19159 7064 19168
rect 7012 19125 7021 19159
rect 7021 19125 7055 19159
rect 7055 19125 7064 19159
rect 7012 19116 7064 19125
rect 12532 19116 12584 19168
rect 13176 19116 13228 19168
rect 13452 19159 13504 19168
rect 13452 19125 13461 19159
rect 13461 19125 13495 19159
rect 13495 19125 13504 19159
rect 13452 19116 13504 19125
rect 18144 19159 18196 19168
rect 18144 19125 18153 19159
rect 18153 19125 18187 19159
rect 18187 19125 18196 19159
rect 18144 19116 18196 19125
rect 22100 19116 22152 19168
rect 22652 19159 22704 19168
rect 22652 19125 22661 19159
rect 22661 19125 22695 19159
rect 22695 19125 22704 19159
rect 22652 19116 22704 19125
rect 24400 19159 24452 19168
rect 24400 19125 24409 19159
rect 24409 19125 24443 19159
rect 24443 19125 24452 19159
rect 24400 19116 24452 19125
rect 32956 19116 33008 19168
rect 34796 19116 34848 19168
rect 35992 19116 36044 19168
rect 36084 19116 36136 19168
rect 36452 19116 36504 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 7288 18912 7340 18964
rect 12348 18912 12400 18964
rect 14648 18912 14700 18964
rect 20076 18912 20128 18964
rect 23296 18912 23348 18964
rect 24400 18955 24452 18964
rect 24400 18921 24409 18955
rect 24409 18921 24443 18955
rect 24443 18921 24452 18955
rect 24400 18912 24452 18921
rect 29736 18912 29788 18964
rect 30472 18912 30524 18964
rect 5172 18776 5224 18828
rect 7380 18776 7432 18828
rect 7748 18819 7800 18828
rect 7748 18785 7757 18819
rect 7757 18785 7791 18819
rect 7791 18785 7800 18819
rect 7748 18776 7800 18785
rect 12716 18776 12768 18828
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 5080 18751 5132 18760
rect 5080 18717 5089 18751
rect 5089 18717 5123 18751
rect 5123 18717 5132 18751
rect 5080 18708 5132 18717
rect 5724 18751 5776 18760
rect 5724 18717 5733 18751
rect 5733 18717 5767 18751
rect 5767 18717 5776 18751
rect 5724 18708 5776 18717
rect 7012 18708 7064 18760
rect 9128 18708 9180 18760
rect 10876 18708 10928 18760
rect 18144 18776 18196 18828
rect 4620 18640 4672 18692
rect 7472 18640 7524 18692
rect 8208 18640 8260 18692
rect 12532 18640 12584 18692
rect 2596 18572 2648 18624
rect 5632 18572 5684 18624
rect 5816 18572 5868 18624
rect 12440 18572 12492 18624
rect 17592 18751 17644 18760
rect 17592 18717 17601 18751
rect 17601 18717 17635 18751
rect 17635 18717 17644 18751
rect 17592 18708 17644 18717
rect 18420 18708 18472 18760
rect 18880 18708 18932 18760
rect 18972 18708 19024 18760
rect 19892 18776 19944 18828
rect 20720 18751 20772 18760
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 27620 18844 27672 18896
rect 34796 18912 34848 18964
rect 35440 18912 35492 18964
rect 36820 18955 36872 18964
rect 36820 18921 36829 18955
rect 36829 18921 36863 18955
rect 36863 18921 36872 18955
rect 36820 18912 36872 18921
rect 34520 18844 34572 18896
rect 24308 18776 24360 18828
rect 29552 18776 29604 18828
rect 36452 18776 36504 18828
rect 22744 18708 22796 18760
rect 24124 18708 24176 18760
rect 24584 18708 24636 18760
rect 19340 18572 19392 18624
rect 20628 18615 20680 18624
rect 20628 18581 20637 18615
rect 20637 18581 20671 18615
rect 20671 18581 20680 18615
rect 20628 18572 20680 18581
rect 21824 18615 21876 18624
rect 21824 18581 21833 18615
rect 21833 18581 21867 18615
rect 21867 18581 21876 18615
rect 21824 18572 21876 18581
rect 26424 18751 26476 18760
rect 26424 18717 26433 18751
rect 26433 18717 26467 18751
rect 26467 18717 26476 18751
rect 26424 18708 26476 18717
rect 29000 18751 29052 18760
rect 29000 18717 29009 18751
rect 29009 18717 29043 18751
rect 29043 18717 29052 18751
rect 29000 18708 29052 18717
rect 32588 18751 32640 18760
rect 32588 18717 32597 18751
rect 32597 18717 32631 18751
rect 32631 18717 32640 18751
rect 32588 18708 32640 18717
rect 25964 18615 26016 18624
rect 25964 18581 25973 18615
rect 25973 18581 26007 18615
rect 26007 18581 26016 18615
rect 25964 18572 26016 18581
rect 30840 18640 30892 18692
rect 31208 18640 31260 18692
rect 29828 18572 29880 18624
rect 32772 18708 32824 18760
rect 32956 18751 33008 18760
rect 32956 18717 32965 18751
rect 32965 18717 32999 18751
rect 32999 18717 33008 18751
rect 33784 18751 33836 18760
rect 32956 18708 33008 18717
rect 33784 18717 33793 18751
rect 33793 18717 33827 18751
rect 33827 18717 33836 18751
rect 33784 18708 33836 18717
rect 34612 18708 34664 18760
rect 35532 18708 35584 18760
rect 37924 18751 37976 18760
rect 37924 18717 37933 18751
rect 37933 18717 37967 18751
rect 37967 18717 37976 18751
rect 37924 18708 37976 18717
rect 35348 18640 35400 18692
rect 35808 18640 35860 18692
rect 36820 18640 36872 18692
rect 35440 18572 35492 18624
rect 36912 18572 36964 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2872 18368 2924 18420
rect 2320 18232 2372 18284
rect 4712 18275 4764 18284
rect 4712 18241 4721 18275
rect 4721 18241 4755 18275
rect 4755 18241 4764 18275
rect 4712 18232 4764 18241
rect 5724 18232 5776 18284
rect 5816 18275 5868 18284
rect 5816 18241 5825 18275
rect 5825 18241 5859 18275
rect 5859 18241 5868 18275
rect 7012 18300 7064 18352
rect 5816 18232 5868 18241
rect 7472 18232 7524 18284
rect 9128 18275 9180 18284
rect 5172 18164 5224 18216
rect 7380 18207 7432 18216
rect 7380 18173 7389 18207
rect 7389 18173 7423 18207
rect 7423 18173 7432 18207
rect 7380 18164 7432 18173
rect 5540 18096 5592 18148
rect 9128 18241 9137 18275
rect 9137 18241 9171 18275
rect 9171 18241 9180 18275
rect 9128 18232 9180 18241
rect 9588 18164 9640 18216
rect 13176 18343 13228 18352
rect 13176 18309 13185 18343
rect 13185 18309 13219 18343
rect 13219 18309 13228 18343
rect 13176 18300 13228 18309
rect 12716 18232 12768 18284
rect 12440 18164 12492 18216
rect 12624 18164 12676 18216
rect 13452 18164 13504 18216
rect 29828 18411 29880 18420
rect 18696 18300 18748 18352
rect 21824 18300 21876 18352
rect 17592 18275 17644 18284
rect 17592 18241 17601 18275
rect 17601 18241 17635 18275
rect 17635 18241 17644 18275
rect 17592 18232 17644 18241
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 25964 18300 26016 18352
rect 27804 18300 27856 18352
rect 28816 18343 28868 18352
rect 28816 18309 28825 18343
rect 28825 18309 28859 18343
rect 28859 18309 28868 18343
rect 28816 18300 28868 18309
rect 29828 18377 29837 18411
rect 29837 18377 29871 18411
rect 29871 18377 29880 18411
rect 29828 18368 29880 18377
rect 29920 18411 29972 18420
rect 29920 18377 29929 18411
rect 29929 18377 29963 18411
rect 29963 18377 29972 18411
rect 29920 18368 29972 18377
rect 32772 18411 32824 18420
rect 32772 18377 32781 18411
rect 32781 18377 32815 18411
rect 32815 18377 32824 18411
rect 32772 18368 32824 18377
rect 35348 18411 35400 18420
rect 35348 18377 35357 18411
rect 35357 18377 35391 18411
rect 35391 18377 35400 18411
rect 35348 18368 35400 18377
rect 35532 18368 35584 18420
rect 36084 18411 36136 18420
rect 36084 18377 36093 18411
rect 36093 18377 36127 18411
rect 36127 18377 36136 18411
rect 36084 18368 36136 18377
rect 37924 18368 37976 18420
rect 32312 18300 32364 18352
rect 32496 18300 32548 18352
rect 17960 18164 18012 18216
rect 18236 18207 18288 18216
rect 18236 18173 18245 18207
rect 18245 18173 18279 18207
rect 18279 18173 18288 18207
rect 18236 18164 18288 18173
rect 24400 18207 24452 18216
rect 24400 18173 24409 18207
rect 24409 18173 24443 18207
rect 24443 18173 24452 18207
rect 24400 18164 24452 18173
rect 27620 18164 27672 18216
rect 29736 18207 29788 18216
rect 29736 18173 29745 18207
rect 29745 18173 29779 18207
rect 29779 18173 29788 18207
rect 29736 18164 29788 18173
rect 31668 18164 31720 18216
rect 33968 18164 34020 18216
rect 34612 18232 34664 18284
rect 36912 18300 36964 18352
rect 35808 18232 35860 18284
rect 36452 18275 36504 18284
rect 36452 18241 36461 18275
rect 36461 18241 36495 18275
rect 36495 18241 36504 18275
rect 36452 18232 36504 18241
rect 36268 18164 36320 18216
rect 3240 18071 3292 18080
rect 3240 18037 3249 18071
rect 3249 18037 3283 18071
rect 3283 18037 3292 18071
rect 3240 18028 3292 18037
rect 5356 18071 5408 18080
rect 5356 18037 5365 18071
rect 5365 18037 5399 18071
rect 5399 18037 5408 18071
rect 5356 18028 5408 18037
rect 32588 18096 32640 18148
rect 37832 18232 37884 18284
rect 6552 18028 6604 18080
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 7748 18071 7800 18080
rect 7748 18037 7757 18071
rect 7757 18037 7791 18071
rect 7791 18037 7800 18071
rect 7748 18028 7800 18037
rect 12348 18071 12400 18080
rect 12348 18037 12357 18071
rect 12357 18037 12391 18071
rect 12391 18037 12400 18071
rect 12348 18028 12400 18037
rect 12440 18028 12492 18080
rect 13176 18028 13228 18080
rect 20076 18071 20128 18080
rect 20076 18037 20085 18071
rect 20085 18037 20119 18071
rect 20119 18037 20128 18071
rect 20076 18028 20128 18037
rect 22284 18071 22336 18080
rect 22284 18037 22293 18071
rect 22293 18037 22327 18071
rect 22327 18037 22336 18071
rect 22284 18028 22336 18037
rect 30564 18028 30616 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1584 17824 1636 17876
rect 2136 17824 2188 17876
rect 3056 17824 3108 17876
rect 5080 17824 5132 17876
rect 7472 17824 7524 17876
rect 8392 17867 8444 17876
rect 8392 17833 8401 17867
rect 8401 17833 8435 17867
rect 8435 17833 8444 17867
rect 8392 17824 8444 17833
rect 9404 17867 9456 17876
rect 9404 17833 9413 17867
rect 9413 17833 9447 17867
rect 9447 17833 9456 17867
rect 9404 17824 9456 17833
rect 9588 17824 9640 17876
rect 12348 17867 12400 17876
rect 12348 17833 12357 17867
rect 12357 17833 12391 17867
rect 12391 17833 12400 17867
rect 12348 17824 12400 17833
rect 3608 17756 3660 17808
rect 4068 17799 4120 17808
rect 4068 17765 4077 17799
rect 4077 17765 4111 17799
rect 4111 17765 4120 17799
rect 4068 17756 4120 17765
rect 2596 17731 2648 17740
rect 2596 17697 2605 17731
rect 2605 17697 2639 17731
rect 2639 17697 2648 17731
rect 2596 17688 2648 17697
rect 3240 17688 3292 17740
rect 5172 17756 5224 17808
rect 9680 17756 9732 17808
rect 5540 17731 5592 17740
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 2504 17663 2556 17672
rect 2504 17629 2513 17663
rect 2513 17629 2547 17663
rect 2547 17629 2556 17663
rect 2504 17620 2556 17629
rect 5540 17697 5549 17731
rect 5549 17697 5583 17731
rect 5583 17697 5592 17731
rect 5540 17688 5592 17697
rect 8392 17688 8444 17740
rect 9588 17663 9640 17672
rect 9588 17629 9597 17663
rect 9597 17629 9631 17663
rect 9631 17629 9640 17663
rect 9588 17620 9640 17629
rect 2596 17484 2648 17536
rect 5080 17552 5132 17604
rect 5448 17552 5500 17604
rect 9312 17595 9364 17604
rect 9312 17561 9321 17595
rect 9321 17561 9355 17595
rect 9355 17561 9364 17595
rect 9312 17552 9364 17561
rect 12532 17756 12584 17808
rect 15200 17824 15252 17876
rect 16304 17824 16356 17876
rect 16856 17824 16908 17876
rect 18604 17824 18656 17876
rect 20260 17824 20312 17876
rect 29920 17824 29972 17876
rect 30840 17824 30892 17876
rect 32588 17867 32640 17876
rect 32588 17833 32597 17867
rect 32597 17833 32631 17867
rect 32631 17833 32640 17867
rect 32588 17824 32640 17833
rect 38016 17867 38068 17876
rect 38016 17833 38025 17867
rect 38025 17833 38059 17867
rect 38059 17833 38068 17867
rect 38016 17824 38068 17833
rect 18144 17756 18196 17808
rect 18788 17756 18840 17808
rect 27160 17756 27212 17808
rect 12624 17688 12676 17740
rect 12716 17688 12768 17740
rect 12348 17620 12400 17672
rect 12532 17663 12584 17672
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 18512 17688 18564 17740
rect 20076 17731 20128 17740
rect 20076 17697 20085 17731
rect 20085 17697 20119 17731
rect 20119 17697 20128 17731
rect 20076 17688 20128 17697
rect 23848 17688 23900 17740
rect 13176 17663 13228 17672
rect 13176 17629 13185 17663
rect 13185 17629 13219 17663
rect 13219 17629 13228 17663
rect 13176 17620 13228 17629
rect 13360 17620 13412 17672
rect 16304 17663 16356 17672
rect 16304 17629 16313 17663
rect 16313 17629 16347 17663
rect 16347 17629 16356 17663
rect 16304 17620 16356 17629
rect 30564 17663 30616 17672
rect 4988 17484 5040 17536
rect 9864 17484 9916 17536
rect 12900 17552 12952 17604
rect 19248 17595 19300 17604
rect 12808 17484 12860 17536
rect 13544 17484 13596 17536
rect 17776 17484 17828 17536
rect 19248 17561 19257 17595
rect 19257 17561 19291 17595
rect 19291 17561 19300 17595
rect 19248 17552 19300 17561
rect 30564 17629 30573 17663
rect 30573 17629 30607 17663
rect 30607 17629 30616 17663
rect 30564 17620 30616 17629
rect 31208 17663 31260 17672
rect 31208 17629 31217 17663
rect 31217 17629 31251 17663
rect 31251 17629 31260 17663
rect 31208 17620 31260 17629
rect 35624 17620 35676 17672
rect 37740 17620 37792 17672
rect 20260 17595 20312 17604
rect 20260 17561 20269 17595
rect 20269 17561 20303 17595
rect 20303 17561 20312 17595
rect 20260 17552 20312 17561
rect 31484 17595 31536 17604
rect 31484 17561 31518 17595
rect 31518 17561 31536 17595
rect 31484 17552 31536 17561
rect 22744 17484 22796 17536
rect 30564 17484 30616 17536
rect 31392 17484 31444 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 5448 17323 5500 17332
rect 1400 17255 1452 17264
rect 1400 17221 1409 17255
rect 1409 17221 1443 17255
rect 1443 17221 1452 17255
rect 1400 17212 1452 17221
rect 2964 17255 3016 17264
rect 2964 17221 2973 17255
rect 2973 17221 3007 17255
rect 3007 17221 3016 17255
rect 2964 17212 3016 17221
rect 5448 17289 5457 17323
rect 5457 17289 5491 17323
rect 5491 17289 5500 17323
rect 5448 17280 5500 17289
rect 9312 17280 9364 17332
rect 10140 17280 10192 17332
rect 18788 17323 18840 17332
rect 18788 17289 18797 17323
rect 18797 17289 18831 17323
rect 18831 17289 18840 17323
rect 18788 17280 18840 17289
rect 20720 17280 20772 17332
rect 29552 17323 29604 17332
rect 13544 17255 13596 17264
rect 13544 17221 13553 17255
rect 13553 17221 13587 17255
rect 13587 17221 13596 17255
rect 13544 17212 13596 17221
rect 18144 17255 18196 17264
rect 18144 17221 18153 17255
rect 18153 17221 18187 17255
rect 18187 17221 18196 17255
rect 18144 17212 18196 17221
rect 23112 17212 23164 17264
rect 23388 17255 23440 17264
rect 23388 17221 23397 17255
rect 23397 17221 23431 17255
rect 23431 17221 23440 17255
rect 23388 17212 23440 17221
rect 2504 17144 2556 17196
rect 2688 17144 2740 17196
rect 3148 17144 3200 17196
rect 5632 17187 5684 17196
rect 2320 17076 2372 17128
rect 3056 17119 3108 17128
rect 3056 17085 3065 17119
rect 3065 17085 3099 17119
rect 3099 17085 3108 17119
rect 3056 17076 3108 17085
rect 3976 17076 4028 17128
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 9680 17144 9732 17196
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 12900 17144 12952 17196
rect 13360 17187 13412 17196
rect 13360 17153 13369 17187
rect 13369 17153 13403 17187
rect 13403 17153 13412 17187
rect 13360 17144 13412 17153
rect 22744 17187 22796 17196
rect 22744 17153 22753 17187
rect 22753 17153 22787 17187
rect 22787 17153 22796 17187
rect 22744 17144 22796 17153
rect 23204 17144 23256 17196
rect 5540 17076 5592 17128
rect 12624 17119 12676 17128
rect 12624 17085 12633 17119
rect 12633 17085 12667 17119
rect 12667 17085 12676 17119
rect 12624 17076 12676 17085
rect 15108 17119 15160 17128
rect 15108 17085 15117 17119
rect 15117 17085 15151 17119
rect 15151 17085 15160 17119
rect 15108 17076 15160 17085
rect 18236 17076 18288 17128
rect 18512 17119 18564 17128
rect 18512 17085 18521 17119
rect 18521 17085 18555 17119
rect 18555 17085 18564 17119
rect 18512 17076 18564 17085
rect 23480 17119 23532 17128
rect 23480 17085 23489 17119
rect 23489 17085 23523 17119
rect 23523 17085 23532 17119
rect 23480 17076 23532 17085
rect 24308 17076 24360 17128
rect 29552 17289 29561 17323
rect 29561 17289 29595 17323
rect 29595 17289 29604 17323
rect 29552 17280 29604 17289
rect 30564 17280 30616 17332
rect 31484 17280 31536 17332
rect 35624 17323 35676 17332
rect 35624 17289 35633 17323
rect 35633 17289 35667 17323
rect 35667 17289 35676 17323
rect 35624 17280 35676 17289
rect 29000 17212 29052 17264
rect 32588 17212 32640 17264
rect 27252 17187 27304 17196
rect 27252 17153 27261 17187
rect 27261 17153 27295 17187
rect 27295 17153 27304 17187
rect 27252 17144 27304 17153
rect 30196 17144 30248 17196
rect 30656 17144 30708 17196
rect 22284 17008 22336 17060
rect 2136 16983 2188 16992
rect 2136 16949 2145 16983
rect 2145 16949 2179 16983
rect 2179 16949 2188 16983
rect 2136 16940 2188 16949
rect 2412 16940 2464 16992
rect 2872 16940 2924 16992
rect 4068 16983 4120 16992
rect 4068 16949 4077 16983
rect 4077 16949 4111 16983
rect 4111 16949 4120 16983
rect 4068 16940 4120 16949
rect 8392 16940 8444 16992
rect 9128 16983 9180 16992
rect 9128 16949 9137 16983
rect 9137 16949 9171 16983
rect 9171 16949 9180 16983
rect 9128 16940 9180 16949
rect 12716 16983 12768 16992
rect 12716 16949 12725 16983
rect 12725 16949 12759 16983
rect 12759 16949 12768 16983
rect 12716 16940 12768 16949
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 18328 16983 18380 16992
rect 18328 16949 18352 16983
rect 18352 16949 18380 16983
rect 18328 16940 18380 16949
rect 18420 16983 18472 16992
rect 18420 16949 18429 16983
rect 18429 16949 18463 16983
rect 18463 16949 18472 16983
rect 27160 17008 27212 17060
rect 29736 17008 29788 17060
rect 18420 16940 18472 16949
rect 22928 16983 22980 16992
rect 22928 16949 22937 16983
rect 22937 16949 22971 16983
rect 22971 16949 22980 16983
rect 22928 16940 22980 16949
rect 23388 16983 23440 16992
rect 23388 16949 23397 16983
rect 23397 16949 23431 16983
rect 23431 16949 23440 16983
rect 23388 16940 23440 16949
rect 23848 16983 23900 16992
rect 23848 16949 23857 16983
rect 23857 16949 23891 16983
rect 23891 16949 23900 16983
rect 23848 16940 23900 16949
rect 26884 16940 26936 16992
rect 30288 16940 30340 16992
rect 31024 17076 31076 17128
rect 32680 16940 32732 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2964 16779 3016 16788
rect 2964 16745 2973 16779
rect 2973 16745 3007 16779
rect 3007 16745 3016 16779
rect 2964 16736 3016 16745
rect 3976 16779 4028 16788
rect 3976 16745 4000 16779
rect 4000 16745 4028 16779
rect 3976 16736 4028 16745
rect 4068 16779 4120 16788
rect 4068 16745 4077 16779
rect 4077 16745 4111 16779
rect 4111 16745 4120 16779
rect 12716 16779 12768 16788
rect 4068 16736 4120 16745
rect 12716 16745 12725 16779
rect 12725 16745 12759 16779
rect 12759 16745 12768 16779
rect 12716 16736 12768 16745
rect 18604 16736 18656 16788
rect 23388 16779 23440 16788
rect 23388 16745 23397 16779
rect 23397 16745 23431 16779
rect 23431 16745 23440 16779
rect 23388 16736 23440 16745
rect 8392 16668 8444 16720
rect 15936 16668 15988 16720
rect 18420 16668 18472 16720
rect 4620 16600 4672 16652
rect 9128 16643 9180 16652
rect 9128 16609 9137 16643
rect 9137 16609 9171 16643
rect 9171 16609 9180 16643
rect 9128 16600 9180 16609
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 2504 16532 2556 16584
rect 2872 16532 2924 16584
rect 7748 16575 7800 16584
rect 7748 16541 7757 16575
rect 7757 16541 7791 16575
rect 7791 16541 7800 16575
rect 7748 16532 7800 16541
rect 12624 16600 12676 16652
rect 18328 16643 18380 16652
rect 18328 16609 18337 16643
rect 18337 16609 18371 16643
rect 18371 16609 18380 16643
rect 18328 16600 18380 16609
rect 18972 16600 19024 16652
rect 19984 16600 20036 16652
rect 20260 16600 20312 16652
rect 23480 16600 23532 16652
rect 27620 16736 27672 16788
rect 31208 16736 31260 16788
rect 34704 16736 34756 16788
rect 35532 16736 35584 16788
rect 30656 16668 30708 16720
rect 35624 16600 35676 16652
rect 2412 16464 2464 16516
rect 8208 16464 8260 16516
rect 9404 16464 9456 16516
rect 12440 16464 12492 16516
rect 12992 16532 13044 16584
rect 18144 16575 18196 16584
rect 18144 16541 18153 16575
rect 18153 16541 18187 16575
rect 18187 16541 18196 16575
rect 18144 16532 18196 16541
rect 18512 16532 18564 16584
rect 23112 16575 23164 16584
rect 23112 16541 23121 16575
rect 23121 16541 23155 16575
rect 23155 16541 23164 16575
rect 23112 16532 23164 16541
rect 23204 16532 23256 16584
rect 26884 16575 26936 16584
rect 26884 16541 26918 16575
rect 26918 16541 26936 16575
rect 26884 16532 26936 16541
rect 15108 16464 15160 16516
rect 7564 16439 7616 16448
rect 7564 16405 7573 16439
rect 7573 16405 7607 16439
rect 7607 16405 7616 16439
rect 7564 16396 7616 16405
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 16212 16396 16264 16448
rect 18604 16439 18656 16448
rect 18604 16405 18613 16439
rect 18613 16405 18647 16439
rect 18647 16405 18656 16439
rect 18604 16396 18656 16405
rect 24860 16396 24912 16448
rect 27712 16396 27764 16448
rect 29092 16396 29144 16448
rect 30288 16575 30340 16584
rect 30288 16541 30297 16575
rect 30297 16541 30331 16575
rect 30331 16541 30340 16575
rect 30288 16532 30340 16541
rect 36268 16464 36320 16516
rect 37188 16439 37240 16448
rect 37188 16405 37197 16439
rect 37197 16405 37231 16439
rect 37231 16405 37240 16439
rect 37188 16396 37240 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 9404 16235 9456 16244
rect 9404 16201 9413 16235
rect 9413 16201 9447 16235
rect 9447 16201 9456 16235
rect 9404 16192 9456 16201
rect 27252 16192 27304 16244
rect 27712 16192 27764 16244
rect 36268 16235 36320 16244
rect 36268 16201 36277 16235
rect 36277 16201 36311 16235
rect 36311 16201 36320 16235
rect 36268 16192 36320 16201
rect 27804 16124 27856 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 3148 16099 3200 16108
rect 3148 16065 3157 16099
rect 3157 16065 3191 16099
rect 3191 16065 3200 16099
rect 3148 16056 3200 16065
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 9588 16099 9640 16108
rect 9588 16065 9597 16099
rect 9597 16065 9631 16099
rect 9631 16065 9640 16099
rect 9588 16056 9640 16065
rect 12900 16099 12952 16108
rect 12900 16065 12909 16099
rect 12909 16065 12943 16099
rect 12943 16065 12952 16099
rect 12900 16056 12952 16065
rect 15936 16056 15988 16108
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 17868 16056 17920 16108
rect 24860 16099 24912 16108
rect 24860 16065 24869 16099
rect 24869 16065 24903 16099
rect 24903 16065 24912 16099
rect 24860 16056 24912 16065
rect 18328 15988 18380 16040
rect 22560 16031 22612 16040
rect 22560 15997 22569 16031
rect 22569 15997 22603 16031
rect 22603 15997 22612 16031
rect 22560 15988 22612 15997
rect 23204 15988 23256 16040
rect 23480 16031 23532 16040
rect 23480 15997 23489 16031
rect 23489 15997 23523 16031
rect 23523 15997 23532 16031
rect 23480 15988 23532 15997
rect 4620 15920 4672 15972
rect 17960 15963 18012 15972
rect 17960 15929 17969 15963
rect 17969 15929 18003 15963
rect 18003 15929 18012 15963
rect 17960 15920 18012 15929
rect 2504 15852 2556 15904
rect 6368 15895 6420 15904
rect 6368 15861 6377 15895
rect 6377 15861 6411 15895
rect 6411 15861 6420 15895
rect 6368 15852 6420 15861
rect 12716 15895 12768 15904
rect 12716 15861 12725 15895
rect 12725 15861 12759 15895
rect 12759 15861 12768 15895
rect 12716 15852 12768 15861
rect 13268 15852 13320 15904
rect 13820 15852 13872 15904
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 17408 15852 17460 15904
rect 20812 15895 20864 15904
rect 20812 15861 20821 15895
rect 20821 15861 20855 15895
rect 20855 15861 20864 15895
rect 20812 15852 20864 15861
rect 26056 15852 26108 15904
rect 32496 16056 32548 16108
rect 30196 15988 30248 16040
rect 35532 16056 35584 16108
rect 36084 16124 36136 16176
rect 36452 16124 36504 16176
rect 37188 16056 37240 16108
rect 29092 15852 29144 15904
rect 35348 15852 35400 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 13084 15512 13136 15564
rect 4160 15444 4212 15496
rect 6184 15487 6236 15496
rect 6184 15453 6193 15487
rect 6193 15453 6227 15487
rect 6227 15453 6236 15487
rect 6184 15444 6236 15453
rect 7380 15444 7432 15496
rect 8668 15444 8720 15496
rect 12532 15444 12584 15496
rect 4620 15376 4672 15428
rect 16212 15623 16264 15632
rect 16212 15589 16221 15623
rect 16221 15589 16255 15623
rect 16255 15589 16264 15623
rect 16212 15580 16264 15589
rect 16948 15648 17000 15700
rect 18052 15648 18104 15700
rect 18328 15648 18380 15700
rect 23204 15691 23256 15700
rect 23204 15657 23213 15691
rect 23213 15657 23247 15691
rect 23247 15657 23256 15691
rect 23204 15648 23256 15657
rect 32680 15691 32732 15700
rect 32680 15657 32689 15691
rect 32689 15657 32723 15691
rect 32723 15657 32732 15691
rect 32680 15648 32732 15657
rect 35900 15648 35952 15700
rect 36084 15691 36136 15700
rect 36084 15657 36093 15691
rect 36093 15657 36127 15691
rect 36127 15657 36136 15691
rect 36084 15648 36136 15657
rect 24676 15580 24728 15632
rect 17960 15512 18012 15564
rect 20812 15555 20864 15564
rect 20812 15521 20821 15555
rect 20821 15521 20855 15555
rect 20855 15521 20864 15555
rect 20812 15512 20864 15521
rect 22192 15555 22244 15564
rect 22192 15521 22201 15555
rect 22201 15521 22235 15555
rect 22235 15521 22244 15555
rect 22192 15512 22244 15521
rect 23848 15512 23900 15564
rect 35808 15555 35860 15564
rect 35808 15521 35817 15555
rect 35817 15521 35851 15555
rect 35851 15521 35860 15555
rect 35808 15512 35860 15521
rect 13268 15487 13320 15496
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 13268 15444 13320 15453
rect 15936 15487 15988 15496
rect 13360 15376 13412 15428
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 19432 15444 19484 15496
rect 22928 15444 22980 15496
rect 25412 15487 25464 15496
rect 25412 15453 25421 15487
rect 25421 15453 25455 15487
rect 25455 15453 25464 15487
rect 25412 15444 25464 15453
rect 29736 15444 29788 15496
rect 32220 15444 32272 15496
rect 35440 15444 35492 15496
rect 20720 15376 20772 15428
rect 20996 15419 21048 15428
rect 20996 15385 21005 15419
rect 21005 15385 21039 15419
rect 21039 15385 21048 15419
rect 20996 15376 21048 15385
rect 30196 15419 30248 15428
rect 30196 15385 30205 15419
rect 30205 15385 30239 15419
rect 30239 15385 30248 15419
rect 30196 15376 30248 15385
rect 15292 15308 15344 15360
rect 16212 15308 16264 15360
rect 16856 15308 16908 15360
rect 17868 15351 17920 15360
rect 17868 15317 17877 15351
rect 17877 15317 17911 15351
rect 17911 15317 17920 15351
rect 17868 15308 17920 15317
rect 27804 15351 27856 15360
rect 27804 15317 27813 15351
rect 27813 15317 27847 15351
rect 27847 15317 27856 15351
rect 27804 15308 27856 15317
rect 29092 15308 29144 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 9588 15104 9640 15156
rect 19984 15104 20036 15156
rect 20996 15104 21048 15156
rect 25412 15104 25464 15156
rect 29736 15147 29788 15156
rect 4160 15079 4212 15088
rect 4160 15045 4169 15079
rect 4169 15045 4203 15079
rect 4203 15045 4212 15079
rect 4160 15036 4212 15045
rect 7564 15079 7616 15088
rect 7564 15045 7573 15079
rect 7573 15045 7607 15079
rect 7607 15045 7616 15079
rect 7564 15036 7616 15045
rect 10140 15079 10192 15088
rect 10140 15045 10149 15079
rect 10149 15045 10183 15079
rect 10183 15045 10192 15079
rect 10140 15036 10192 15045
rect 12716 15079 12768 15088
rect 12716 15045 12725 15079
rect 12725 15045 12759 15079
rect 12759 15045 12768 15079
rect 12716 15036 12768 15045
rect 24400 15079 24452 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 9496 14968 9548 15020
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 3240 14900 3292 14952
rect 10048 14943 10100 14952
rect 4068 14832 4120 14884
rect 10048 14909 10057 14943
rect 10057 14909 10091 14943
rect 10091 14909 10100 14943
rect 10048 14900 10100 14909
rect 12992 14943 13044 14952
rect 12992 14909 13001 14943
rect 13001 14909 13035 14943
rect 13035 14909 13044 14943
rect 12992 14900 13044 14909
rect 16948 14943 17000 14952
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 2780 14764 2832 14816
rect 3884 14764 3936 14816
rect 9772 14832 9824 14884
rect 19616 14968 19668 15020
rect 19800 14968 19852 15020
rect 19432 14943 19484 14952
rect 19432 14909 19441 14943
rect 19441 14909 19475 14943
rect 19475 14909 19484 14943
rect 19432 14900 19484 14909
rect 24400 15045 24409 15079
rect 24409 15045 24443 15079
rect 24443 15045 24452 15079
rect 24400 15036 24452 15045
rect 26056 15079 26108 15088
rect 26056 15045 26065 15079
rect 26065 15045 26099 15079
rect 26099 15045 26108 15079
rect 26056 15036 26108 15045
rect 29736 15113 29745 15147
rect 29745 15113 29779 15147
rect 29779 15113 29788 15147
rect 29736 15104 29788 15113
rect 29276 15036 29328 15088
rect 35900 15036 35952 15088
rect 36452 15036 36504 15088
rect 22560 14968 22612 15020
rect 34796 14968 34848 15020
rect 35532 15011 35584 15020
rect 35532 14977 35541 15011
rect 35541 14977 35575 15011
rect 35575 14977 35584 15011
rect 35532 14968 35584 14977
rect 22192 14900 22244 14952
rect 19524 14832 19576 14884
rect 20536 14832 20588 14884
rect 27896 14900 27948 14952
rect 30380 14832 30432 14884
rect 35348 14832 35400 14884
rect 9312 14764 9364 14816
rect 19340 14807 19392 14816
rect 19340 14773 19349 14807
rect 19349 14773 19383 14807
rect 19383 14773 19392 14807
rect 19340 14764 19392 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3240 14603 3292 14612
rect 3240 14569 3249 14603
rect 3249 14569 3283 14603
rect 3283 14569 3292 14603
rect 3240 14560 3292 14569
rect 9312 14560 9364 14612
rect 19340 14603 19392 14612
rect 19340 14569 19349 14603
rect 19349 14569 19383 14603
rect 19383 14569 19392 14603
rect 19340 14560 19392 14569
rect 19800 14603 19852 14612
rect 19800 14569 19809 14603
rect 19809 14569 19843 14603
rect 19843 14569 19852 14603
rect 19800 14560 19852 14569
rect 34336 14560 34388 14612
rect 3976 14492 4028 14544
rect 5356 14467 5408 14476
rect 5356 14433 5365 14467
rect 5365 14433 5399 14467
rect 5399 14433 5408 14467
rect 5356 14424 5408 14433
rect 6184 14424 6236 14476
rect 18604 14492 18656 14544
rect 9128 14424 9180 14476
rect 10048 14424 10100 14476
rect 10600 14424 10652 14476
rect 19432 14467 19484 14476
rect 19432 14433 19441 14467
rect 19441 14433 19475 14467
rect 19475 14433 19484 14467
rect 19432 14424 19484 14433
rect 5172 14356 5224 14408
rect 9496 14356 9548 14408
rect 23664 14424 23716 14476
rect 27160 14467 27212 14476
rect 27160 14433 27169 14467
rect 27169 14433 27203 14467
rect 27203 14433 27212 14467
rect 27160 14424 27212 14433
rect 30196 14424 30248 14476
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 19984 14356 20036 14408
rect 5356 14288 5408 14340
rect 6368 14288 6420 14340
rect 10232 14288 10284 14340
rect 17316 14288 17368 14340
rect 19248 14288 19300 14340
rect 19524 14288 19576 14340
rect 21824 14331 21876 14340
rect 21824 14297 21833 14331
rect 21833 14297 21867 14331
rect 21867 14297 21876 14331
rect 21824 14288 21876 14297
rect 29276 14356 29328 14408
rect 29552 14288 29604 14340
rect 31852 14356 31904 14408
rect 32220 14356 32272 14408
rect 35532 14560 35584 14612
rect 36452 14424 36504 14476
rect 30380 14288 30432 14340
rect 34980 14399 35032 14408
rect 34980 14365 34989 14399
rect 34989 14365 35023 14399
rect 35023 14365 35032 14399
rect 34980 14356 35032 14365
rect 38016 14331 38068 14340
rect 38016 14297 38025 14331
rect 38025 14297 38059 14331
rect 38059 14297 38068 14331
rect 38016 14288 38068 14297
rect 9220 14263 9272 14272
rect 9220 14229 9229 14263
rect 9229 14229 9263 14263
rect 9263 14229 9272 14263
rect 9220 14220 9272 14229
rect 10140 14263 10192 14272
rect 10140 14229 10149 14263
rect 10149 14229 10183 14263
rect 10183 14229 10192 14263
rect 10140 14220 10192 14229
rect 26148 14263 26200 14272
rect 26148 14229 26157 14263
rect 26157 14229 26191 14263
rect 26191 14229 26200 14263
rect 26148 14220 26200 14229
rect 26608 14263 26660 14272
rect 26608 14229 26617 14263
rect 26617 14229 26651 14263
rect 26651 14229 26660 14263
rect 26608 14220 26660 14229
rect 27896 14220 27948 14272
rect 29184 14220 29236 14272
rect 33140 14263 33192 14272
rect 33140 14229 33149 14263
rect 33149 14229 33183 14263
rect 33183 14229 33192 14263
rect 33140 14220 33192 14229
rect 34428 14220 34480 14272
rect 34704 14263 34756 14272
rect 34704 14229 34713 14263
rect 34713 14229 34747 14263
rect 34747 14229 34756 14263
rect 34704 14220 34756 14229
rect 37924 14263 37976 14272
rect 37924 14229 37933 14263
rect 37933 14229 37967 14263
rect 37967 14229 37976 14263
rect 37924 14220 37976 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 16120 14016 16172 14068
rect 16948 14016 17000 14068
rect 17316 14059 17368 14068
rect 17316 14025 17325 14059
rect 17325 14025 17359 14059
rect 17359 14025 17368 14059
rect 17316 14016 17368 14025
rect 19248 14059 19300 14068
rect 19248 14025 19257 14059
rect 19257 14025 19291 14059
rect 19291 14025 19300 14059
rect 19248 14016 19300 14025
rect 21824 14016 21876 14068
rect 27160 14016 27212 14068
rect 30380 14016 30432 14068
rect 32220 14059 32272 14068
rect 32220 14025 32229 14059
rect 32229 14025 32263 14059
rect 32263 14025 32272 14059
rect 32220 14016 32272 14025
rect 34980 14016 35032 14068
rect 35808 14016 35860 14068
rect 5172 13991 5224 14000
rect 5172 13957 5181 13991
rect 5181 13957 5215 13991
rect 5215 13957 5224 13991
rect 5172 13948 5224 13957
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 10140 13948 10192 14000
rect 12992 13991 13044 14000
rect 5356 13880 5408 13889
rect 8668 13923 8720 13932
rect 8668 13889 8677 13923
rect 8677 13889 8711 13923
rect 8711 13889 8720 13923
rect 8668 13880 8720 13889
rect 3976 13855 4028 13864
rect 3976 13821 3985 13855
rect 3985 13821 4019 13855
rect 4019 13821 4028 13855
rect 3976 13812 4028 13821
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 8852 13855 8904 13864
rect 8852 13821 8861 13855
rect 8861 13821 8895 13855
rect 8895 13821 8904 13855
rect 8852 13812 8904 13821
rect 9128 13855 9180 13864
rect 9128 13821 9137 13855
rect 9137 13821 9171 13855
rect 9171 13821 9180 13855
rect 12992 13957 13001 13991
rect 13001 13957 13035 13991
rect 13035 13957 13044 13991
rect 12992 13948 13044 13957
rect 10600 13880 10652 13932
rect 17224 13880 17276 13932
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 20996 13923 21048 13932
rect 20996 13889 21005 13923
rect 21005 13889 21039 13923
rect 21039 13889 21048 13923
rect 20996 13880 21048 13889
rect 29092 13948 29144 14000
rect 29184 13923 29236 13932
rect 29184 13889 29193 13923
rect 29193 13889 29227 13923
rect 29227 13889 29236 13923
rect 29184 13880 29236 13889
rect 9128 13812 9180 13821
rect 12532 13812 12584 13864
rect 14648 13855 14700 13864
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 14832 13855 14884 13864
rect 14832 13821 14841 13855
rect 14841 13821 14875 13855
rect 14875 13821 14884 13855
rect 14832 13812 14884 13821
rect 27896 13744 27948 13796
rect 33324 13923 33376 13932
rect 33324 13889 33342 13923
rect 33342 13889 33376 13923
rect 33324 13880 33376 13889
rect 30380 13744 30432 13796
rect 31484 13812 31536 13864
rect 33600 13855 33652 13864
rect 33600 13821 33609 13855
rect 33609 13821 33643 13855
rect 33643 13821 33652 13855
rect 33600 13812 33652 13821
rect 30932 13744 30984 13796
rect 34336 13923 34388 13932
rect 34336 13889 34345 13923
rect 34345 13889 34379 13923
rect 34379 13889 34388 13923
rect 34336 13880 34388 13889
rect 35256 13880 35308 13932
rect 35532 13880 35584 13932
rect 37280 13923 37332 13932
rect 37280 13889 37289 13923
rect 37289 13889 37323 13923
rect 37323 13889 37332 13923
rect 37280 13880 37332 13889
rect 34520 13812 34572 13864
rect 29368 13719 29420 13728
rect 29368 13685 29377 13719
rect 29377 13685 29411 13719
rect 29411 13685 29420 13719
rect 29368 13676 29420 13685
rect 37648 13676 37700 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 8852 13472 8904 13524
rect 10048 13515 10100 13524
rect 10048 13481 10057 13515
rect 10057 13481 10091 13515
rect 10091 13481 10100 13515
rect 10048 13472 10100 13481
rect 10232 13472 10284 13524
rect 10508 13472 10560 13524
rect 14832 13472 14884 13524
rect 16764 13515 16816 13524
rect 16764 13481 16773 13515
rect 16773 13481 16807 13515
rect 16807 13481 16816 13515
rect 16764 13472 16816 13481
rect 17224 13515 17276 13524
rect 17224 13481 17233 13515
rect 17233 13481 17267 13515
rect 17267 13481 17276 13515
rect 17224 13472 17276 13481
rect 19340 13472 19392 13524
rect 20996 13472 21048 13524
rect 7012 13404 7064 13456
rect 8208 13404 8260 13456
rect 4160 13336 4212 13388
rect 5540 13336 5592 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 8392 13311 8444 13320
rect 7012 13268 7064 13277
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 10508 13268 10560 13320
rect 17500 13404 17552 13456
rect 16028 13379 16080 13388
rect 16028 13345 16037 13379
rect 16037 13345 16071 13379
rect 16071 13345 16080 13379
rect 16028 13336 16080 13345
rect 19432 13336 19484 13388
rect 20536 13336 20588 13388
rect 27620 13472 27672 13524
rect 30932 13515 30984 13524
rect 30932 13481 30941 13515
rect 30941 13481 30975 13515
rect 30975 13481 30984 13515
rect 30932 13472 30984 13481
rect 33324 13472 33376 13524
rect 36452 13515 36504 13524
rect 36452 13481 36461 13515
rect 36461 13481 36495 13515
rect 36495 13481 36504 13515
rect 36452 13472 36504 13481
rect 27896 13447 27948 13456
rect 27896 13413 27905 13447
rect 27905 13413 27939 13447
rect 27939 13413 27948 13447
rect 27896 13404 27948 13413
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 15200 13268 15252 13320
rect 18236 13268 18288 13320
rect 19984 13311 20036 13320
rect 19984 13277 19993 13311
rect 19993 13277 20027 13311
rect 20027 13277 20036 13311
rect 19984 13268 20036 13277
rect 22284 13268 22336 13320
rect 26608 13268 26660 13320
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 12900 13200 12952 13252
rect 20444 13200 20496 13252
rect 25872 13243 25924 13252
rect 25872 13209 25881 13243
rect 25881 13209 25915 13243
rect 25915 13209 25924 13243
rect 25872 13200 25924 13209
rect 26976 13200 27028 13252
rect 33140 13311 33192 13320
rect 33140 13277 33149 13311
rect 33149 13277 33183 13311
rect 33183 13277 33192 13311
rect 33140 13268 33192 13277
rect 33600 13268 33652 13320
rect 29828 13243 29880 13252
rect 29828 13209 29862 13243
rect 29862 13209 29880 13243
rect 29828 13200 29880 13209
rect 31668 13200 31720 13252
rect 34520 13200 34572 13252
rect 34796 13200 34848 13252
rect 35440 13200 35492 13252
rect 16856 13132 16908 13184
rect 27160 13132 27212 13184
rect 29000 13175 29052 13184
rect 29000 13141 29009 13175
rect 29009 13141 29043 13175
rect 29043 13141 29052 13175
rect 29000 13132 29052 13141
rect 34428 13132 34480 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 10508 12928 10560 12980
rect 11428 12928 11480 12980
rect 2504 12903 2556 12912
rect 2504 12869 2513 12903
rect 2513 12869 2547 12903
rect 2547 12869 2556 12903
rect 2504 12860 2556 12869
rect 2780 12835 2832 12844
rect 2780 12801 2789 12835
rect 2789 12801 2823 12835
rect 2823 12801 2832 12835
rect 2780 12792 2832 12801
rect 7012 12792 7064 12844
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 8392 12792 8444 12801
rect 15200 12928 15252 12980
rect 17040 12971 17092 12980
rect 17040 12937 17049 12971
rect 17049 12937 17083 12971
rect 17083 12937 17092 12971
rect 17040 12928 17092 12937
rect 16764 12860 16816 12912
rect 19340 12928 19392 12980
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 14648 12835 14700 12844
rect 14648 12801 14657 12835
rect 14657 12801 14691 12835
rect 14691 12801 14700 12835
rect 14648 12792 14700 12801
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 19432 12792 19484 12844
rect 20168 12928 20220 12980
rect 26976 12971 27028 12980
rect 26976 12937 26985 12971
rect 26985 12937 27019 12971
rect 27019 12937 27028 12971
rect 26976 12928 27028 12937
rect 29828 12971 29880 12980
rect 29828 12937 29837 12971
rect 29837 12937 29871 12971
rect 29871 12937 29880 12971
rect 29828 12928 29880 12937
rect 34704 12928 34756 12980
rect 20352 12792 20404 12844
rect 22284 12835 22336 12844
rect 22284 12801 22293 12835
rect 22293 12801 22327 12835
rect 22327 12801 22336 12835
rect 22284 12792 22336 12801
rect 27160 12835 27212 12844
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 29368 12792 29420 12844
rect 34428 12835 34480 12844
rect 34428 12801 34437 12835
rect 34437 12801 34471 12835
rect 34471 12801 34480 12835
rect 34428 12792 34480 12801
rect 34704 12835 34756 12844
rect 34704 12801 34713 12835
rect 34713 12801 34747 12835
rect 34747 12801 34756 12835
rect 34704 12792 34756 12801
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 8576 12767 8628 12776
rect 8576 12733 8585 12767
rect 8585 12733 8619 12767
rect 8619 12733 8628 12767
rect 8576 12724 8628 12733
rect 9772 12767 9824 12776
rect 9772 12733 9781 12767
rect 9781 12733 9815 12767
rect 9815 12733 9824 12767
rect 9772 12724 9824 12733
rect 17868 12724 17920 12776
rect 18604 12724 18656 12776
rect 22468 12767 22520 12776
rect 22468 12733 22477 12767
rect 22477 12733 22511 12767
rect 22511 12733 22520 12767
rect 22468 12724 22520 12733
rect 23480 12767 23532 12776
rect 23480 12733 23489 12767
rect 23489 12733 23523 12767
rect 23523 12733 23532 12767
rect 23480 12724 23532 12733
rect 20444 12656 20496 12708
rect 34796 12656 34848 12708
rect 1584 12588 1636 12640
rect 2412 12588 2464 12640
rect 3976 12588 4028 12640
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 35440 12588 35492 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2596 12427 2648 12436
rect 2596 12393 2605 12427
rect 2605 12393 2639 12427
rect 2639 12393 2648 12427
rect 2596 12384 2648 12393
rect 10416 12384 10468 12436
rect 2412 12248 2464 12300
rect 4804 12248 4856 12300
rect 5540 12248 5592 12300
rect 8576 12248 8628 12300
rect 10600 12248 10652 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 15108 12384 15160 12436
rect 20352 12384 20404 12436
rect 22468 12384 22520 12436
rect 35440 12427 35492 12436
rect 35440 12393 35449 12427
rect 35449 12393 35483 12427
rect 35483 12393 35492 12427
rect 35440 12384 35492 12393
rect 37280 12384 37332 12436
rect 18236 12291 18288 12300
rect 18236 12257 18245 12291
rect 18245 12257 18279 12291
rect 18279 12257 18288 12291
rect 18236 12248 18288 12257
rect 26148 12248 26200 12300
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 20904 12180 20956 12232
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 35348 12180 35400 12232
rect 6368 12112 6420 12164
rect 10048 12112 10100 12164
rect 14648 12112 14700 12164
rect 21916 12112 21968 12164
rect 22100 12155 22152 12164
rect 22100 12121 22109 12155
rect 22109 12121 22143 12155
rect 22143 12121 22152 12155
rect 22100 12112 22152 12121
rect 25504 12112 25556 12164
rect 25872 12155 25924 12164
rect 25872 12121 25881 12155
rect 25881 12121 25915 12155
rect 25915 12121 25924 12155
rect 25872 12112 25924 12121
rect 30380 12112 30432 12164
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 2964 12044 3016 12096
rect 10692 12044 10744 12096
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 20260 12044 20312 12096
rect 26976 12044 27028 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 6368 11883 6420 11892
rect 6368 11849 6377 11883
rect 6377 11849 6411 11883
rect 6411 11849 6420 11883
rect 6368 11840 6420 11849
rect 11428 11840 11480 11892
rect 17868 11840 17920 11892
rect 1400 11815 1452 11824
rect 1400 11781 1409 11815
rect 1409 11781 1443 11815
rect 1443 11781 1452 11815
rect 1400 11772 1452 11781
rect 10692 11704 10744 11756
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 14004 11772 14056 11824
rect 18512 11772 18564 11824
rect 10784 11704 10836 11713
rect 13360 11704 13412 11756
rect 16856 11704 16908 11756
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 19432 11704 19484 11756
rect 20628 11840 20680 11892
rect 23020 11840 23072 11892
rect 25504 11883 25556 11892
rect 25504 11849 25513 11883
rect 25513 11849 25547 11883
rect 25547 11849 25556 11883
rect 25504 11840 25556 11849
rect 20260 11772 20312 11824
rect 21916 11772 21968 11824
rect 29092 11772 29144 11824
rect 22008 11747 22060 11756
rect 10600 11679 10652 11688
rect 10600 11645 10609 11679
rect 10609 11645 10643 11679
rect 10643 11645 10652 11679
rect 10600 11636 10652 11645
rect 11888 11636 11940 11688
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 16672 11636 16724 11688
rect 17132 11636 17184 11688
rect 22008 11713 22017 11747
rect 22017 11713 22051 11747
rect 22051 11713 22060 11747
rect 22008 11704 22060 11713
rect 15384 11568 15436 11620
rect 10416 11500 10468 11552
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 10968 11543 11020 11552
rect 10968 11509 10977 11543
rect 10977 11509 11011 11543
rect 11011 11509 11020 11543
rect 10968 11500 11020 11509
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 20628 11568 20680 11620
rect 25228 11704 25280 11756
rect 26148 11704 26200 11756
rect 26976 11747 27028 11756
rect 26976 11713 26985 11747
rect 26985 11713 27019 11747
rect 27019 11713 27028 11747
rect 26976 11704 27028 11713
rect 30472 11704 30524 11756
rect 31116 11840 31168 11892
rect 25964 11679 26016 11688
rect 25964 11645 25973 11679
rect 25973 11645 26007 11679
rect 26007 11645 26016 11679
rect 25964 11636 26016 11645
rect 25412 11568 25464 11620
rect 20352 11500 20404 11552
rect 27160 11543 27212 11552
rect 27160 11509 27169 11543
rect 27169 11509 27203 11543
rect 27203 11509 27212 11543
rect 27160 11500 27212 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1584 11296 1636 11348
rect 2596 11296 2648 11348
rect 10600 11296 10652 11348
rect 11888 11339 11940 11348
rect 11888 11305 11897 11339
rect 11897 11305 11931 11339
rect 11931 11305 11940 11339
rect 11888 11296 11940 11305
rect 15384 11339 15436 11348
rect 15384 11305 15393 11339
rect 15393 11305 15427 11339
rect 15427 11305 15436 11339
rect 15384 11296 15436 11305
rect 10876 11228 10928 11280
rect 15108 11228 15160 11280
rect 2504 11160 2556 11212
rect 12532 11160 12584 11212
rect 14004 11160 14056 11212
rect 16672 11296 16724 11348
rect 16856 11339 16908 11348
rect 16856 11305 16865 11339
rect 16865 11305 16899 11339
rect 16899 11305 16908 11339
rect 16856 11296 16908 11305
rect 17592 11296 17644 11348
rect 20352 11339 20404 11348
rect 20352 11305 20361 11339
rect 20361 11305 20395 11339
rect 20395 11305 20404 11339
rect 20352 11296 20404 11305
rect 2228 11092 2280 11144
rect 10508 11092 10560 11144
rect 10784 11092 10836 11144
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 13084 11092 13136 11144
rect 13820 11092 13872 11144
rect 2688 11024 2740 11076
rect 4068 11024 4120 11076
rect 8024 11024 8076 11076
rect 12164 11067 12216 11076
rect 12164 11033 12173 11067
rect 12173 11033 12207 11067
rect 12207 11033 12216 11067
rect 12164 11024 12216 11033
rect 15936 11228 15988 11280
rect 21640 11228 21692 11280
rect 17592 11092 17644 11144
rect 18604 11024 18656 11076
rect 20628 11135 20680 11144
rect 20628 11101 20637 11135
rect 20637 11101 20671 11135
rect 20671 11101 20680 11135
rect 20628 11092 20680 11101
rect 20260 11024 20312 11076
rect 22008 11160 22060 11212
rect 25964 11296 26016 11348
rect 30288 11296 30340 11348
rect 33876 11296 33928 11348
rect 34704 11296 34756 11348
rect 30104 11228 30156 11280
rect 25228 11160 25280 11212
rect 29000 11092 29052 11144
rect 21640 11024 21692 11076
rect 22192 11067 22244 11076
rect 22192 11033 22201 11067
rect 22201 11033 22235 11067
rect 22235 11033 22244 11067
rect 22192 11024 22244 11033
rect 3056 10956 3108 11008
rect 11704 10999 11756 11008
rect 11704 10965 11713 10999
rect 11713 10965 11747 10999
rect 11747 10965 11756 10999
rect 11704 10956 11756 10965
rect 13176 10956 13228 11008
rect 15200 10956 15252 11008
rect 19432 10999 19484 11008
rect 19432 10965 19441 10999
rect 19441 10965 19475 10999
rect 19475 10965 19484 10999
rect 19432 10956 19484 10965
rect 20812 10999 20864 11008
rect 20812 10965 20821 10999
rect 20821 10965 20855 10999
rect 20855 10965 20864 10999
rect 20812 10956 20864 10965
rect 22652 10999 22704 11008
rect 22652 10965 22661 10999
rect 22661 10965 22695 10999
rect 22695 10965 22704 10999
rect 22652 10956 22704 10965
rect 27160 11024 27212 11076
rect 30380 11092 30432 11144
rect 29920 10956 29972 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 15292 10752 15344 10804
rect 10692 10684 10744 10736
rect 12164 10684 12216 10736
rect 12900 10684 12952 10736
rect 15016 10684 15068 10736
rect 16028 10752 16080 10804
rect 22192 10752 22244 10804
rect 30380 10795 30432 10804
rect 30380 10761 30389 10795
rect 30389 10761 30423 10795
rect 30423 10761 30432 10795
rect 30380 10752 30432 10761
rect 31668 10752 31720 10804
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 2872 10659 2924 10668
rect 2872 10625 2881 10659
rect 2881 10625 2915 10659
rect 2915 10625 2924 10659
rect 2872 10616 2924 10625
rect 2964 10616 3016 10668
rect 3332 10616 3384 10668
rect 4620 10616 4672 10668
rect 10508 10659 10560 10668
rect 10508 10625 10517 10659
rect 10517 10625 10551 10659
rect 10551 10625 10560 10659
rect 10508 10616 10560 10625
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 15200 10659 15252 10668
rect 15200 10625 15209 10659
rect 15209 10625 15243 10659
rect 15243 10625 15252 10659
rect 18052 10684 18104 10736
rect 18604 10684 18656 10736
rect 15200 10616 15252 10625
rect 17592 10659 17644 10668
rect 17592 10625 17601 10659
rect 17601 10625 17635 10659
rect 17635 10625 17644 10659
rect 17592 10616 17644 10625
rect 17868 10659 17920 10668
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 18420 10659 18472 10668
rect 18420 10625 18429 10659
rect 18429 10625 18463 10659
rect 18463 10625 18472 10659
rect 18420 10616 18472 10625
rect 30104 10684 30156 10736
rect 20812 10616 20864 10668
rect 30932 10659 30984 10668
rect 30932 10625 30941 10659
rect 30941 10625 30975 10659
rect 30975 10625 30984 10659
rect 30932 10616 30984 10625
rect 34704 10659 34756 10668
rect 34704 10625 34713 10659
rect 34713 10625 34747 10659
rect 34747 10625 34756 10659
rect 34704 10616 34756 10625
rect 34796 10616 34848 10668
rect 1952 10548 2004 10600
rect 3976 10548 4028 10600
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 2504 10480 2556 10532
rect 4712 10480 4764 10532
rect 12532 10548 12584 10600
rect 13820 10548 13872 10600
rect 18512 10548 18564 10600
rect 17224 10523 17276 10532
rect 3056 10455 3108 10464
rect 3056 10421 3080 10455
rect 3080 10421 3108 10455
rect 3056 10412 3108 10421
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 12072 10455 12124 10464
rect 12072 10421 12081 10455
rect 12081 10421 12115 10455
rect 12115 10421 12124 10455
rect 12072 10412 12124 10421
rect 12716 10412 12768 10464
rect 17224 10489 17233 10523
rect 17233 10489 17267 10523
rect 17267 10489 17276 10523
rect 17224 10480 17276 10489
rect 34336 10480 34388 10532
rect 15108 10455 15160 10464
rect 15108 10421 15117 10455
rect 15117 10421 15151 10455
rect 15151 10421 15160 10455
rect 15108 10412 15160 10421
rect 15476 10412 15528 10464
rect 19708 10455 19760 10464
rect 19708 10421 19717 10455
rect 19717 10421 19751 10455
rect 19751 10421 19760 10455
rect 19708 10412 19760 10421
rect 20352 10455 20404 10464
rect 20352 10421 20361 10455
rect 20361 10421 20395 10455
rect 20395 10421 20404 10455
rect 20352 10412 20404 10421
rect 26056 10412 26108 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 2228 10208 2280 10260
rect 4068 10208 4120 10260
rect 4712 10208 4764 10260
rect 11888 10208 11940 10260
rect 15108 10251 15160 10260
rect 15108 10217 15117 10251
rect 15117 10217 15151 10251
rect 15151 10217 15160 10251
rect 15108 10208 15160 10217
rect 16028 10251 16080 10260
rect 16028 10217 16037 10251
rect 16037 10217 16071 10251
rect 16071 10217 16080 10251
rect 16028 10208 16080 10217
rect 20352 10208 20404 10260
rect 2596 10115 2648 10124
rect 2596 10081 2605 10115
rect 2605 10081 2639 10115
rect 2639 10081 2648 10115
rect 2596 10072 2648 10081
rect 11060 10115 11112 10124
rect 11060 10081 11069 10115
rect 11069 10081 11103 10115
rect 11103 10081 11112 10115
rect 11060 10072 11112 10081
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 2780 10004 2832 10013
rect 3884 10004 3936 10056
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 2596 9936 2648 9988
rect 5540 9979 5592 9988
rect 5540 9945 5574 9979
rect 5574 9945 5592 9979
rect 10324 9979 10376 9988
rect 5540 9936 5592 9945
rect 10324 9945 10333 9979
rect 10333 9945 10367 9979
rect 10367 9945 10376 9979
rect 10324 9936 10376 9945
rect 19432 10072 19484 10124
rect 24400 10115 24452 10124
rect 24400 10081 24409 10115
rect 24409 10081 24443 10115
rect 24443 10081 24452 10115
rect 24400 10072 24452 10081
rect 26056 10115 26108 10124
rect 26056 10081 26065 10115
rect 26065 10081 26099 10115
rect 26099 10081 26108 10115
rect 26056 10072 26108 10081
rect 30288 10072 30340 10124
rect 13820 10004 13872 10056
rect 15016 10047 15068 10056
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 20812 10004 20864 10056
rect 30840 10047 30892 10056
rect 30840 10013 30849 10047
rect 30849 10013 30883 10047
rect 30883 10013 30892 10047
rect 30840 10004 30892 10013
rect 31300 10072 31352 10124
rect 31484 10047 31536 10056
rect 31484 10013 31493 10047
rect 31493 10013 31527 10047
rect 31527 10013 31536 10047
rect 31484 10004 31536 10013
rect 34336 10004 34388 10056
rect 17868 9936 17920 9988
rect 20260 9936 20312 9988
rect 20444 9936 20496 9988
rect 31392 9979 31444 9988
rect 31392 9945 31401 9979
rect 31401 9945 31435 9979
rect 31435 9945 31444 9979
rect 31392 9936 31444 9945
rect 38108 10047 38160 10056
rect 38108 10013 38117 10047
rect 38117 10013 38151 10047
rect 38151 10013 38160 10047
rect 38108 10004 38160 10013
rect 35072 9936 35124 9988
rect 6552 9868 6604 9920
rect 10140 9868 10192 9920
rect 13084 9911 13136 9920
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 13084 9868 13136 9877
rect 15844 9868 15896 9920
rect 18420 9868 18472 9920
rect 18604 9911 18656 9920
rect 18604 9877 18613 9911
rect 18613 9877 18647 9911
rect 18647 9877 18656 9911
rect 18604 9868 18656 9877
rect 19984 9868 20036 9920
rect 21548 9868 21600 9920
rect 21732 9911 21784 9920
rect 21732 9877 21741 9911
rect 21741 9877 21775 9911
rect 21775 9877 21784 9911
rect 21732 9868 21784 9877
rect 29920 9911 29972 9920
rect 29920 9877 29929 9911
rect 29929 9877 29963 9911
rect 29963 9877 29972 9911
rect 29920 9868 29972 9877
rect 30748 9911 30800 9920
rect 30748 9877 30757 9911
rect 30757 9877 30791 9911
rect 30791 9877 30800 9911
rect 30748 9868 30800 9877
rect 34520 9868 34572 9920
rect 36360 9911 36412 9920
rect 36360 9877 36369 9911
rect 36369 9877 36403 9911
rect 36403 9877 36412 9911
rect 36360 9868 36412 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2780 9664 2832 9716
rect 2872 9664 2924 9716
rect 4068 9664 4120 9716
rect 5816 9664 5868 9716
rect 10324 9664 10376 9716
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 4620 9596 4672 9648
rect 9312 9596 9364 9648
rect 20444 9596 20496 9648
rect 22100 9596 22152 9648
rect 30840 9664 30892 9716
rect 34796 9664 34848 9716
rect 35072 9596 35124 9648
rect 35348 9596 35400 9648
rect 5632 9571 5684 9580
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 2412 9392 2464 9444
rect 5632 9537 5641 9571
rect 5641 9537 5675 9571
rect 5675 9537 5684 9571
rect 5632 9528 5684 9537
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 12072 9528 12124 9580
rect 15476 9571 15528 9580
rect 15476 9537 15485 9571
rect 15485 9537 15519 9571
rect 15519 9537 15528 9571
rect 15476 9528 15528 9537
rect 15844 9528 15896 9580
rect 20628 9528 20680 9580
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 22652 9528 22704 9580
rect 28632 9571 28684 9580
rect 7380 9460 7432 9512
rect 9496 9503 9548 9512
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 11796 9503 11848 9512
rect 11796 9469 11805 9503
rect 11805 9469 11839 9503
rect 11839 9469 11848 9503
rect 11796 9460 11848 9469
rect 17408 9460 17460 9512
rect 26608 9460 26660 9512
rect 5540 9392 5592 9444
rect 5816 9392 5868 9444
rect 11060 9392 11112 9444
rect 27528 9460 27580 9512
rect 3056 9324 3108 9376
rect 4896 9324 4948 9376
rect 15292 9367 15344 9376
rect 15292 9333 15301 9367
rect 15301 9333 15335 9367
rect 15335 9333 15344 9367
rect 15292 9324 15344 9333
rect 15568 9324 15620 9376
rect 20352 9324 20404 9376
rect 28632 9537 28641 9571
rect 28641 9537 28675 9571
rect 28675 9537 28684 9571
rect 28632 9528 28684 9537
rect 29368 9460 29420 9512
rect 29920 9460 29972 9512
rect 34244 9571 34296 9580
rect 34244 9537 34253 9571
rect 34253 9537 34287 9571
rect 34287 9537 34296 9571
rect 34244 9528 34296 9537
rect 34428 9571 34480 9580
rect 34428 9537 34437 9571
rect 34437 9537 34471 9571
rect 34471 9537 34480 9571
rect 34428 9528 34480 9537
rect 34336 9503 34388 9512
rect 34336 9469 34345 9503
rect 34345 9469 34379 9503
rect 34379 9469 34388 9503
rect 34336 9460 34388 9469
rect 34520 9460 34572 9512
rect 33508 9367 33560 9376
rect 33508 9333 33517 9367
rect 33517 9333 33551 9367
rect 33551 9333 33560 9367
rect 33508 9324 33560 9333
rect 34612 9392 34664 9444
rect 34704 9324 34756 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3332 9120 3384 9172
rect 5632 9120 5684 9172
rect 20352 9120 20404 9172
rect 29552 9120 29604 9172
rect 29920 9120 29972 9172
rect 34520 9120 34572 9172
rect 1400 9095 1452 9104
rect 1400 9061 1409 9095
rect 1409 9061 1443 9095
rect 1443 9061 1452 9095
rect 1400 9052 1452 9061
rect 5172 9052 5224 9104
rect 9496 9052 9548 9104
rect 31300 9095 31352 9104
rect 31300 9061 31309 9095
rect 31309 9061 31343 9095
rect 31343 9061 31352 9095
rect 31300 9052 31352 9061
rect 34244 9052 34296 9104
rect 35624 9052 35676 9104
rect 5724 8984 5776 9036
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 16580 9027 16632 9036
rect 16580 8993 16589 9027
rect 16589 8993 16623 9027
rect 16623 8993 16632 9027
rect 16580 8984 16632 8993
rect 20628 8984 20680 9036
rect 27068 9027 27120 9036
rect 27068 8993 27077 9027
rect 27077 8993 27111 9027
rect 27111 8993 27120 9027
rect 27068 8984 27120 8993
rect 29092 8984 29144 9036
rect 30748 8984 30800 9036
rect 4896 8916 4948 8968
rect 5264 8916 5316 8968
rect 10968 8959 11020 8968
rect 10968 8925 10977 8959
rect 10977 8925 11011 8959
rect 11011 8925 11020 8959
rect 10968 8916 11020 8925
rect 11704 8916 11756 8968
rect 12624 8916 12676 8968
rect 15384 8959 15436 8968
rect 15384 8925 15393 8959
rect 15393 8925 15427 8959
rect 15427 8925 15436 8959
rect 15384 8916 15436 8925
rect 19984 8916 20036 8968
rect 20812 8916 20864 8968
rect 25228 8959 25280 8968
rect 25228 8925 25237 8959
rect 25237 8925 25271 8959
rect 25271 8925 25280 8959
rect 25228 8916 25280 8925
rect 30840 8916 30892 8968
rect 34796 8984 34848 9036
rect 35900 8984 35952 9036
rect 34704 8916 34756 8968
rect 35164 8959 35216 8968
rect 35164 8925 35173 8959
rect 35173 8925 35207 8959
rect 35207 8925 35216 8959
rect 35164 8916 35216 8925
rect 35256 8916 35308 8968
rect 36360 8984 36412 9036
rect 2596 8891 2648 8900
rect 2596 8857 2605 8891
rect 2605 8857 2639 8891
rect 2639 8857 2648 8891
rect 2596 8848 2648 8857
rect 2688 8848 2740 8900
rect 6552 8848 6604 8900
rect 20444 8848 20496 8900
rect 24032 8848 24084 8900
rect 29552 8848 29604 8900
rect 34612 8848 34664 8900
rect 5632 8780 5684 8832
rect 6920 8780 6972 8832
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 12164 8780 12216 8832
rect 19432 8780 19484 8832
rect 23756 8780 23808 8832
rect 30380 8823 30432 8832
rect 30380 8789 30389 8823
rect 30389 8789 30423 8823
rect 30423 8789 30432 8823
rect 30380 8780 30432 8789
rect 31668 8823 31720 8832
rect 31668 8789 31677 8823
rect 31677 8789 31711 8823
rect 31711 8789 31720 8823
rect 31668 8780 31720 8789
rect 34520 8780 34572 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 5632 8551 5684 8560
rect 5632 8517 5641 8551
rect 5641 8517 5675 8551
rect 5675 8517 5684 8551
rect 5632 8508 5684 8517
rect 5356 8440 5408 8492
rect 5816 8576 5868 8628
rect 6920 8619 6972 8628
rect 6920 8585 6929 8619
rect 6929 8585 6963 8619
rect 6963 8585 6972 8619
rect 6920 8576 6972 8585
rect 9220 8576 9272 8628
rect 11796 8508 11848 8560
rect 12164 8551 12216 8560
rect 12164 8517 12173 8551
rect 12173 8517 12207 8551
rect 12207 8517 12216 8551
rect 12164 8508 12216 8517
rect 13728 8508 13780 8560
rect 25136 8576 25188 8628
rect 25228 8576 25280 8628
rect 26056 8576 26108 8628
rect 28632 8576 28684 8628
rect 35348 8576 35400 8628
rect 22100 8508 22152 8560
rect 8300 8440 8352 8492
rect 23756 8483 23808 8492
rect 23756 8449 23765 8483
rect 23765 8449 23799 8483
rect 23799 8449 23808 8483
rect 23756 8440 23808 8449
rect 24032 8483 24084 8492
rect 24032 8449 24041 8483
rect 24041 8449 24075 8483
rect 24075 8449 24084 8483
rect 24032 8440 24084 8449
rect 5264 8372 5316 8424
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 4068 8304 4120 8356
rect 5172 8304 5224 8356
rect 6644 8236 6696 8288
rect 8760 8372 8812 8424
rect 10968 8415 11020 8424
rect 10968 8381 10977 8415
rect 10977 8381 11011 8415
rect 11011 8381 11020 8415
rect 10968 8372 11020 8381
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 16672 8347 16724 8356
rect 16672 8313 16681 8347
rect 16681 8313 16715 8347
rect 16715 8313 16724 8347
rect 16672 8304 16724 8313
rect 20720 8236 20772 8288
rect 25412 8440 25464 8492
rect 25872 8483 25924 8492
rect 25872 8449 25881 8483
rect 25881 8449 25915 8483
rect 25915 8449 25924 8483
rect 25872 8440 25924 8449
rect 25964 8440 26016 8492
rect 27252 8483 27304 8492
rect 27252 8449 27286 8483
rect 27286 8449 27304 8483
rect 27252 8440 27304 8449
rect 35164 8508 35216 8560
rect 35532 8551 35584 8560
rect 35532 8517 35541 8551
rect 35541 8517 35575 8551
rect 35575 8517 35584 8551
rect 35532 8508 35584 8517
rect 35900 8508 35952 8560
rect 30380 8440 30432 8492
rect 30932 8440 30984 8492
rect 34520 8483 34572 8492
rect 34520 8449 34529 8483
rect 34529 8449 34563 8483
rect 34563 8449 34572 8483
rect 34520 8440 34572 8449
rect 30472 8372 30524 8424
rect 33508 8372 33560 8424
rect 34152 8372 34204 8424
rect 35348 8440 35400 8492
rect 25044 8304 25096 8356
rect 28816 8347 28868 8356
rect 28816 8313 28825 8347
rect 28825 8313 28859 8347
rect 28859 8313 28868 8347
rect 28816 8304 28868 8313
rect 29368 8304 29420 8356
rect 33600 8304 33652 8356
rect 35440 8304 35492 8356
rect 35716 8347 35768 8356
rect 35716 8313 35725 8347
rect 35725 8313 35759 8347
rect 35759 8313 35768 8347
rect 35716 8304 35768 8313
rect 26976 8236 27028 8288
rect 30748 8279 30800 8288
rect 30748 8245 30757 8279
rect 30757 8245 30791 8279
rect 30791 8245 30800 8279
rect 30748 8236 30800 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2228 8032 2280 8084
rect 19340 8032 19392 8084
rect 3516 7964 3568 8016
rect 19432 7964 19484 8016
rect 5816 7896 5868 7948
rect 6644 7939 6696 7948
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 7564 7896 7616 7948
rect 11152 7939 11204 7948
rect 11152 7905 11161 7939
rect 11161 7905 11195 7939
rect 11195 7905 11204 7939
rect 11152 7896 11204 7905
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 15752 7939 15804 7948
rect 15752 7905 15761 7939
rect 15761 7905 15795 7939
rect 15795 7905 15804 7939
rect 15752 7896 15804 7905
rect 17132 7896 17184 7948
rect 28172 8032 28224 8084
rect 30472 8032 30524 8084
rect 35532 8032 35584 8084
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 10048 7760 10100 7812
rect 14556 7828 14608 7880
rect 16856 7760 16908 7812
rect 5448 7692 5500 7744
rect 18328 7692 18380 7744
rect 18604 7828 18656 7880
rect 19984 7896 20036 7948
rect 21732 7896 21784 7948
rect 25320 7939 25372 7948
rect 25320 7905 25329 7939
rect 25329 7905 25363 7939
rect 25363 7905 25372 7939
rect 25320 7896 25372 7905
rect 26608 7896 26660 7948
rect 25596 7828 25648 7880
rect 28724 7828 28776 7880
rect 35164 7871 35216 7880
rect 35164 7837 35173 7871
rect 35173 7837 35207 7871
rect 35207 7837 35216 7871
rect 35164 7828 35216 7837
rect 35348 7871 35400 7880
rect 35348 7837 35357 7871
rect 35357 7837 35391 7871
rect 35391 7837 35400 7871
rect 35348 7828 35400 7837
rect 35624 7828 35676 7880
rect 20444 7760 20496 7812
rect 21272 7760 21324 7812
rect 25964 7760 26016 7812
rect 20168 7692 20220 7744
rect 22284 7692 22336 7744
rect 35900 7692 35952 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 10048 7531 10100 7540
rect 10048 7497 10057 7531
rect 10057 7497 10091 7531
rect 10091 7497 10100 7531
rect 10048 7488 10100 7497
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 11428 7488 11480 7540
rect 19340 7488 19392 7540
rect 19984 7531 20036 7540
rect 19984 7497 19993 7531
rect 19993 7497 20027 7531
rect 20027 7497 20036 7531
rect 19984 7488 20036 7497
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 23112 7488 23164 7540
rect 24400 7488 24452 7540
rect 25872 7488 25924 7540
rect 26056 7531 26108 7540
rect 26056 7497 26065 7531
rect 26065 7497 26099 7531
rect 26099 7497 26108 7531
rect 26056 7488 26108 7497
rect 12624 7463 12676 7472
rect 12624 7429 12633 7463
rect 12633 7429 12667 7463
rect 12667 7429 12676 7463
rect 12624 7420 12676 7429
rect 14188 7420 14240 7472
rect 27252 7488 27304 7540
rect 5264 7352 5316 7404
rect 5448 7352 5500 7404
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 15568 7352 15620 7404
rect 17132 7352 17184 7404
rect 20628 7352 20680 7404
rect 21548 7352 21600 7404
rect 23112 7395 23164 7404
rect 23112 7361 23121 7395
rect 23121 7361 23155 7395
rect 23155 7361 23164 7395
rect 23112 7352 23164 7361
rect 27528 7420 27580 7472
rect 29184 7420 29236 7472
rect 29644 7463 29696 7472
rect 29644 7429 29653 7463
rect 29653 7429 29687 7463
rect 29687 7429 29696 7463
rect 29644 7420 29696 7429
rect 26608 7352 26660 7404
rect 26976 7395 27028 7404
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 7564 7216 7616 7268
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 20720 7327 20772 7336
rect 20720 7293 20729 7327
rect 20729 7293 20763 7327
rect 20763 7293 20772 7327
rect 20720 7284 20772 7293
rect 22100 7327 22152 7336
rect 22100 7293 22109 7327
rect 22109 7293 22143 7327
rect 22143 7293 22152 7327
rect 22100 7284 22152 7293
rect 15568 7216 15620 7268
rect 19340 7216 19392 7268
rect 25412 7284 25464 7336
rect 26976 7361 26985 7395
rect 26985 7361 27019 7395
rect 27019 7361 27028 7395
rect 26976 7352 27028 7361
rect 29276 7352 29328 7404
rect 35164 7488 35216 7540
rect 33600 7463 33652 7472
rect 33600 7429 33609 7463
rect 33609 7429 33643 7463
rect 33643 7429 33652 7463
rect 33600 7420 33652 7429
rect 30380 7395 30432 7404
rect 30380 7361 30389 7395
rect 30389 7361 30423 7395
rect 30423 7361 30432 7395
rect 30380 7352 30432 7361
rect 30472 7395 30524 7404
rect 30472 7361 30481 7395
rect 30481 7361 30515 7395
rect 30515 7361 30524 7395
rect 30472 7352 30524 7361
rect 30748 7352 30800 7404
rect 27068 7284 27120 7336
rect 28080 7284 28132 7336
rect 33600 7216 33652 7268
rect 4804 7148 4856 7200
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 23296 7191 23348 7200
rect 23296 7157 23305 7191
rect 23305 7157 23339 7191
rect 23339 7157 23348 7191
rect 23296 7148 23348 7157
rect 28632 7148 28684 7200
rect 29552 7148 29604 7200
rect 36176 7191 36228 7200
rect 36176 7157 36185 7191
rect 36185 7157 36219 7191
rect 36219 7157 36228 7191
rect 36176 7148 36228 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 23296 6944 23348 6996
rect 28632 6944 28684 6996
rect 30472 6944 30524 6996
rect 30564 6987 30616 6996
rect 30564 6953 30573 6987
rect 30573 6953 30607 6987
rect 30607 6953 30616 6987
rect 30564 6944 30616 6953
rect 28080 6876 28132 6928
rect 29276 6876 29328 6928
rect 30380 6876 30432 6928
rect 5172 6851 5224 6860
rect 5172 6817 5181 6851
rect 5181 6817 5215 6851
rect 5215 6817 5224 6851
rect 5172 6808 5224 6817
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4620 6740 4672 6792
rect 5356 6740 5408 6792
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8300 6783 8352 6792
rect 8024 6740 8076 6749
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 2688 6604 2740 6656
rect 2872 6604 2924 6656
rect 10232 6808 10284 6860
rect 15568 6851 15620 6860
rect 15568 6817 15577 6851
rect 15577 6817 15611 6851
rect 15611 6817 15620 6851
rect 15568 6808 15620 6817
rect 16488 6808 16540 6860
rect 26608 6851 26660 6860
rect 9680 6740 9732 6792
rect 15660 6740 15712 6792
rect 16856 6740 16908 6792
rect 17224 6740 17276 6792
rect 18420 6783 18472 6792
rect 18420 6749 18429 6783
rect 18429 6749 18463 6783
rect 18463 6749 18472 6783
rect 18420 6740 18472 6749
rect 26608 6817 26617 6851
rect 26617 6817 26651 6851
rect 26651 6817 26660 6851
rect 26608 6808 26660 6817
rect 33324 6808 33376 6860
rect 34152 6851 34204 6860
rect 34152 6817 34161 6851
rect 34161 6817 34195 6851
rect 34195 6817 34204 6851
rect 34152 6808 34204 6817
rect 22192 6783 22244 6792
rect 4896 6604 4948 6656
rect 5540 6604 5592 6656
rect 7932 6604 7984 6656
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 11980 6604 12032 6656
rect 15384 6604 15436 6656
rect 17868 6647 17920 6656
rect 17868 6613 17877 6647
rect 17877 6613 17911 6647
rect 17911 6613 17920 6647
rect 17868 6604 17920 6613
rect 20168 6715 20220 6724
rect 20168 6681 20177 6715
rect 20177 6681 20211 6715
rect 20211 6681 20220 6715
rect 20168 6672 20220 6681
rect 20720 6672 20772 6724
rect 21824 6672 21876 6724
rect 22192 6749 22201 6783
rect 22201 6749 22235 6783
rect 22235 6749 22244 6783
rect 22192 6740 22244 6749
rect 26148 6783 26200 6792
rect 26148 6749 26157 6783
rect 26157 6749 26191 6783
rect 26191 6749 26200 6783
rect 26148 6740 26200 6749
rect 27712 6740 27764 6792
rect 28724 6740 28776 6792
rect 30380 6783 30432 6792
rect 23296 6672 23348 6724
rect 30380 6749 30389 6783
rect 30389 6749 30423 6783
rect 30423 6749 30432 6783
rect 30380 6740 30432 6749
rect 30748 6740 30800 6792
rect 31760 6740 31812 6792
rect 32864 6672 32916 6724
rect 33600 6740 33652 6792
rect 34060 6783 34112 6792
rect 34060 6749 34069 6783
rect 34069 6749 34103 6783
rect 34103 6749 34112 6783
rect 34060 6740 34112 6749
rect 35716 6851 35768 6860
rect 35716 6817 35725 6851
rect 35725 6817 35759 6851
rect 35759 6817 35768 6851
rect 35716 6808 35768 6817
rect 35900 6851 35952 6860
rect 35900 6817 35909 6851
rect 35909 6817 35943 6851
rect 35943 6817 35952 6851
rect 35900 6808 35952 6817
rect 35624 6783 35676 6792
rect 35624 6749 35633 6783
rect 35633 6749 35667 6783
rect 35667 6749 35676 6783
rect 35624 6740 35676 6749
rect 20076 6647 20128 6656
rect 20076 6613 20085 6647
rect 20085 6613 20119 6647
rect 20119 6613 20128 6647
rect 20076 6604 20128 6613
rect 20444 6604 20496 6656
rect 25964 6647 26016 6656
rect 25964 6613 25973 6647
rect 25973 6613 26007 6647
rect 26007 6613 26016 6647
rect 25964 6604 26016 6613
rect 32220 6604 32272 6656
rect 36176 6672 36228 6724
rect 36452 6672 36504 6724
rect 35992 6604 36044 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 5816 6400 5868 6452
rect 8024 6400 8076 6452
rect 13728 6400 13780 6452
rect 14556 6443 14608 6452
rect 14556 6409 14565 6443
rect 14565 6409 14599 6443
rect 14599 6409 14608 6443
rect 14556 6400 14608 6409
rect 14924 6400 14976 6452
rect 15660 6400 15712 6452
rect 21824 6443 21876 6452
rect 21824 6409 21833 6443
rect 21833 6409 21867 6443
rect 21867 6409 21876 6443
rect 21824 6400 21876 6409
rect 3884 6332 3936 6384
rect 4804 6375 4856 6384
rect 4804 6341 4813 6375
rect 4813 6341 4847 6375
rect 4847 6341 4856 6375
rect 4804 6332 4856 6341
rect 2504 6307 2556 6316
rect 2504 6273 2538 6307
rect 2538 6273 2556 6307
rect 4620 6307 4672 6316
rect 2504 6264 2556 6273
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 5172 6332 5224 6384
rect 8300 6332 8352 6384
rect 14372 6332 14424 6384
rect 18420 6332 18472 6384
rect 20076 6332 20128 6384
rect 25596 6375 25648 6384
rect 25596 6341 25605 6375
rect 25605 6341 25639 6375
rect 25639 6341 25648 6375
rect 25596 6332 25648 6341
rect 34060 6400 34112 6452
rect 35624 6400 35676 6452
rect 36452 6443 36504 6452
rect 5540 6264 5592 6316
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 22284 6264 22336 6316
rect 23940 6307 23992 6316
rect 23940 6273 23949 6307
rect 23949 6273 23983 6307
rect 23983 6273 23992 6307
rect 23940 6264 23992 6273
rect 32220 6307 32272 6316
rect 32220 6273 32229 6307
rect 32229 6273 32263 6307
rect 32263 6273 32272 6307
rect 32220 6264 32272 6273
rect 35900 6332 35952 6384
rect 34796 6264 34848 6316
rect 35348 6264 35400 6316
rect 35992 6307 36044 6316
rect 10232 6196 10284 6248
rect 15568 6196 15620 6248
rect 16488 6196 16540 6248
rect 4160 6128 4212 6180
rect 4712 6128 4764 6180
rect 10968 6128 11020 6180
rect 14464 6128 14516 6180
rect 17040 6171 17092 6180
rect 17040 6137 17049 6171
rect 17049 6137 17083 6171
rect 17083 6137 17092 6171
rect 17040 6128 17092 6137
rect 21088 6128 21140 6180
rect 22192 6128 22244 6180
rect 30288 6196 30340 6248
rect 32496 6196 32548 6248
rect 33600 6196 33652 6248
rect 35992 6273 36001 6307
rect 36001 6273 36035 6307
rect 36035 6273 36044 6307
rect 35992 6264 36044 6273
rect 36452 6409 36461 6443
rect 36461 6409 36495 6443
rect 36495 6409 36504 6443
rect 36452 6400 36504 6409
rect 37832 6307 37884 6316
rect 37832 6273 37841 6307
rect 37841 6273 37875 6307
rect 37875 6273 37884 6307
rect 37832 6264 37884 6273
rect 29828 6128 29880 6180
rect 4620 6060 4672 6112
rect 14280 6060 14332 6112
rect 20720 6060 20772 6112
rect 20904 6103 20956 6112
rect 20904 6069 20913 6103
rect 20913 6069 20947 6103
rect 20947 6069 20956 6103
rect 20904 6060 20956 6069
rect 32220 6103 32272 6112
rect 32220 6069 32229 6103
rect 32229 6069 32263 6103
rect 32263 6069 32272 6103
rect 32220 6060 32272 6069
rect 38016 6103 38068 6112
rect 38016 6069 38025 6103
rect 38025 6069 38059 6103
rect 38059 6069 38068 6103
rect 38016 6060 38068 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2504 5856 2556 5908
rect 3976 5856 4028 5908
rect 10968 5856 11020 5908
rect 19708 5856 19760 5908
rect 4528 5788 4580 5840
rect 4896 5788 4948 5840
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 4712 5720 4764 5772
rect 5632 5720 5684 5772
rect 25964 5856 26016 5908
rect 20720 5788 20772 5840
rect 32220 5788 32272 5840
rect 5540 5652 5592 5704
rect 5816 5652 5868 5704
rect 3884 5559 3936 5568
rect 3884 5525 3893 5559
rect 3893 5525 3927 5559
rect 3927 5525 3936 5559
rect 3884 5516 3936 5525
rect 5172 5584 5224 5636
rect 15660 5720 15712 5772
rect 19432 5720 19484 5772
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 6736 5584 6788 5636
rect 14464 5627 14516 5636
rect 14464 5593 14473 5627
rect 14473 5593 14507 5627
rect 14507 5593 14516 5627
rect 14464 5584 14516 5593
rect 19340 5652 19392 5704
rect 19708 5695 19760 5704
rect 19708 5661 19717 5695
rect 19717 5661 19751 5695
rect 19751 5661 19760 5695
rect 19708 5652 19760 5661
rect 5816 5559 5868 5568
rect 5816 5525 5825 5559
rect 5825 5525 5859 5559
rect 5859 5525 5868 5559
rect 6644 5559 6696 5568
rect 5816 5516 5868 5525
rect 6644 5525 6653 5559
rect 6653 5525 6687 5559
rect 6687 5525 6696 5559
rect 6644 5516 6696 5525
rect 7932 5516 7984 5568
rect 10324 5559 10376 5568
rect 10324 5525 10333 5559
rect 10333 5525 10367 5559
rect 10367 5525 10376 5559
rect 10324 5516 10376 5525
rect 14280 5516 14332 5568
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 19248 5559 19300 5568
rect 19248 5525 19257 5559
rect 19257 5525 19291 5559
rect 19291 5525 19300 5559
rect 19248 5516 19300 5525
rect 19340 5516 19392 5568
rect 19892 5720 19944 5772
rect 23756 5720 23808 5772
rect 26148 5720 26200 5772
rect 20444 5695 20496 5704
rect 20444 5661 20453 5695
rect 20453 5661 20487 5695
rect 20487 5661 20496 5695
rect 20444 5652 20496 5661
rect 19892 5584 19944 5636
rect 20720 5584 20772 5636
rect 26792 5652 26844 5704
rect 29092 5720 29144 5772
rect 30288 5763 30340 5772
rect 30288 5729 30297 5763
rect 30297 5729 30331 5763
rect 30331 5729 30340 5763
rect 30288 5720 30340 5729
rect 30564 5720 30616 5772
rect 30380 5652 30432 5704
rect 20628 5559 20680 5568
rect 20628 5525 20637 5559
rect 20637 5525 20671 5559
rect 20671 5525 20680 5559
rect 20628 5516 20680 5525
rect 22192 5627 22244 5636
rect 22192 5593 22201 5627
rect 22201 5593 22235 5627
rect 22235 5593 22244 5627
rect 22192 5584 22244 5593
rect 24768 5584 24820 5636
rect 27804 5584 27856 5636
rect 29828 5584 29880 5636
rect 23480 5516 23532 5568
rect 30656 5584 30708 5636
rect 31024 5516 31076 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2596 5312 2648 5364
rect 4528 5355 4580 5364
rect 4528 5321 4537 5355
rect 4537 5321 4571 5355
rect 4571 5321 4580 5355
rect 4528 5312 4580 5321
rect 8760 5355 8812 5364
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 14556 5312 14608 5364
rect 15476 5355 15528 5364
rect 15476 5321 15485 5355
rect 15485 5321 15519 5355
rect 15519 5321 15528 5355
rect 15476 5312 15528 5321
rect 19432 5312 19484 5364
rect 20720 5355 20772 5364
rect 20720 5321 20729 5355
rect 20729 5321 20763 5355
rect 20763 5321 20772 5355
rect 20720 5312 20772 5321
rect 26332 5355 26384 5364
rect 26332 5321 26341 5355
rect 26341 5321 26375 5355
rect 26375 5321 26384 5355
rect 26332 5312 26384 5321
rect 28448 5355 28500 5364
rect 28448 5321 28457 5355
rect 28457 5321 28491 5355
rect 28491 5321 28500 5355
rect 28448 5312 28500 5321
rect 29828 5355 29880 5364
rect 29828 5321 29837 5355
rect 29837 5321 29871 5355
rect 29871 5321 29880 5355
rect 29828 5312 29880 5321
rect 30564 5312 30616 5364
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 4620 5176 4672 5228
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 5540 5219 5592 5228
rect 4160 5108 4212 5160
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 6644 5176 6696 5228
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 5724 5108 5776 5160
rect 6736 5108 6788 5160
rect 4528 5040 4580 5092
rect 9036 5151 9088 5160
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 10324 5151 10376 5160
rect 9036 5108 9088 5117
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 9772 5040 9824 5092
rect 10784 5176 10836 5228
rect 12532 5176 12584 5228
rect 19248 5244 19300 5296
rect 19340 5244 19392 5296
rect 20260 5244 20312 5296
rect 15844 5176 15896 5228
rect 17040 5176 17092 5228
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 19708 5176 19760 5228
rect 15660 5108 15712 5160
rect 25044 5108 25096 5160
rect 27712 5151 27764 5160
rect 27712 5117 27721 5151
rect 27721 5117 27755 5151
rect 27755 5117 27764 5151
rect 27712 5108 27764 5117
rect 29092 5108 29144 5160
rect 3240 4972 3292 5024
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 10692 4972 10744 5024
rect 15200 5040 15252 5092
rect 26332 5040 26384 5092
rect 15292 4972 15344 5024
rect 15936 5015 15988 5024
rect 15936 4981 15945 5015
rect 15945 4981 15979 5015
rect 15979 4981 15988 5015
rect 15936 4972 15988 4981
rect 19156 4972 19208 5024
rect 26976 4972 27028 5024
rect 34704 5015 34756 5024
rect 34704 4981 34713 5015
rect 34713 4981 34747 5015
rect 34747 4981 34756 5015
rect 34704 4972 34756 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4620 4768 4672 4820
rect 5816 4768 5868 4820
rect 5172 4700 5224 4752
rect 14464 4768 14516 4820
rect 15844 4811 15896 4820
rect 15844 4777 15853 4811
rect 15853 4777 15887 4811
rect 15887 4777 15896 4811
rect 15844 4768 15896 4777
rect 19708 4811 19760 4820
rect 19708 4777 19717 4811
rect 19717 4777 19751 4811
rect 19751 4777 19760 4811
rect 19708 4768 19760 4777
rect 23756 4811 23808 4820
rect 23756 4777 23765 4811
rect 23765 4777 23799 4811
rect 23799 4777 23808 4811
rect 23756 4768 23808 4777
rect 24768 4768 24820 4820
rect 35900 4768 35952 4820
rect 6644 4632 6696 4684
rect 7380 4632 7432 4684
rect 9036 4632 9088 4684
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 4988 4564 5040 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 10784 4632 10836 4684
rect 7288 4564 7340 4573
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10692 4607 10744 4616
rect 10508 4564 10560 4573
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 12440 4743 12492 4752
rect 12440 4709 12449 4743
rect 12449 4709 12483 4743
rect 12483 4709 12492 4743
rect 12440 4700 12492 4709
rect 17132 4700 17184 4752
rect 14648 4632 14700 4684
rect 15200 4675 15252 4684
rect 15200 4641 15209 4675
rect 15209 4641 15243 4675
rect 15243 4641 15252 4675
rect 15200 4632 15252 4641
rect 15936 4632 15988 4684
rect 22928 4632 22980 4684
rect 25044 4675 25096 4684
rect 25044 4641 25053 4675
rect 25053 4641 25087 4675
rect 25087 4641 25096 4675
rect 25044 4632 25096 4641
rect 11888 4607 11940 4616
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14556 4564 14608 4616
rect 17868 4564 17920 4616
rect 18236 4607 18288 4616
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 20996 4607 21048 4616
rect 20996 4573 21005 4607
rect 21005 4573 21039 4607
rect 21039 4573 21048 4607
rect 37740 4700 37792 4752
rect 26792 4675 26844 4684
rect 26792 4641 26801 4675
rect 26801 4641 26835 4675
rect 26835 4641 26844 4675
rect 26792 4632 26844 4641
rect 28080 4675 28132 4684
rect 28080 4641 28089 4675
rect 28089 4641 28123 4675
rect 28123 4641 28132 4675
rect 28080 4632 28132 4641
rect 29092 4632 29144 4684
rect 34612 4632 34664 4684
rect 26976 4607 27028 4616
rect 20996 4564 21048 4573
rect 26976 4573 26985 4607
rect 26985 4573 27019 4607
rect 27019 4573 27028 4607
rect 26976 4564 27028 4573
rect 31024 4607 31076 4616
rect 31024 4573 31033 4607
rect 31033 4573 31067 4607
rect 31067 4573 31076 4607
rect 31024 4564 31076 4573
rect 34796 4607 34848 4616
rect 34796 4573 34838 4607
rect 34838 4573 34848 4607
rect 34796 4564 34848 4573
rect 5448 4496 5500 4548
rect 3148 4428 3200 4480
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 7380 4496 7432 4548
rect 10784 4539 10836 4548
rect 10784 4505 10793 4539
rect 10793 4505 10827 4539
rect 10827 4505 10836 4539
rect 10784 4496 10836 4505
rect 16396 4496 16448 4548
rect 16856 4496 16908 4548
rect 23480 4496 23532 4548
rect 29184 4496 29236 4548
rect 11520 4471 11572 4480
rect 11520 4437 11529 4471
rect 11529 4437 11563 4471
rect 11563 4437 11572 4471
rect 11520 4428 11572 4437
rect 13820 4428 13872 4480
rect 17316 4428 17368 4480
rect 24676 4428 24728 4480
rect 24768 4471 24820 4480
rect 24768 4437 24777 4471
rect 24777 4437 24811 4471
rect 24811 4437 24820 4471
rect 27620 4471 27672 4480
rect 24768 4428 24820 4437
rect 27620 4437 27629 4471
rect 27629 4437 27663 4471
rect 27663 4437 27672 4471
rect 27620 4428 27672 4437
rect 29092 4428 29144 4480
rect 31208 4471 31260 4480
rect 31208 4437 31217 4471
rect 31217 4437 31251 4471
rect 31251 4437 31260 4471
rect 31208 4428 31260 4437
rect 34520 4428 34572 4480
rect 34796 4428 34848 4480
rect 35808 4471 35860 4480
rect 35808 4437 35817 4471
rect 35817 4437 35851 4471
rect 35851 4437 35860 4471
rect 35808 4428 35860 4437
rect 36268 4428 36320 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 5448 4224 5500 4276
rect 11612 4224 11664 4276
rect 11888 4224 11940 4276
rect 14648 4267 14700 4276
rect 14648 4233 14657 4267
rect 14657 4233 14691 4267
rect 14691 4233 14700 4267
rect 14648 4224 14700 4233
rect 15476 4224 15528 4276
rect 27712 4224 27764 4276
rect 4068 4156 4120 4208
rect 10784 4156 10836 4208
rect 15292 4156 15344 4208
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 3148 4131 3200 4140
rect 3148 4097 3182 4131
rect 3182 4097 3200 4131
rect 3148 4088 3200 4097
rect 4436 4088 4488 4140
rect 7932 4131 7984 4140
rect 7932 4097 7941 4131
rect 7941 4097 7975 4131
rect 7975 4097 7984 4131
rect 7932 4088 7984 4097
rect 11520 4088 11572 4140
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 15384 4131 15436 4140
rect 15384 4097 15393 4131
rect 15393 4097 15427 4131
rect 15427 4097 15436 4131
rect 15384 4088 15436 4097
rect 17316 4131 17368 4140
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 17316 4088 17368 4097
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 23480 4131 23532 4140
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 15200 4063 15252 4072
rect 15200 4029 15209 4063
rect 15209 4029 15243 4063
rect 15243 4029 15252 4063
rect 15200 4020 15252 4029
rect 18236 4020 18288 4072
rect 2412 3952 2464 4004
rect 15660 3952 15712 4004
rect 23480 4097 23489 4131
rect 23489 4097 23523 4131
rect 23523 4097 23532 4131
rect 23480 4088 23532 4097
rect 23664 4131 23716 4140
rect 23664 4097 23673 4131
rect 23673 4097 23707 4131
rect 23707 4097 23716 4131
rect 23664 4088 23716 4097
rect 24676 4131 24728 4140
rect 24676 4097 24685 4131
rect 24685 4097 24719 4131
rect 24719 4097 24728 4131
rect 24676 4088 24728 4097
rect 23756 4063 23808 4072
rect 23756 4029 23765 4063
rect 23765 4029 23799 4063
rect 23799 4029 23808 4063
rect 23756 4020 23808 4029
rect 26792 4088 26844 4140
rect 27620 4088 27672 4140
rect 28816 4088 28868 4140
rect 29092 4131 29144 4140
rect 29092 4097 29110 4131
rect 29110 4097 29144 4131
rect 29092 4088 29144 4097
rect 29644 4088 29696 4140
rect 33876 4131 33928 4140
rect 33876 4097 33885 4131
rect 33885 4097 33919 4131
rect 33919 4097 33928 4131
rect 33876 4088 33928 4097
rect 34520 4088 34572 4140
rect 35440 4088 35492 4140
rect 31116 4020 31168 4072
rect 31760 4020 31812 4072
rect 34704 4020 34756 4072
rect 4712 3927 4764 3936
rect 4712 3893 4721 3927
rect 4721 3893 4755 3927
rect 4755 3893 4764 3927
rect 4712 3884 4764 3893
rect 5724 3884 5776 3936
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 10876 3884 10928 3936
rect 13452 3884 13504 3936
rect 17500 3927 17552 3936
rect 17500 3893 17509 3927
rect 17509 3893 17543 3927
rect 17543 3893 17552 3927
rect 17500 3884 17552 3893
rect 19892 3884 19944 3936
rect 24584 3884 24636 3936
rect 27620 3884 27672 3936
rect 34060 3927 34112 3936
rect 34060 3893 34069 3927
rect 34069 3893 34103 3927
rect 34103 3893 34112 3927
rect 34060 3884 34112 3893
rect 36268 3927 36320 3936
rect 36268 3893 36277 3927
rect 36277 3893 36311 3927
rect 36311 3893 36320 3927
rect 36268 3884 36320 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 6828 3612 6880 3664
rect 9772 3655 9824 3664
rect 9772 3621 9781 3655
rect 9781 3621 9815 3655
rect 9815 3621 9824 3655
rect 9772 3612 9824 3621
rect 11244 3680 11296 3732
rect 15752 3680 15804 3732
rect 16396 3723 16448 3732
rect 16396 3689 16405 3723
rect 16405 3689 16439 3723
rect 16439 3689 16448 3723
rect 16396 3680 16448 3689
rect 19340 3680 19392 3732
rect 20996 3723 21048 3732
rect 20996 3689 21005 3723
rect 21005 3689 21039 3723
rect 21039 3689 21048 3723
rect 20996 3680 21048 3689
rect 22928 3723 22980 3732
rect 22928 3689 22937 3723
rect 22937 3689 22971 3723
rect 22971 3689 22980 3723
rect 22928 3680 22980 3689
rect 29644 3723 29696 3732
rect 13084 3544 13136 3596
rect 23756 3612 23808 3664
rect 23480 3587 23532 3596
rect 23480 3553 23489 3587
rect 23489 3553 23523 3587
rect 23523 3553 23532 3587
rect 23480 3544 23532 3553
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 2872 3476 2924 3528
rect 3884 3476 3936 3528
rect 5724 3476 5776 3528
rect 10876 3519 10928 3528
rect 10876 3485 10894 3519
rect 10894 3485 10928 3519
rect 10876 3476 10928 3485
rect 4712 3408 4764 3460
rect 3976 3340 4028 3392
rect 11244 3408 11296 3460
rect 17500 3519 17552 3528
rect 17500 3485 17518 3519
rect 17518 3485 17552 3519
rect 17776 3519 17828 3528
rect 17500 3476 17552 3485
rect 17776 3485 17785 3519
rect 17785 3485 17819 3519
rect 17819 3485 17828 3519
rect 17776 3476 17828 3485
rect 19892 3519 19944 3528
rect 19892 3485 19926 3519
rect 19926 3485 19944 3519
rect 19892 3476 19944 3485
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 29644 3689 29653 3723
rect 29653 3689 29687 3723
rect 29687 3689 29696 3723
rect 29644 3680 29696 3689
rect 32496 3723 32548 3732
rect 29276 3612 29328 3664
rect 32496 3689 32505 3723
rect 32505 3689 32539 3723
rect 32539 3689 32548 3723
rect 32496 3680 32548 3689
rect 34612 3680 34664 3732
rect 35440 3680 35492 3732
rect 31116 3587 31168 3596
rect 31116 3553 31125 3587
rect 31125 3553 31159 3587
rect 31159 3553 31168 3587
rect 31116 3544 31168 3553
rect 36268 3544 36320 3596
rect 23664 3408 23716 3460
rect 5724 3383 5776 3392
rect 5724 3349 5733 3383
rect 5733 3349 5767 3383
rect 5767 3349 5776 3383
rect 5724 3340 5776 3349
rect 11704 3383 11756 3392
rect 11704 3349 11713 3383
rect 11713 3349 11747 3383
rect 11747 3349 11756 3383
rect 11704 3340 11756 3349
rect 24400 3383 24452 3392
rect 24400 3349 24409 3383
rect 24409 3349 24443 3383
rect 24443 3349 24452 3383
rect 24400 3340 24452 3349
rect 27896 3451 27948 3460
rect 27896 3417 27930 3451
rect 27930 3417 27948 3451
rect 27896 3408 27948 3417
rect 31208 3408 31260 3460
rect 34704 3408 34756 3460
rect 33876 3340 33928 3392
rect 35808 3476 35860 3528
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 9312 3136 9364 3188
rect 14556 3179 14608 3188
rect 14556 3145 14565 3179
rect 14565 3145 14599 3179
rect 14599 3145 14608 3179
rect 14556 3136 14608 3145
rect 5724 3068 5776 3120
rect 11704 3068 11756 3120
rect 2780 2864 2832 2916
rect 2688 2796 2740 2848
rect 2964 2796 3016 2848
rect 7748 3043 7800 3052
rect 7748 3009 7782 3043
rect 7782 3009 7800 3043
rect 7748 3000 7800 3009
rect 16672 3068 16724 3120
rect 17776 3068 17828 3120
rect 20904 3068 20956 3120
rect 13452 3043 13504 3052
rect 13452 3009 13486 3043
rect 13486 3009 13504 3043
rect 13452 3000 13504 3009
rect 23480 3136 23532 3188
rect 27896 3136 27948 3188
rect 31116 3136 31168 3188
rect 34704 3179 34756 3188
rect 24400 3068 24452 3120
rect 31392 3068 31444 3120
rect 27620 3043 27672 3052
rect 27620 3009 27629 3043
rect 27629 3009 27663 3043
rect 27663 3009 27672 3043
rect 27620 3000 27672 3009
rect 34704 3145 34713 3179
rect 34713 3145 34747 3179
rect 34747 3145 34756 3179
rect 34704 3136 34756 3145
rect 34060 3068 34112 3120
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3056 2592 3108 2644
rect 2964 2456 3016 2508
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 34612 2388 34664 2440
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 13360 2320 13412 2372
rect 38016 2295 38068 2304
rect 38016 2261 38025 2295
rect 38025 2261 38059 2295
rect 38059 2261 38068 2295
rect 38016 2252 38068 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 3422 39672 3478 39681
rect 3422 39607 3478 39616
rect 3148 36576 3200 36582
rect 3148 36518 3200 36524
rect 3160 34610 3188 36518
rect 3332 36100 3384 36106
rect 3332 36042 3384 36048
rect 3344 35290 3372 36042
rect 3332 35284 3384 35290
rect 3332 35226 3384 35232
rect 3148 34604 3200 34610
rect 3148 34546 3200 34552
rect 2780 34400 2832 34406
rect 2780 34342 2832 34348
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1412 33561 1440 33934
rect 2688 33856 2740 33862
rect 2688 33798 2740 33804
rect 1398 33552 1454 33561
rect 1398 33487 1454 33496
rect 1400 32428 1452 32434
rect 1400 32370 1452 32376
rect 1412 32201 1440 32370
rect 1584 32224 1636 32230
rect 1398 32192 1454 32201
rect 1584 32166 1636 32172
rect 1398 32127 1454 32136
rect 1596 31414 1624 32166
rect 1584 31408 1636 31414
rect 1584 31350 1636 31356
rect 1400 31340 1452 31346
rect 1400 31282 1452 31288
rect 1412 30870 1440 31282
rect 2700 31142 2728 33798
rect 2792 33454 2820 34342
rect 2780 33448 2832 33454
rect 2780 33390 2832 33396
rect 2964 33448 3016 33454
rect 2964 33390 3016 33396
rect 2976 32978 3004 33390
rect 2964 32972 3016 32978
rect 2964 32914 3016 32920
rect 2872 32360 2924 32366
rect 2872 32302 2924 32308
rect 3056 32360 3108 32366
rect 3056 32302 3108 32308
rect 2884 32026 2912 32302
rect 2872 32020 2924 32026
rect 2872 31962 2924 31968
rect 3068 31482 3096 32302
rect 3056 31476 3108 31482
rect 3056 31418 3108 31424
rect 2688 31136 2740 31142
rect 2688 31078 2740 31084
rect 2780 31136 2832 31142
rect 2780 31078 2832 31084
rect 1400 30864 1452 30870
rect 1398 30832 1400 30841
rect 1452 30832 1454 30841
rect 1398 30767 1454 30776
rect 2792 29850 2820 31078
rect 2780 29844 2832 29850
rect 2780 29786 2832 29792
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1412 29481 1440 29582
rect 1398 29472 1454 29481
rect 1398 29407 1454 29416
rect 3238 28792 3294 28801
rect 3238 28727 3294 28736
rect 1400 28552 1452 28558
rect 1400 28494 1452 28500
rect 2780 28552 2832 28558
rect 2780 28494 2832 28500
rect 1412 28150 1440 28494
rect 2596 28416 2648 28422
rect 2596 28358 2648 28364
rect 1400 28144 1452 28150
rect 1398 28112 1400 28121
rect 1452 28112 1454 28121
rect 1398 28047 1454 28056
rect 1400 26988 1452 26994
rect 1400 26930 1452 26936
rect 1412 26761 1440 26930
rect 1584 26784 1636 26790
rect 1398 26752 1454 26761
rect 1584 26726 1636 26732
rect 1398 26687 1454 26696
rect 1596 25906 1624 26726
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1412 25430 1440 25842
rect 2608 25702 2636 28358
rect 2792 28082 2820 28494
rect 2780 28076 2832 28082
rect 2780 28018 2832 28024
rect 3252 28014 3280 28727
rect 2964 28008 3016 28014
rect 2964 27950 3016 27956
rect 3240 28008 3292 28014
rect 3240 27950 3292 27956
rect 2976 27674 3004 27950
rect 2964 27668 3016 27674
rect 2964 27610 3016 27616
rect 2964 26036 3016 26042
rect 2964 25978 3016 25984
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 2596 25696 2648 25702
rect 2596 25638 2648 25644
rect 1400 25424 1452 25430
rect 1398 25392 1400 25401
rect 1452 25392 1454 25401
rect 1398 25327 1454 25336
rect 2596 25288 2648 25294
rect 2596 25230 2648 25236
rect 2608 24818 2636 25230
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 2792 24886 2820 25094
rect 2780 24880 2832 24886
rect 2780 24822 2832 24828
rect 2596 24812 2648 24818
rect 2596 24754 2648 24760
rect 2884 24410 2912 25842
rect 2872 24404 2924 24410
rect 2872 24346 2924 24352
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 24041 1440 24142
rect 1398 24032 1454 24041
rect 1398 23967 1454 23976
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 2976 23066 3004 25978
rect 3240 25288 3292 25294
rect 3240 25230 3292 25236
rect 3056 24744 3108 24750
rect 3054 24712 3056 24721
rect 3108 24712 3110 24721
rect 3054 24647 3110 24656
rect 3068 24342 3096 24647
rect 3252 24410 3280 25230
rect 3436 24614 3464 39607
rect 9692 39222 9904 39250
rect 3606 38992 3662 39001
rect 3606 38927 3662 38936
rect 3620 31414 3648 38927
rect 3698 38312 3754 38321
rect 3698 38247 3754 38256
rect 3712 34406 3740 38247
rect 3974 37632 4030 37641
rect 3974 37567 4030 37576
rect 3790 36952 3846 36961
rect 3790 36887 3846 36896
rect 3804 36310 3832 36887
rect 3988 36854 4016 37567
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 3976 36848 4028 36854
rect 3976 36790 4028 36796
rect 4068 36644 4120 36650
rect 4068 36586 4120 36592
rect 3884 36576 3936 36582
rect 3884 36518 3936 36524
rect 3792 36304 3844 36310
rect 3792 36246 3844 36252
rect 3792 35624 3844 35630
rect 3792 35566 3844 35572
rect 3804 35290 3832 35566
rect 3792 35284 3844 35290
rect 3792 35226 3844 35232
rect 3896 34678 3924 36518
rect 4080 36281 4108 36586
rect 4712 36576 4764 36582
rect 4712 36518 4764 36524
rect 8944 36576 8996 36582
rect 8944 36518 8996 36524
rect 9128 36576 9180 36582
rect 9128 36518 9180 36524
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4066 36272 4122 36281
rect 4066 36207 4122 36216
rect 4066 35592 4122 35601
rect 4066 35527 4068 35536
rect 4120 35527 4122 35536
rect 4068 35498 4120 35504
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4724 35018 4752 36518
rect 8956 36242 8984 36518
rect 5264 36236 5316 36242
rect 5264 36178 5316 36184
rect 8944 36236 8996 36242
rect 8944 36178 8996 36184
rect 5276 35766 5304 36178
rect 7564 36168 7616 36174
rect 7564 36110 7616 36116
rect 5264 35760 5316 35766
rect 5264 35702 5316 35708
rect 4344 35012 4396 35018
rect 4344 34954 4396 34960
rect 4712 35012 4764 35018
rect 4712 34954 4764 34960
rect 4068 34944 4120 34950
rect 4066 34912 4068 34921
rect 4120 34912 4122 34921
rect 4066 34847 4122 34856
rect 3884 34672 3936 34678
rect 3884 34614 3936 34620
rect 4356 34542 4384 34954
rect 4344 34536 4396 34542
rect 4344 34478 4396 34484
rect 4620 34536 4672 34542
rect 4620 34478 4672 34484
rect 4068 34468 4120 34474
rect 4068 34410 4120 34416
rect 3700 34400 3752 34406
rect 3700 34342 3752 34348
rect 4080 34241 4108 34410
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4066 34232 4122 34241
rect 4214 34224 4522 34244
rect 4066 34167 4122 34176
rect 4632 34066 4660 34478
rect 4620 34060 4672 34066
rect 4620 34002 4672 34008
rect 4632 33590 4660 34002
rect 4620 33584 4672 33590
rect 4620 33526 4672 33532
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 3792 32904 3844 32910
rect 3792 32846 3844 32852
rect 4066 32872 4122 32881
rect 3608 31408 3660 31414
rect 3608 31350 3660 31356
rect 3608 31136 3660 31142
rect 3608 31078 3660 31084
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3240 24404 3292 24410
rect 3240 24346 3292 24352
rect 3056 24336 3108 24342
rect 3056 24278 3108 24284
rect 3238 23352 3294 23361
rect 3238 23287 3294 23296
rect 1412 22710 1440 23054
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1400 22704 1452 22710
rect 1398 22672 1400 22681
rect 1452 22672 1454 22681
rect 1398 22607 1454 22616
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 21321 1440 21490
rect 1398 21312 1454 21321
rect 1398 21247 1454 21256
rect 1400 20460 1452 20466
rect 1400 20402 1452 20408
rect 1412 19961 1440 20402
rect 1398 19952 1454 19961
rect 1398 19887 1454 19896
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1412 18601 1440 18702
rect 1398 18592 1454 18601
rect 1398 18527 1454 18536
rect 1596 17882 1624 22918
rect 2792 22642 2820 23054
rect 2976 23038 3096 23066
rect 2964 22976 3016 22982
rect 2964 22918 3016 22924
rect 2976 22710 3004 22918
rect 2964 22704 3016 22710
rect 2964 22646 3016 22652
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2700 21554 2728 21966
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2332 18290 2360 20198
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2424 19378 2452 19790
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 2136 17876 2188 17882
rect 2136 17818 2188 17824
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1412 17270 1440 17614
rect 1400 17264 1452 17270
rect 1398 17232 1400 17241
rect 1452 17232 1454 17241
rect 1398 17167 1454 17176
rect 2148 16998 2176 17818
rect 2332 17134 2360 18226
rect 2516 17678 2544 21286
rect 2596 20256 2648 20262
rect 2596 20198 2648 20204
rect 2608 19446 2636 20198
rect 2596 19440 2648 19446
rect 2596 19382 2648 19388
rect 2872 19304 2924 19310
rect 2870 19272 2872 19281
rect 2924 19272 2926 19281
rect 2870 19207 2926 19216
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2608 17746 2636 18566
rect 2884 18426 2912 19207
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 3068 17882 3096 23038
rect 3252 22574 3280 23287
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2608 17626 2636 17682
rect 2516 17202 2544 17614
rect 2608 17598 2728 17626
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2320 17128 2372 17134
rect 2320 17070 2372 17076
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2424 16522 2452 16934
rect 2516 16590 2544 17138
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2412 16516 2464 16522
rect 2412 16458 2464 16464
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 15881 1440 16050
rect 2504 15904 2556 15910
rect 1398 15872 1454 15881
rect 2504 15846 2556 15852
rect 1398 15807 1454 15816
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1412 14521 1440 14962
rect 1398 14512 1454 14521
rect 1398 14447 1454 14456
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 13161 1440 13262
rect 1584 13184 1636 13190
rect 1398 13152 1454 13161
rect 1584 13126 1636 13132
rect 1398 13087 1454 13096
rect 1596 12646 1624 13126
rect 2516 12918 2544 15846
rect 2504 12912 2556 12918
rect 2504 12854 2556 12860
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2424 12306 2452 12582
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2516 12238 2544 12854
rect 2608 12782 2636 17478
rect 2700 17202 2728 17598
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2884 16590 2912 16934
rect 2976 16794 3004 17206
rect 3068 17134 3096 17818
rect 3252 17746 3280 18022
rect 3620 17814 3648 31078
rect 3804 29850 3832 32846
rect 4066 32807 4122 32816
rect 3884 31340 3936 31346
rect 3884 31282 3936 31288
rect 3896 30394 3924 31282
rect 4080 31210 4108 32807
rect 5276 32502 5304 35702
rect 7576 35698 7604 36110
rect 7564 35692 7616 35698
rect 7564 35634 7616 35640
rect 8024 35624 8076 35630
rect 8024 35566 8076 35572
rect 8036 35290 8064 35566
rect 8024 35284 8076 35290
rect 8024 35226 8076 35232
rect 9140 35154 9168 36518
rect 9312 35488 9364 35494
rect 9312 35430 9364 35436
rect 9324 35154 9352 35430
rect 6000 35148 6052 35154
rect 6000 35090 6052 35096
rect 9128 35148 9180 35154
rect 9128 35090 9180 35096
rect 9312 35148 9364 35154
rect 9312 35090 9364 35096
rect 6012 34202 6040 35090
rect 6736 35080 6788 35086
rect 6736 35022 6788 35028
rect 8116 35080 8168 35086
rect 8116 35022 8168 35028
rect 6748 34746 6776 35022
rect 8128 34746 8156 35022
rect 6736 34740 6788 34746
rect 6736 34682 6788 34688
rect 8116 34740 8168 34746
rect 8116 34682 8168 34688
rect 8024 34672 8076 34678
rect 8024 34614 8076 34620
rect 7472 34604 7524 34610
rect 7472 34546 7524 34552
rect 6276 34400 6328 34406
rect 6276 34342 6328 34348
rect 6000 34196 6052 34202
rect 6000 34138 6052 34144
rect 6288 34066 6316 34342
rect 6276 34060 6328 34066
rect 6276 34002 6328 34008
rect 7484 33998 7512 34546
rect 7932 34468 7984 34474
rect 7932 34410 7984 34416
rect 7656 34400 7708 34406
rect 7708 34360 7788 34388
rect 7656 34342 7708 34348
rect 7760 34202 7788 34360
rect 7748 34196 7800 34202
rect 7748 34138 7800 34144
rect 7472 33992 7524 33998
rect 7472 33934 7524 33940
rect 6092 33924 6144 33930
rect 6092 33866 6144 33872
rect 5264 32496 5316 32502
rect 5264 32438 5316 32444
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 5276 31890 5304 32438
rect 5816 32224 5868 32230
rect 5816 32166 5868 32172
rect 5828 31890 5856 32166
rect 6104 31890 6132 33866
rect 7484 33522 7512 33934
rect 7472 33516 7524 33522
rect 7472 33458 7524 33464
rect 7760 33386 7788 34138
rect 7944 34066 7972 34410
rect 7932 34060 7984 34066
rect 7932 34002 7984 34008
rect 7944 33454 7972 34002
rect 8036 33930 8064 34614
rect 8024 33924 8076 33930
rect 8024 33866 8076 33872
rect 8036 33590 8064 33866
rect 8024 33584 8076 33590
rect 8024 33526 8076 33532
rect 7932 33448 7984 33454
rect 7932 33390 7984 33396
rect 7748 33380 7800 33386
rect 7748 33322 7800 33328
rect 7104 33312 7156 33318
rect 7104 33254 7156 33260
rect 7564 33312 7616 33318
rect 7564 33254 7616 33260
rect 7116 32434 7144 33254
rect 7576 32910 7604 33254
rect 7564 32904 7616 32910
rect 7564 32846 7616 32852
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 7392 32502 7420 32710
rect 7380 32496 7432 32502
rect 7380 32438 7432 32444
rect 7104 32428 7156 32434
rect 7104 32370 7156 32376
rect 4160 31884 4212 31890
rect 4160 31826 4212 31832
rect 5264 31884 5316 31890
rect 5264 31826 5316 31832
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 6092 31884 6144 31890
rect 6092 31826 6144 31832
rect 4172 31521 4200 31826
rect 7944 31754 7972 33390
rect 9036 32360 9088 32366
rect 9036 32302 9088 32308
rect 5540 31748 5592 31754
rect 5540 31690 5592 31696
rect 7932 31748 7984 31754
rect 7932 31690 7984 31696
rect 4158 31512 4214 31521
rect 4158 31447 4214 31456
rect 5552 31346 5580 31690
rect 9048 31414 9076 32302
rect 9036 31408 9088 31414
rect 9036 31350 9088 31356
rect 4804 31340 4856 31346
rect 4804 31282 4856 31288
rect 5540 31340 5592 31346
rect 5540 31282 5592 31288
rect 4068 31204 4120 31210
rect 4068 31146 4120 31152
rect 3976 31136 4028 31142
rect 3976 31078 4028 31084
rect 3988 30802 4016 31078
rect 4080 30802 4108 31146
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 3976 30796 4028 30802
rect 3976 30738 4028 30744
rect 4068 30796 4120 30802
rect 4068 30738 4120 30744
rect 4816 30394 4844 31282
rect 5816 31272 5868 31278
rect 5816 31214 5868 31220
rect 7472 31272 7524 31278
rect 7472 31214 7524 31220
rect 5828 30870 5856 31214
rect 7484 30938 7512 31214
rect 9048 31210 9076 31350
rect 8300 31204 8352 31210
rect 8300 31146 8352 31152
rect 9036 31204 9088 31210
rect 9036 31146 9088 31152
rect 7472 30932 7524 30938
rect 7472 30874 7524 30880
rect 5816 30864 5868 30870
rect 5816 30806 5868 30812
rect 3884 30388 3936 30394
rect 3884 30330 3936 30336
rect 4804 30388 4856 30394
rect 4804 30330 4856 30336
rect 4712 30320 4764 30326
rect 4712 30262 4764 30268
rect 4068 30252 4120 30258
rect 4068 30194 4120 30200
rect 3882 30152 3938 30161
rect 3882 30087 3938 30096
rect 3792 29844 3844 29850
rect 3792 29786 3844 29792
rect 3896 29102 3924 30087
rect 4080 29646 4108 30194
rect 4620 30048 4672 30054
rect 4620 29990 4672 29996
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4632 29850 4660 29990
rect 4620 29844 4672 29850
rect 4620 29786 4672 29792
rect 4724 29646 4752 30262
rect 8312 30190 8340 31146
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 9324 30598 9352 30670
rect 9496 30660 9548 30666
rect 9496 30602 9548 30608
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 9324 30274 9352 30534
rect 9324 30246 9444 30274
rect 5080 30184 5132 30190
rect 4816 30132 5080 30138
rect 4816 30126 5132 30132
rect 8300 30184 8352 30190
rect 8300 30126 8352 30132
rect 9128 30184 9180 30190
rect 9128 30126 9180 30132
rect 9312 30184 9364 30190
rect 9312 30126 9364 30132
rect 4816 30122 5120 30126
rect 4804 30116 5120 30122
rect 4856 30110 5120 30116
rect 4804 30058 4856 30064
rect 4816 29714 4844 30058
rect 4804 29708 4856 29714
rect 4804 29650 4856 29656
rect 4068 29640 4120 29646
rect 4068 29582 4120 29588
rect 4712 29640 4764 29646
rect 4712 29582 4764 29588
rect 3700 29096 3752 29102
rect 3700 29038 3752 29044
rect 3884 29096 3936 29102
rect 3884 29038 3936 29044
rect 3712 28762 3740 29038
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 3700 28756 3752 28762
rect 3700 28698 3752 28704
rect 4620 28756 4672 28762
rect 4620 28698 4672 28704
rect 4160 28552 4212 28558
rect 4160 28494 4212 28500
rect 4172 27962 4200 28494
rect 4080 27934 4200 27962
rect 4080 27554 4108 27934
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4632 27674 4660 28698
rect 4724 28558 4752 29582
rect 4816 28626 4844 29650
rect 8116 29572 8168 29578
rect 8116 29514 8168 29520
rect 4804 28620 4856 28626
rect 4804 28562 4856 28568
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 4724 28218 4752 28494
rect 4712 28212 4764 28218
rect 4712 28154 4764 28160
rect 4620 27668 4672 27674
rect 4620 27610 4672 27616
rect 4080 27526 4200 27554
rect 3974 27432 4030 27441
rect 4172 27402 4200 27526
rect 4620 27532 4672 27538
rect 4620 27474 4672 27480
rect 3974 27367 4030 27376
rect 4160 27396 4212 27402
rect 3988 26858 4016 27367
rect 4160 27338 4212 27344
rect 4172 26874 4200 27338
rect 3976 26852 4028 26858
rect 3976 26794 4028 26800
rect 4080 26846 4200 26874
rect 4080 26466 4108 26846
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4632 26586 4660 27474
rect 4724 27470 4752 28154
rect 4816 27538 4844 28562
rect 8128 28558 8156 29514
rect 9140 29306 9168 30126
rect 9324 29850 9352 30126
rect 9312 29844 9364 29850
rect 9312 29786 9364 29792
rect 9128 29300 9180 29306
rect 9128 29242 9180 29248
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 8680 28626 8708 28902
rect 8668 28620 8720 28626
rect 8668 28562 8720 28568
rect 5264 28552 5316 28558
rect 5264 28494 5316 28500
rect 8116 28552 8168 28558
rect 8116 28494 8168 28500
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 4804 27532 4856 27538
rect 4804 27474 4856 27480
rect 4712 27464 4764 27470
rect 4712 27406 4764 27412
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 4080 26438 4200 26466
rect 4172 25906 4200 26438
rect 4160 25900 4212 25906
rect 4160 25842 4212 25848
rect 4172 25786 4200 25842
rect 4080 25758 4200 25786
rect 4620 25832 4672 25838
rect 4620 25774 4672 25780
rect 4080 25378 4108 25758
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4080 25350 4200 25378
rect 4632 25362 4660 25774
rect 4724 25362 4752 26726
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4172 25294 4200 25350
rect 4620 25356 4672 25362
rect 4620 25298 4672 25304
rect 4712 25356 4764 25362
rect 4712 25298 4764 25304
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4632 24274 4660 25298
rect 4816 25242 4844 25842
rect 5000 25838 5028 28358
rect 5276 28082 5304 28494
rect 9140 28082 9168 28902
rect 9220 28484 9272 28490
rect 9220 28426 9272 28432
rect 5264 28076 5316 28082
rect 5264 28018 5316 28024
rect 9128 28076 9180 28082
rect 9128 28018 9180 28024
rect 5080 27668 5132 27674
rect 5080 27610 5132 27616
rect 4988 25832 5040 25838
rect 4988 25774 5040 25780
rect 5092 25770 5120 27610
rect 5172 26784 5224 26790
rect 5172 26726 5224 26732
rect 5184 26450 5212 26726
rect 5172 26444 5224 26450
rect 5172 26386 5224 26392
rect 5172 25900 5224 25906
rect 5172 25842 5224 25848
rect 5080 25764 5132 25770
rect 5080 25706 5132 25712
rect 4988 25696 5040 25702
rect 4988 25638 5040 25644
rect 5000 25362 5028 25638
rect 5092 25430 5120 25706
rect 5184 25498 5212 25842
rect 5172 25492 5224 25498
rect 5172 25434 5224 25440
rect 5080 25424 5132 25430
rect 5080 25366 5132 25372
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 4724 25226 4844 25242
rect 4712 25220 4844 25226
rect 4764 25214 4844 25220
rect 4712 25162 4764 25168
rect 4620 24268 4672 24274
rect 4620 24210 4672 24216
rect 4632 24070 4660 24210
rect 4724 24138 4752 25162
rect 4804 25152 4856 25158
rect 4804 25094 4856 25100
rect 4816 24206 4844 25094
rect 5092 24818 5120 25366
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 4908 24274 4936 24550
rect 5092 24410 5120 24754
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 4896 24268 4948 24274
rect 4896 24210 4948 24216
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4712 24132 4764 24138
rect 4712 24074 4764 24080
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4632 23186 4660 24006
rect 4724 23526 4752 24074
rect 5276 23730 5304 28018
rect 9232 27470 9260 28426
rect 9312 28008 9364 28014
rect 9312 27950 9364 27956
rect 9324 27606 9352 27950
rect 9312 27600 9364 27606
rect 9312 27542 9364 27548
rect 9036 27464 9088 27470
rect 9036 27406 9088 27412
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 5540 26852 5592 26858
rect 5540 26794 5592 26800
rect 5552 26518 5580 26794
rect 5540 26512 5592 26518
rect 5540 26454 5592 26460
rect 5356 26308 5408 26314
rect 5356 26250 5408 26256
rect 5368 26042 5396 26250
rect 5448 26240 5500 26246
rect 5448 26182 5500 26188
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 5356 25832 5408 25838
rect 5356 25774 5408 25780
rect 4988 23724 5040 23730
rect 4988 23666 5040 23672
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4172 22778 4200 23054
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 4172 22522 4200 22714
rect 4080 22494 4200 22522
rect 4080 22216 4108 22494
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4080 22188 4292 22216
rect 4172 21690 4200 22188
rect 4264 22030 4292 22188
rect 4632 22098 4660 23122
rect 4724 23050 4752 23462
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4712 23044 4764 23050
rect 4712 22986 4764 22992
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4526 21992 4582 22001
rect 4724 21962 4752 22986
rect 4816 22166 4844 23258
rect 5000 23118 5028 23666
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 4804 22160 4856 22166
rect 4804 22102 4856 22108
rect 4526 21927 4582 21936
rect 4712 21956 4764 21962
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 4172 21332 4200 21626
rect 4540 21593 4568 21927
rect 4712 21898 4764 21904
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4526 21584 4582 21593
rect 4526 21519 4528 21528
rect 4580 21519 4582 21528
rect 4528 21490 4580 21496
rect 4080 21304 4200 21332
rect 4080 21026 4108 21304
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4080 20998 4200 21026
rect 4172 20942 4200 20998
rect 4632 20942 4660 21830
rect 4816 21146 4844 22102
rect 5000 22030 5028 23054
rect 5264 22636 5316 22642
rect 5264 22578 5316 22584
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 5092 21622 5120 22374
rect 5276 22234 5304 22578
rect 5264 22228 5316 22234
rect 5264 22170 5316 22176
rect 5080 21616 5132 21622
rect 5080 21558 5132 21564
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 4988 21480 5040 21486
rect 4988 21422 5040 21428
rect 4804 21140 4856 21146
rect 4804 21082 4856 21088
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4066 20632 4122 20641
rect 4066 20567 4122 20576
rect 4080 20534 4108 20567
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 4172 20466 4200 20742
rect 4632 20466 4660 20878
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4632 18698 4660 20402
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4712 18284 4764 18290
rect 4712 18226 4764 18232
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 3608 17808 3660 17814
rect 3608 17750 3660 17756
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 3160 16114 3188 17138
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3988 16794 4016 17070
rect 4080 16998 4108 17750
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4080 16794 4108 16934
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4066 16552 4122 16561
rect 4066 16487 4122 16496
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3974 15192 4030 15201
rect 3974 15127 4030 15136
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2792 12850 2820 14758
rect 3252 14618 3280 14894
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3896 13841 3924 14758
rect 3988 14550 4016 15127
rect 4080 14890 4108 16487
rect 4632 15978 4660 16594
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4172 15094 4200 15438
rect 4632 15434 4660 15914
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3976 13864 4028 13870
rect 3882 13832 3938 13841
rect 4080 13852 4108 14826
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4028 13824 4108 13852
rect 3976 13806 4028 13812
rect 3882 13767 3938 13776
rect 4080 13410 4108 13824
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4080 13394 4200 13410
rect 4080 13388 4212 13394
rect 4080 13382 4160 13388
rect 4160 13330 4212 13336
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2608 12442 2636 12718
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 1412 11830 1440 12174
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1400 11824 1452 11830
rect 1398 11792 1400 11801
rect 1452 11792 1454 11801
rect 1398 11727 1454 11736
rect 1596 11354 1624 12038
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10441 1440 10610
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 1964 10266 1992 10542
rect 2240 10266 2268 11086
rect 2516 10538 2544 11154
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 9110 1440 9522
rect 1400 9104 1452 9110
rect 1398 9072 1400 9081
rect 1452 9072 1454 9081
rect 1398 9007 1454 9016
rect 2240 8090 2268 10202
rect 2516 10062 2544 10474
rect 2608 10130 2636 11290
rect 2792 11098 2820 12786
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3514 12472 3570 12481
rect 3514 12407 3570 12416
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2700 11082 2820 11098
rect 2688 11076 2820 11082
rect 2740 11070 2820 11076
rect 2688 11018 2740 11024
rect 2976 10674 3004 12038
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7721 1440 7822
rect 1398 7712 1454 7721
rect 1398 7647 1454 7656
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6361 1440 6734
rect 1398 6352 1454 6361
rect 1398 6287 1454 6296
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1412 5001 1440 5170
rect 1398 4992 1454 5001
rect 1398 4927 1454 4936
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1412 3641 1440 4082
rect 2424 4010 2452 9386
rect 2608 8906 2636 9930
rect 2792 9722 2820 9998
rect 2884 9722 2912 10610
rect 3068 10470 3096 10950
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2700 8906 2728 9454
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2516 5914 2544 6258
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2608 5370 2636 8842
rect 2700 6662 2728 8842
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2884 5710 2912 6598
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2412 4004 2464 4010
rect 2412 3946 2464 3952
rect 1398 3632 1454 3641
rect 1398 3567 1454 3576
rect 2884 3534 2912 4014
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 1412 921 1440 3470
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2700 2446 2728 2790
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 1601 1900 2314
rect 2700 2281 2728 2382
rect 2686 2272 2742 2281
rect 2686 2207 2742 2216
rect 1858 1592 1914 1601
rect 1858 1527 1914 1536
rect 1398 912 1454 921
rect 1398 847 1454 856
rect 2792 377 2820 2858
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2976 2514 3004 2790
rect 3068 2650 3096 9318
rect 3344 9178 3372 10610
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3528 8022 3556 12407
rect 3988 10606 4016 12582
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4066 11112 4122 11121
rect 4066 11047 4068 11056
rect 4120 11047 4122 11056
rect 4068 11018 4120 11024
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 10266 4108 10406
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3516 8016 3568 8022
rect 3516 7958 3568 7964
rect 3896 6390 3924 9998
rect 4066 9752 4122 9761
rect 4066 9687 4068 9696
rect 4120 9687 4122 9696
rect 4068 9658 4120 9664
rect 4632 9654 4660 10610
rect 4724 10538 4752 18226
rect 5000 17542 5028 21422
rect 5184 21078 5212 21558
rect 5368 21486 5396 25774
rect 5460 24206 5488 26182
rect 5552 25362 5580 26454
rect 5632 26308 5684 26314
rect 5632 26250 5684 26256
rect 5644 26081 5672 26250
rect 5630 26072 5686 26081
rect 9048 26042 9076 27406
rect 9416 26926 9444 30246
rect 9508 27062 9536 30602
rect 9496 27056 9548 27062
rect 9496 26998 9548 27004
rect 9220 26920 9272 26926
rect 9220 26862 9272 26868
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 5630 26007 5686 26016
rect 9036 26036 9088 26042
rect 9036 25978 9088 25984
rect 9232 25838 9260 26862
rect 9404 26784 9456 26790
rect 9404 26726 9456 26732
rect 9312 26308 9364 26314
rect 9312 26250 9364 26256
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 5540 25356 5592 25362
rect 5540 25298 5592 25304
rect 9128 25220 9180 25226
rect 9128 25162 9180 25168
rect 9140 24954 9168 25162
rect 9128 24948 9180 24954
rect 9128 24890 9180 24896
rect 5816 24608 5868 24614
rect 5816 24550 5868 24556
rect 5448 24200 5500 24206
rect 5448 24142 5500 24148
rect 5460 23730 5488 24142
rect 5448 23724 5500 23730
rect 5448 23666 5500 23672
rect 5828 22438 5856 24550
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6656 23322 6684 24142
rect 6736 23724 6788 23730
rect 6736 23666 6788 23672
rect 6644 23316 6696 23322
rect 6644 23258 6696 23264
rect 6656 22642 6684 23258
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5828 22030 5856 22374
rect 6656 22234 6684 22578
rect 6644 22228 6696 22234
rect 6644 22170 6696 22176
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5448 21548 5500 21554
rect 5448 21490 5500 21496
rect 5356 21480 5408 21486
rect 5356 21422 5408 21428
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 5356 21344 5408 21350
rect 5356 21286 5408 21292
rect 5172 21072 5224 21078
rect 5172 21014 5224 21020
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 5092 20058 5120 20878
rect 5184 20466 5212 21014
rect 5276 21010 5304 21286
rect 5368 21146 5396 21286
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5264 20868 5316 20874
rect 5264 20810 5316 20816
rect 5276 20466 5304 20810
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 5184 19514 5212 20402
rect 5368 20262 5396 21082
rect 5460 20602 5488 21490
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5448 20596 5500 20602
rect 5448 20538 5500 20544
rect 5552 20534 5580 20946
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5552 20330 5580 20470
rect 5540 20324 5592 20330
rect 5540 20266 5592 20272
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5184 18834 5212 19450
rect 6748 19446 6776 23666
rect 7748 23588 7800 23594
rect 7748 23530 7800 23536
rect 7656 22704 7708 22710
rect 7656 22646 7708 22652
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7116 22030 7144 22374
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7116 21865 7144 21966
rect 7392 21894 7420 22170
rect 7668 22030 7696 22646
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7380 21888 7432 21894
rect 7102 21856 7158 21865
rect 7380 21830 7432 21836
rect 7102 21791 7158 21800
rect 7392 21486 7420 21830
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 5092 17882 5120 18702
rect 5184 18222 5212 18770
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 5552 18154 5580 19314
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7024 18766 7052 19110
rect 7300 18970 7328 19790
rect 7392 19310 7420 21422
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7668 20534 7696 21286
rect 7656 20528 7708 20534
rect 7656 20470 7708 20476
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 5080 17604 5132 17610
rect 5184 17592 5212 17750
rect 5132 17564 5212 17592
rect 5080 17546 5132 17552
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5368 14482 5396 18022
rect 5538 17776 5594 17785
rect 5538 17711 5540 17720
rect 5592 17711 5594 17720
rect 5540 17682 5592 17688
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 5460 17338 5488 17546
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5552 17134 5580 17682
rect 5644 17202 5672 18566
rect 5736 18290 5764 18702
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5828 18290 5856 18566
rect 7024 18358 7052 18702
rect 7012 18352 7064 18358
rect 7012 18294 7064 18300
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5816 18284 5868 18290
rect 5816 18226 5868 18232
rect 7300 18086 7328 18906
rect 7760 18834 7788 23530
rect 9232 23186 9260 25774
rect 9324 25770 9352 26250
rect 9416 26042 9444 26726
rect 9404 26036 9456 26042
rect 9404 25978 9456 25984
rect 9508 25922 9536 26998
rect 9588 26988 9640 26994
rect 9588 26930 9640 26936
rect 9600 25974 9628 26930
rect 9416 25906 9536 25922
rect 9588 25968 9640 25974
rect 9588 25910 9640 25916
rect 9404 25900 9536 25906
rect 9456 25894 9536 25900
rect 9404 25842 9456 25848
rect 9312 25764 9364 25770
rect 9312 25706 9364 25712
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 7840 23044 7892 23050
rect 7840 22986 7892 22992
rect 7852 22778 7880 22986
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7852 21146 7880 21830
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 7852 20058 7880 21082
rect 7944 20398 7972 21286
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7392 18222 7420 18770
rect 8220 18698 8248 22714
rect 9416 22642 9444 25842
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 8404 19514 8432 22034
rect 9416 21010 9444 22170
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9600 21554 9628 21966
rect 9588 21548 9640 21554
rect 9508 21508 9588 21536
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 7484 18290 7512 18634
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 6564 16114 6592 18022
rect 7484 17882 7512 18226
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7760 16590 7788 18022
rect 8404 17882 8432 19450
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9140 18290 9168 18702
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9416 17882 9444 20946
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 8404 17746 8432 17818
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9324 17338 9352 17546
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 8404 16726 8432 16934
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 9140 16658 9168 16934
rect 9128 16652 9180 16658
rect 9416 16640 9444 17818
rect 9128 16594 9180 16600
rect 9324 16612 9444 16640
rect 9508 17660 9536 21508
rect 9588 21490 9640 21496
rect 9692 20330 9720 39222
rect 9876 39114 9904 39222
rect 9954 39200 10010 40000
rect 29918 39200 29974 40000
rect 9968 39114 9996 39200
rect 9876 39086 9996 39114
rect 29932 37262 29960 39200
rect 38014 37904 38070 37913
rect 38014 37839 38070 37848
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 38028 37466 38056 37839
rect 38016 37460 38068 37466
rect 38016 37402 38068 37408
rect 29920 37256 29972 37262
rect 29920 37198 29972 37204
rect 37832 37256 37884 37262
rect 37832 37198 37884 37204
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 29932 36922 29960 37198
rect 30196 37120 30248 37126
rect 30196 37062 30248 37068
rect 29920 36916 29972 36922
rect 29920 36858 29972 36864
rect 12348 36780 12400 36786
rect 12348 36722 12400 36728
rect 9772 36236 9824 36242
rect 9772 36178 9824 36184
rect 9784 35630 9812 36178
rect 11980 36100 12032 36106
rect 11980 36042 12032 36048
rect 11520 35692 11572 35698
rect 11520 35634 11572 35640
rect 9772 35624 9824 35630
rect 9772 35566 9824 35572
rect 9784 29102 9812 35566
rect 10140 35488 10192 35494
rect 10140 35430 10192 35436
rect 10152 35222 10180 35430
rect 10140 35216 10192 35222
rect 10140 35158 10192 35164
rect 11532 34746 11560 35634
rect 11888 35624 11940 35630
rect 11888 35566 11940 35572
rect 11796 35012 11848 35018
rect 11796 34954 11848 34960
rect 11520 34740 11572 34746
rect 11520 34682 11572 34688
rect 11808 34610 11836 34954
rect 11796 34604 11848 34610
rect 11796 34546 11848 34552
rect 11900 34542 11928 35566
rect 11992 35154 12020 36042
rect 12360 35290 12388 36722
rect 16396 36712 16448 36718
rect 16396 36654 16448 36660
rect 17500 36712 17552 36718
rect 17500 36654 17552 36660
rect 17960 36712 18012 36718
rect 17960 36654 18012 36660
rect 18052 36712 18104 36718
rect 18052 36654 18104 36660
rect 24584 36712 24636 36718
rect 24584 36654 24636 36660
rect 24768 36712 24820 36718
rect 24768 36654 24820 36660
rect 15200 36644 15252 36650
rect 15200 36586 15252 36592
rect 12624 36576 12676 36582
rect 12624 36518 12676 36524
rect 12532 36372 12584 36378
rect 12532 36314 12584 36320
rect 12440 36236 12492 36242
rect 12440 36178 12492 36184
rect 12452 35698 12480 36178
rect 12440 35692 12492 35698
rect 12440 35634 12492 35640
rect 12544 35494 12572 36314
rect 12636 35766 12664 36518
rect 13820 36236 13872 36242
rect 13820 36178 13872 36184
rect 12808 36168 12860 36174
rect 12808 36110 12860 36116
rect 12716 36032 12768 36038
rect 12716 35974 12768 35980
rect 12624 35760 12676 35766
rect 12624 35702 12676 35708
rect 12532 35488 12584 35494
rect 12532 35430 12584 35436
rect 12348 35284 12400 35290
rect 12348 35226 12400 35232
rect 12544 35222 12572 35430
rect 12532 35216 12584 35222
rect 12532 35158 12584 35164
rect 11980 35148 12032 35154
rect 11980 35090 12032 35096
rect 12440 35080 12492 35086
rect 12440 35022 12492 35028
rect 12452 34746 12480 35022
rect 12440 34740 12492 34746
rect 12440 34682 12492 34688
rect 11980 34604 12032 34610
rect 11980 34546 12032 34552
rect 11888 34536 11940 34542
rect 11888 34478 11940 34484
rect 11152 33856 11204 33862
rect 11152 33798 11204 33804
rect 10508 33516 10560 33522
rect 10508 33458 10560 33464
rect 10520 33318 10548 33458
rect 11164 33454 11192 33798
rect 11152 33448 11204 33454
rect 11152 33390 11204 33396
rect 11060 33380 11112 33386
rect 11060 33322 11112 33328
rect 10508 33312 10560 33318
rect 10508 33254 10560 33260
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9876 30938 9904 31758
rect 9864 30932 9916 30938
rect 9864 30874 9916 30880
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 9784 28626 9812 29038
rect 9772 28620 9824 28626
rect 9772 28562 9824 28568
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 9784 27130 9812 27406
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 10416 26988 10468 26994
rect 10416 26930 10468 26936
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 9784 25702 9812 25978
rect 10048 25968 10100 25974
rect 10048 25910 10100 25916
rect 9956 25900 10008 25906
rect 9956 25842 10008 25848
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 9784 24886 9812 25298
rect 9968 25226 9996 25842
rect 10060 25362 10088 25910
rect 10232 25832 10284 25838
rect 10232 25774 10284 25780
rect 10244 25430 10272 25774
rect 10324 25696 10376 25702
rect 10324 25638 10376 25644
rect 10232 25424 10284 25430
rect 10232 25366 10284 25372
rect 10048 25356 10100 25362
rect 10048 25298 10100 25304
rect 9956 25220 10008 25226
rect 9956 25162 10008 25168
rect 9772 24880 9824 24886
rect 9772 24822 9824 24828
rect 9784 24342 9812 24822
rect 9968 24698 9996 25162
rect 10060 24818 10088 25298
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 10152 24698 10180 24754
rect 10244 24750 10272 25366
rect 9968 24670 10180 24698
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 9772 24336 9824 24342
rect 9772 24278 9824 24284
rect 9864 22568 9916 22574
rect 9864 22510 9916 22516
rect 9876 21894 9904 22510
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9784 21690 9812 21830
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9784 20874 9812 21626
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 9876 19378 9904 21830
rect 9968 21690 9996 24670
rect 10244 21690 10272 24686
rect 10336 24614 10364 25638
rect 10428 25498 10456 26930
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10324 24608 10376 24614
rect 10324 24550 10376 24556
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 9968 21078 9996 21422
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9600 17882 9628 18158
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9692 17870 9904 17898
rect 9692 17814 9720 17870
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9588 17672 9640 17678
rect 9508 17632 9588 17660
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6196 14482 6224 15438
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5184 14006 5212 14350
rect 6380 14346 6408 15846
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7392 15026 7420 15438
rect 7576 15094 7604 16390
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5368 13938 5396 14282
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7024 13462 7052 13806
rect 8220 13462 8248 16458
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8680 13938 8708 15438
rect 9324 14822 9352 16612
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 16250 9444 16458
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9508 15026 9536 17632
rect 9588 17614 9640 17620
rect 9876 17542 9904 17870
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9692 16658 9720 17138
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9600 15162 9628 16050
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 10152 15094 10180 17274
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14618 9352 14758
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 9140 13870 9168 14418
rect 9508 14414 9536 14962
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 8864 13530 8892 13806
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4816 12306 4844 12582
rect 5552 12306 5580 13330
rect 9232 13326 9260 14214
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 7024 12850 7052 13262
rect 8404 12850 8432 13262
rect 9784 12889 9812 14826
rect 10060 14482 10088 14894
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10152 14362 10180 15030
rect 10152 14346 10272 14362
rect 10152 14340 10284 14346
rect 10152 14334 10232 14340
rect 10232 14282 10284 14288
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10152 14006 10180 14214
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10244 13530 10272 14282
rect 10520 13530 10548 33254
rect 11072 33114 11100 33322
rect 11060 33108 11112 33114
rect 11060 33050 11112 33056
rect 11164 32910 11192 33390
rect 11900 32978 11928 34478
rect 11992 33658 12020 34546
rect 12544 34406 12572 35158
rect 12728 35018 12756 35974
rect 12820 35630 12848 36110
rect 13544 36032 13596 36038
rect 13544 35974 13596 35980
rect 12808 35624 12860 35630
rect 12808 35566 12860 35572
rect 12820 35086 12848 35566
rect 12808 35080 12860 35086
rect 12808 35022 12860 35028
rect 12716 35012 12768 35018
rect 12716 34954 12768 34960
rect 12532 34400 12584 34406
rect 12532 34342 12584 34348
rect 12544 34202 12572 34342
rect 12532 34196 12584 34202
rect 12532 34138 12584 34144
rect 12348 33992 12400 33998
rect 12348 33934 12400 33940
rect 11980 33652 12032 33658
rect 11980 33594 12032 33600
rect 12360 33114 12388 33934
rect 12728 33930 12756 34954
rect 12820 34678 12848 35022
rect 13556 35018 13584 35974
rect 13832 35222 13860 36178
rect 14096 36168 14148 36174
rect 14096 36110 14148 36116
rect 13820 35216 13872 35222
rect 13820 35158 13872 35164
rect 14108 35154 14136 36110
rect 15212 35766 15240 36586
rect 16028 36168 16080 36174
rect 16028 36110 16080 36116
rect 15200 35760 15252 35766
rect 15200 35702 15252 35708
rect 14280 35488 14332 35494
rect 14280 35430 14332 35436
rect 14096 35148 14148 35154
rect 14096 35090 14148 35096
rect 13544 35012 13596 35018
rect 13544 34954 13596 34960
rect 12808 34672 12860 34678
rect 12808 34614 12860 34620
rect 12900 34604 12952 34610
rect 12900 34546 12952 34552
rect 13544 34604 13596 34610
rect 13544 34546 13596 34552
rect 12716 33924 12768 33930
rect 12716 33866 12768 33872
rect 12728 33522 12756 33866
rect 12716 33516 12768 33522
rect 12716 33458 12768 33464
rect 12348 33108 12400 33114
rect 12348 33050 12400 33056
rect 11888 32972 11940 32978
rect 11888 32914 11940 32920
rect 11152 32904 11204 32910
rect 11152 32846 11204 32852
rect 12440 32904 12492 32910
rect 12440 32846 12492 32852
rect 11520 32768 11572 32774
rect 11520 32710 11572 32716
rect 11532 31890 11560 32710
rect 12452 32366 12480 32846
rect 12912 32774 12940 34546
rect 13556 33862 13584 34546
rect 13268 33856 13320 33862
rect 13268 33798 13320 33804
rect 13544 33856 13596 33862
rect 13544 33798 13596 33804
rect 12900 32768 12952 32774
rect 12900 32710 12952 32716
rect 12440 32360 12492 32366
rect 12440 32302 12492 32308
rect 11520 31884 11572 31890
rect 11520 31826 11572 31832
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 12440 31816 12492 31822
rect 12440 31758 12492 31764
rect 13084 31816 13136 31822
rect 13084 31758 13136 31764
rect 11348 30802 11376 31758
rect 12072 31408 12124 31414
rect 12072 31350 12124 31356
rect 11980 31136 12032 31142
rect 11980 31078 12032 31084
rect 11336 30796 11388 30802
rect 11336 30738 11388 30744
rect 11152 30728 11204 30734
rect 11152 30670 11204 30676
rect 11164 30258 11192 30670
rect 11152 30252 11204 30258
rect 11152 30194 11204 30200
rect 11992 30054 12020 31078
rect 12084 30326 12112 31350
rect 12176 31346 12296 31362
rect 12164 31340 12296 31346
rect 12216 31334 12296 31340
rect 12164 31282 12216 31288
rect 12164 31204 12216 31210
rect 12164 31146 12216 31152
rect 12072 30320 12124 30326
rect 12072 30262 12124 30268
rect 11980 30048 12032 30054
rect 11980 29990 12032 29996
rect 11992 29714 12020 29990
rect 12084 29850 12112 30262
rect 12176 30190 12204 31146
rect 12268 30258 12296 31334
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 12164 30184 12216 30190
rect 12164 30126 12216 30132
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 12176 29782 12204 30126
rect 12164 29776 12216 29782
rect 12164 29718 12216 29724
rect 11980 29708 12032 29714
rect 11980 29650 12032 29656
rect 12268 28626 12296 30194
rect 12452 30122 12480 31758
rect 12992 31680 13044 31686
rect 12992 31622 13044 31628
rect 13004 31414 13032 31622
rect 12992 31408 13044 31414
rect 12992 31350 13044 31356
rect 13096 31278 13124 31758
rect 13084 31272 13136 31278
rect 13084 31214 13136 31220
rect 12992 30660 13044 30666
rect 12992 30602 13044 30608
rect 12532 30252 12584 30258
rect 12532 30194 12584 30200
rect 12440 30116 12492 30122
rect 12440 30058 12492 30064
rect 12256 28620 12308 28626
rect 12256 28562 12308 28568
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 11440 26450 11468 27406
rect 11888 26852 11940 26858
rect 11888 26794 11940 26800
rect 11612 26784 11664 26790
rect 11612 26726 11664 26732
rect 11624 26450 11652 26726
rect 11900 26586 11928 26794
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 11612 26444 11664 26450
rect 11612 26386 11664 26392
rect 12544 25974 12572 30194
rect 13004 29102 13032 30602
rect 13280 30054 13308 33798
rect 14292 32434 14320 35430
rect 14648 35216 14700 35222
rect 14648 35158 14700 35164
rect 14462 34504 14518 34513
rect 14462 34439 14464 34448
rect 14516 34439 14518 34448
rect 14464 34410 14516 34416
rect 14660 33289 14688 35158
rect 15212 35154 15240 35702
rect 16040 35698 16068 36110
rect 15936 35692 15988 35698
rect 15936 35634 15988 35640
rect 16028 35692 16080 35698
rect 16028 35634 16080 35640
rect 15200 35148 15252 35154
rect 15200 35090 15252 35096
rect 15948 34746 15976 35634
rect 16408 35290 16436 36654
rect 17512 36378 17540 36654
rect 17972 36378 18000 36654
rect 17500 36372 17552 36378
rect 17500 36314 17552 36320
rect 17960 36372 18012 36378
rect 17960 36314 18012 36320
rect 16856 35828 16908 35834
rect 16856 35770 16908 35776
rect 16396 35284 16448 35290
rect 16396 35226 16448 35232
rect 16868 35086 16896 35770
rect 18064 35494 18092 36654
rect 19432 36576 19484 36582
rect 19432 36518 19484 36524
rect 19444 36242 19472 36518
rect 24596 36378 24624 36654
rect 24584 36372 24636 36378
rect 24584 36314 24636 36320
rect 19432 36236 19484 36242
rect 19432 36178 19484 36184
rect 20904 36236 20956 36242
rect 20904 36178 20956 36184
rect 23572 36236 23624 36242
rect 23572 36178 23624 36184
rect 18144 36168 18196 36174
rect 18144 36110 18196 36116
rect 18052 35488 18104 35494
rect 18052 35430 18104 35436
rect 17776 35284 17828 35290
rect 17776 35226 17828 35232
rect 16580 35080 16632 35086
rect 16580 35022 16632 35028
rect 16672 35080 16724 35086
rect 16672 35022 16724 35028
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 15936 34740 15988 34746
rect 15936 34682 15988 34688
rect 16592 34610 16620 35022
rect 15936 34604 15988 34610
rect 15936 34546 15988 34552
rect 16120 34604 16172 34610
rect 16120 34546 16172 34552
rect 16580 34604 16632 34610
rect 16580 34546 16632 34552
rect 15660 33992 15712 33998
rect 15660 33934 15712 33940
rect 14646 33280 14702 33289
rect 14646 33215 14702 33224
rect 14556 32972 14608 32978
rect 14556 32914 14608 32920
rect 14280 32428 14332 32434
rect 14280 32370 14332 32376
rect 14568 30666 14596 32914
rect 14660 32910 14688 33215
rect 14648 32904 14700 32910
rect 14648 32846 14700 32852
rect 15200 32496 15252 32502
rect 15200 32438 15252 32444
rect 14740 31748 14792 31754
rect 14740 31690 14792 31696
rect 14752 30802 14780 31690
rect 15212 30938 15240 32438
rect 15384 31136 15436 31142
rect 15384 31078 15436 31084
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 14740 30796 14792 30802
rect 14740 30738 14792 30744
rect 15108 30796 15160 30802
rect 15108 30738 15160 30744
rect 14556 30660 14608 30666
rect 14556 30602 14608 30608
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 13268 30048 13320 30054
rect 13268 29990 13320 29996
rect 13912 30048 13964 30054
rect 13912 29990 13964 29996
rect 13280 29238 13308 29990
rect 13268 29232 13320 29238
rect 13268 29174 13320 29180
rect 12992 29096 13044 29102
rect 12992 29038 13044 29044
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13004 28014 13032 29038
rect 13832 28626 13860 29038
rect 13820 28620 13872 28626
rect 13820 28562 13872 28568
rect 13084 28552 13136 28558
rect 13924 28506 13952 29990
rect 14108 29646 14136 30194
rect 14568 30054 14596 30602
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14004 29504 14056 29510
rect 14004 29446 14056 29452
rect 13084 28494 13136 28500
rect 12992 28008 13044 28014
rect 12992 27950 13044 27956
rect 13096 27878 13124 28494
rect 13832 28478 13952 28506
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 12532 25968 12584 25974
rect 12532 25910 12584 25916
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 11704 25696 11756 25702
rect 11704 25638 11756 25644
rect 10980 25362 11008 25638
rect 11716 25498 11744 25638
rect 11704 25492 11756 25498
rect 11704 25434 11756 25440
rect 10968 25356 11020 25362
rect 10968 25298 11020 25304
rect 12544 23322 12572 25910
rect 12900 23520 12952 23526
rect 12900 23462 12952 23468
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12912 23118 12940 23462
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 10598 21992 10654 22001
rect 10598 21927 10654 21936
rect 10612 21894 10640 21927
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10704 21010 10732 21626
rect 10888 21554 10916 23054
rect 11348 22098 11376 23054
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 11520 22500 11572 22506
rect 11520 22442 11572 22448
rect 11336 22092 11388 22098
rect 11336 22034 11388 22040
rect 11428 22092 11480 22098
rect 11428 22034 11480 22040
rect 11440 21962 11468 22034
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10888 19242 10916 21490
rect 11348 20602 11376 21898
rect 11532 21554 11560 22442
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 11716 21622 11744 22374
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 12360 21146 12388 22578
rect 12532 22568 12584 22574
rect 12532 22510 12584 22516
rect 12544 22166 12572 22510
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 12452 21418 12480 21558
rect 12544 21486 12572 22102
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12636 21593 12664 22034
rect 12912 21865 12940 23054
rect 12898 21856 12954 21865
rect 12898 21791 12954 21800
rect 12622 21584 12678 21593
rect 12622 21519 12678 21528
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12636 21418 12664 21519
rect 12440 21412 12492 21418
rect 12440 21354 12492 21360
rect 12624 21412 12676 21418
rect 12624 21354 12676 21360
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11808 20466 11836 20742
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11900 19786 11928 21082
rect 12912 20942 12940 21791
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12728 20602 12756 20878
rect 13096 20806 13124 27814
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13280 23322 13308 25842
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 13832 21894 13860 28478
rect 14016 28370 14044 29446
rect 13924 28342 14044 28370
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13556 21690 13584 21830
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12636 19922 12664 20198
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 12348 19780 12400 19786
rect 12348 19722 12400 19728
rect 10876 19236 10928 19242
rect 10876 19178 10928 19184
rect 10888 18766 10916 19178
rect 12360 18970 12388 19722
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 12360 18086 12388 18906
rect 12544 18698 12572 19110
rect 12728 18834 12756 20538
rect 13096 20466 13124 20742
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 13280 20262 13308 20878
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12452 18222 12480 18566
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12440 18080 12492 18086
rect 12544 18068 12572 18634
rect 12728 18290 12756 18770
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12492 18040 12572 18068
rect 12440 18022 12492 18028
rect 12360 17882 12388 18022
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12348 17672 12400 17678
rect 12452 17660 12480 18022
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12544 17678 12572 17750
rect 12636 17746 12664 18158
rect 12728 17746 12756 18226
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12400 17632 12480 17660
rect 12348 17614 12400 17620
rect 12452 17202 12480 17632
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12452 16522 12480 17138
rect 12636 17134 12664 17682
rect 12820 17542 12848 19314
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13188 18358 13216 19110
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 13188 17678 13216 18022
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12912 17202 12940 17546
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12912 17082 12940 17138
rect 13280 17082 13308 20198
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13464 18222 13492 19110
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13372 17202 13400 17614
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13556 17270 13584 17478
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 12636 16658 12664 17070
rect 12912 17054 13032 17082
rect 13280 17054 13400 17082
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12728 16794 12756 16934
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12912 16114 12940 16934
rect 13004 16590 13032 17054
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12544 15026 12572 15438
rect 12728 15094 12756 15846
rect 13096 15570 13124 16390
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 13280 15502 13308 15846
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10612 13938 10640 14418
rect 13004 14006 13032 14894
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 9770 12880 9826 12889
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 8392 12844 8444 12850
rect 9770 12815 9826 12824
rect 8392 12786 8444 12792
rect 9784 12782 9812 12815
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 8588 12306 8616 12718
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 10060 12170 10088 13466
rect 10520 13326 10548 13466
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10520 12986 10548 13262
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 6380 11898 6408 12106
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 10428 11558 10456 12378
rect 10612 12306 10640 13874
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12544 13326 12572 13806
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10612 11694 10640 12242
rect 11440 12238 11468 12922
rect 12912 12850 12940 13194
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 10692 12232 10744 12238
rect 11428 12232 11480 12238
rect 10744 12192 10824 12220
rect 10692 12174 10744 12180
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11762 10732 12038
rect 10796 11762 10824 12192
rect 11428 12174 11480 12180
rect 11440 11898 11468 12174
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10612 11354 10640 11494
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4724 10266 4752 10474
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 5552 9450 5580 9930
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4908 8974 4936 9318
rect 5644 9178 5672 9522
rect 5828 9450 5856 9658
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4066 8392 4122 8401
rect 4066 8327 4068 8336
rect 4120 8327 4122 8336
rect 4068 8298 4120 8304
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4066 7032 4122 7041
rect 4214 7024 4522 7044
rect 4066 6967 4122 6976
rect 4080 6882 4108 6967
rect 4080 6854 4200 6882
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3896 5574 3924 6326
rect 3988 5914 4016 6734
rect 4172 6186 4200 6854
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4632 6322 4660 6734
rect 4816 6390 4844 7142
rect 4908 6662 4936 8910
rect 5184 8362 5212 9046
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5276 8634 5304 8910
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5644 8566 5672 8774
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5184 6866 5212 8298
rect 5276 7410 5304 8366
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4528 5840 4580 5846
rect 4528 5782 4580 5788
rect 4066 5672 4122 5681
rect 4122 5630 4200 5658
rect 4066 5607 4122 5616
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3252 4622 3280 4966
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3160 4146 3188 4422
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3896 3534 3924 5510
rect 4172 5166 4200 5630
rect 4540 5370 4568 5782
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4540 5114 4568 5306
rect 4632 5234 4660 6054
rect 4724 5778 4752 6122
rect 4908 5846 4936 6598
rect 5184 6390 5212 6802
rect 5368 6798 5396 8434
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7546 5488 7686
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 5184 5234 5212 5578
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 4540 5098 4660 5114
rect 4528 5092 4660 5098
rect 4580 5086 4660 5092
rect 4528 5034 4580 5040
rect 4540 5003 4568 5034
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4632 4826 4660 5086
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 5000 4622 5028 4966
rect 5184 4758 5212 5170
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5460 4554 5488 7346
rect 5632 7336 5684 7342
rect 5736 7324 5764 8978
rect 5828 8634 5856 9386
rect 6564 8906 6592 9862
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5684 7296 5764 7324
rect 5632 7278 5684 7284
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6322 5580 6598
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5552 5710 5580 6258
rect 5644 5778 5672 7278
rect 5828 6458 5856 7890
rect 6564 7886 6592 8842
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8634 6960 8774
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 7392 8430 7420 9454
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7954 6684 8230
rect 7576 7954 7604 8366
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 7576 7274 7604 7890
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 8036 6798 8064 11018
rect 10520 10674 10548 11086
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9324 9654 9352 10542
rect 10612 10470 10640 11290
rect 10704 10742 10732 11698
rect 10796 11150 10824 11698
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10152 9926 10180 9998
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9508 9110 9536 9454
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8312 6798 8340 8434
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5828 5710 5856 6394
rect 7944 5710 7972 6598
rect 8036 6458 8064 6734
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8312 6390 8340 6734
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 5552 5234 5580 5646
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5736 4622 5764 5102
rect 5828 4826 5856 5510
rect 6656 5234 6684 5510
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 6656 4690 6684 5170
rect 6748 5166 6776 5578
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 5724 4616 5776 4622
rect 5722 4584 5724 4593
rect 5776 4584 5778 4593
rect 5448 4548 5500 4554
rect 5722 4519 5778 4528
rect 6840 4570 6868 5170
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7288 4616 7340 4622
rect 6840 4564 7288 4570
rect 6840 4558 7340 4564
rect 6840 4542 7328 4558
rect 7392 4554 7420 4626
rect 7380 4548 7432 4554
rect 5448 4490 5500 4496
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 4080 4214 4108 4247
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4448 4146 4476 4422
rect 5460 4282 5488 4490
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 4724 3466 4752 3878
rect 5736 3534 5764 3878
rect 6840 3670 6868 4542
rect 7380 4490 7432 4496
rect 7944 4146 7972 5510
rect 8772 5370 8800 8366
rect 9232 6644 9260 8570
rect 9312 6656 9364 6662
rect 9232 6616 9312 6644
rect 9312 6598 9364 6604
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9048 4690 9076 5102
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 5736 3398 5764 3470
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 3988 2961 4016 3334
rect 5736 3126 5764 3334
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 7760 3058 7788 3878
rect 9324 3194 9352 6598
rect 9508 6361 9536 9046
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10060 7546 10088 7754
rect 10152 7546 10180 9862
rect 10336 9722 10364 9930
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10888 9586 10916 11222
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10980 8974 11008 11494
rect 11900 11354 11928 11630
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 12544 11218 12572 12038
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 11072 10033 11100 10066
rect 11058 10024 11114 10033
rect 11058 9959 11114 9968
rect 11072 9450 11100 9959
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11716 8974 11744 10950
rect 11900 10266 11928 11086
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12176 10742 12204 11018
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12544 10606 12572 11154
rect 12912 10742 12940 12786
rect 13280 12434 13308 15438
rect 13372 15434 13400 17054
rect 13832 15910 13860 21490
rect 13924 21350 13952 28342
rect 14108 27146 14136 29582
rect 15120 29170 15148 30738
rect 15396 30734 15424 31078
rect 15384 30728 15436 30734
rect 15384 30670 15436 30676
rect 15672 30326 15700 33934
rect 15948 32910 15976 34546
rect 16132 34406 16160 34546
rect 16684 34542 16712 35022
rect 16868 34746 16896 35022
rect 17316 35012 17368 35018
rect 17316 34954 17368 34960
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 16672 34536 16724 34542
rect 16672 34478 16724 34484
rect 16948 34536 17000 34542
rect 16948 34478 17000 34484
rect 16120 34400 16172 34406
rect 16120 34342 16172 34348
rect 16212 34060 16264 34066
rect 16212 34002 16264 34008
rect 16224 33658 16252 34002
rect 16672 33856 16724 33862
rect 16672 33798 16724 33804
rect 16212 33652 16264 33658
rect 16212 33594 16264 33600
rect 15936 32904 15988 32910
rect 15936 32846 15988 32852
rect 15660 30320 15712 30326
rect 15660 30262 15712 30268
rect 15672 29714 15700 30262
rect 15660 29708 15712 29714
rect 15660 29650 15712 29656
rect 15844 29640 15896 29646
rect 15844 29582 15896 29588
rect 15292 29504 15344 29510
rect 15292 29446 15344 29452
rect 15304 29170 15332 29446
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 15292 29164 15344 29170
rect 15292 29106 15344 29112
rect 15856 28966 15884 29582
rect 15936 29028 15988 29034
rect 15936 28970 15988 28976
rect 14832 28960 14884 28966
rect 14832 28902 14884 28908
rect 15844 28960 15896 28966
rect 15844 28902 15896 28908
rect 14844 28626 14872 28902
rect 15856 28762 15884 28902
rect 15844 28756 15896 28762
rect 15844 28698 15896 28704
rect 14832 28620 14884 28626
rect 14832 28562 14884 28568
rect 14924 28076 14976 28082
rect 14924 28018 14976 28024
rect 14280 27872 14332 27878
rect 14280 27814 14332 27820
rect 14464 27872 14516 27878
rect 14464 27814 14516 27820
rect 14292 27538 14320 27814
rect 14280 27532 14332 27538
rect 14280 27474 14332 27480
rect 14016 27118 14136 27146
rect 14016 26042 14044 27118
rect 14476 27062 14504 27814
rect 14464 27056 14516 27062
rect 14464 26998 14516 27004
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14292 26586 14320 26862
rect 14936 26586 14964 28018
rect 15856 27946 15884 28698
rect 15948 28558 15976 28970
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 15948 28082 15976 28494
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 15844 27940 15896 27946
rect 15844 27882 15896 27888
rect 15384 27872 15436 27878
rect 15384 27814 15436 27820
rect 15660 27872 15712 27878
rect 15660 27814 15712 27820
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14924 26580 14976 26586
rect 14924 26522 14976 26528
rect 15396 26450 15424 27814
rect 15672 27538 15700 27814
rect 15660 27532 15712 27538
rect 15660 27474 15712 27480
rect 15752 27532 15804 27538
rect 15752 27474 15804 27480
rect 15764 26926 15792 27474
rect 15948 27470 15976 28018
rect 15936 27464 15988 27470
rect 15936 27406 15988 27412
rect 15752 26920 15804 26926
rect 15752 26862 15804 26868
rect 15384 26444 15436 26450
rect 15384 26386 15436 26392
rect 15948 26382 15976 27406
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 14004 26036 14056 26042
rect 14004 25978 14056 25984
rect 14108 25974 14136 26318
rect 14096 25968 14148 25974
rect 14096 25910 14148 25916
rect 15292 25832 15344 25838
rect 15292 25774 15344 25780
rect 15304 24750 15332 25774
rect 15292 24744 15344 24750
rect 15292 24686 15344 24692
rect 15660 24744 15712 24750
rect 15660 24686 15712 24692
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15672 24274 15700 24686
rect 15856 24410 15884 24686
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 15660 24268 15712 24274
rect 15660 24210 15712 24216
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 15304 23186 15332 23462
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 14016 22438 14044 23054
rect 15292 23044 15344 23050
rect 15292 22986 15344 22992
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 14924 22432 14976 22438
rect 14924 22374 14976 22380
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 14016 21554 14044 22374
rect 14936 22098 14964 22374
rect 15212 22098 15240 22374
rect 15304 22166 15332 22986
rect 16040 22642 16068 23462
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 15200 22092 15252 22098
rect 16224 22094 16252 33594
rect 16684 33522 16712 33798
rect 16672 33516 16724 33522
rect 16672 33458 16724 33464
rect 16960 33454 16988 34478
rect 17132 34400 17184 34406
rect 17132 34342 17184 34348
rect 17144 34134 17172 34342
rect 17132 34128 17184 34134
rect 17132 34070 17184 34076
rect 17224 33992 17276 33998
rect 17224 33934 17276 33940
rect 17236 33522 17264 33934
rect 17328 33930 17356 34954
rect 17682 34640 17738 34649
rect 17682 34575 17738 34584
rect 17696 34542 17724 34575
rect 17684 34536 17736 34542
rect 17684 34478 17736 34484
rect 17788 34406 17816 35226
rect 17960 35148 18012 35154
rect 17960 35090 18012 35096
rect 17868 35080 17920 35086
rect 17868 35022 17920 35028
rect 17880 34610 17908 35022
rect 17868 34604 17920 34610
rect 17868 34546 17920 34552
rect 17776 34400 17828 34406
rect 17776 34342 17828 34348
rect 17972 34066 18000 35090
rect 18052 34740 18104 34746
rect 18156 34728 18184 36110
rect 20916 36038 20944 36178
rect 21732 36168 21784 36174
rect 21732 36110 21784 36116
rect 19432 36032 19484 36038
rect 19432 35974 19484 35980
rect 20904 36032 20956 36038
rect 20904 35974 20956 35980
rect 19444 35834 19472 35974
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 20916 35766 20944 35974
rect 20904 35760 20956 35766
rect 20904 35702 20956 35708
rect 21744 35698 21772 36110
rect 21916 36100 21968 36106
rect 21916 36042 21968 36048
rect 21928 35834 21956 36042
rect 23584 35894 23612 36178
rect 24308 36168 24360 36174
rect 24308 36110 24360 36116
rect 23584 35866 23796 35894
rect 21916 35828 21968 35834
rect 21916 35770 21968 35776
rect 18972 35692 19024 35698
rect 18972 35634 19024 35640
rect 20628 35692 20680 35698
rect 20628 35634 20680 35640
rect 21732 35692 21784 35698
rect 21732 35634 21784 35640
rect 18236 35624 18288 35630
rect 18236 35566 18288 35572
rect 18248 34950 18276 35566
rect 18328 35488 18380 35494
rect 18328 35430 18380 35436
rect 18236 34944 18288 34950
rect 18236 34886 18288 34892
rect 18104 34700 18184 34728
rect 18052 34682 18104 34688
rect 18052 34536 18104 34542
rect 18144 34536 18196 34542
rect 18104 34496 18144 34524
rect 18052 34478 18104 34484
rect 18144 34478 18196 34484
rect 17960 34060 18012 34066
rect 17960 34002 18012 34008
rect 17316 33924 17368 33930
rect 17316 33866 17368 33872
rect 17224 33516 17276 33522
rect 17224 33458 17276 33464
rect 16948 33448 17000 33454
rect 16948 33390 17000 33396
rect 17236 33114 17264 33458
rect 17972 33289 18000 34002
rect 17958 33280 18014 33289
rect 17958 33215 18014 33224
rect 17224 33108 17276 33114
rect 17224 33050 17276 33056
rect 17960 32972 18012 32978
rect 17960 32914 18012 32920
rect 17040 32768 17092 32774
rect 17040 32710 17092 32716
rect 16396 31952 16448 31958
rect 16396 31894 16448 31900
rect 16408 31754 16436 31894
rect 16580 31884 16632 31890
rect 16580 31826 16632 31832
rect 16592 31754 16620 31826
rect 16304 31748 16356 31754
rect 16408 31726 16620 31754
rect 16304 31690 16356 31696
rect 16316 30802 16344 31690
rect 16592 31414 16620 31726
rect 17052 31414 17080 32710
rect 17972 31414 18000 32914
rect 18064 32434 18092 34478
rect 18144 33448 18196 33454
rect 18144 33390 18196 33396
rect 18156 32910 18184 33390
rect 18144 32904 18196 32910
rect 18144 32846 18196 32852
rect 18052 32428 18104 32434
rect 18052 32370 18104 32376
rect 16580 31408 16632 31414
rect 16580 31350 16632 31356
rect 17040 31408 17092 31414
rect 17040 31350 17092 31356
rect 17960 31408 18012 31414
rect 17960 31350 18012 31356
rect 16304 30796 16356 30802
rect 16304 30738 16356 30744
rect 16672 29096 16724 29102
rect 16672 29038 16724 29044
rect 16580 28620 16632 28626
rect 16580 28562 16632 28568
rect 16592 28218 16620 28562
rect 16580 28212 16632 28218
rect 16580 28154 16632 28160
rect 16488 27940 16540 27946
rect 16488 27882 16540 27888
rect 16500 27674 16528 27882
rect 16488 27668 16540 27674
rect 16488 27610 16540 27616
rect 16500 26586 16528 27610
rect 16592 27538 16620 28154
rect 16580 27532 16632 27538
rect 16580 27474 16632 27480
rect 16488 26580 16540 26586
rect 16488 26522 16540 26528
rect 16684 26382 16712 29038
rect 17052 28490 17080 31350
rect 17776 30864 17828 30870
rect 17776 30806 17828 30812
rect 17788 30054 17816 30806
rect 18052 30660 18104 30666
rect 18052 30602 18104 30608
rect 18064 30258 18092 30602
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 17776 30048 17828 30054
rect 17776 29990 17828 29996
rect 17788 29714 17816 29990
rect 18156 29866 18184 32846
rect 18248 31958 18276 34886
rect 18340 32978 18368 35430
rect 18788 35080 18840 35086
rect 18788 35022 18840 35028
rect 18602 34640 18658 34649
rect 18800 34610 18828 35022
rect 18984 34746 19012 35634
rect 20640 35290 20668 35634
rect 23768 35630 23796 35866
rect 23112 35624 23164 35630
rect 23112 35566 23164 35572
rect 23296 35624 23348 35630
rect 23296 35566 23348 35572
rect 23756 35624 23808 35630
rect 23756 35566 23808 35572
rect 21916 35488 21968 35494
rect 21916 35430 21968 35436
rect 20628 35284 20680 35290
rect 20628 35226 20680 35232
rect 21928 35154 21956 35430
rect 21916 35148 21968 35154
rect 21916 35090 21968 35096
rect 21180 35012 21232 35018
rect 21180 34954 21232 34960
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 21192 34746 21220 34954
rect 18972 34740 19024 34746
rect 18972 34682 19024 34688
rect 21180 34740 21232 34746
rect 21180 34682 21232 34688
rect 18602 34575 18658 34584
rect 18788 34604 18840 34610
rect 18616 34542 18644 34575
rect 18788 34546 18840 34552
rect 20168 34604 20220 34610
rect 20168 34546 20220 34552
rect 18604 34536 18656 34542
rect 18418 34504 18474 34513
rect 18656 34496 18736 34524
rect 18604 34478 18656 34484
rect 18418 34439 18420 34448
rect 18472 34439 18474 34448
rect 18420 34410 18472 34416
rect 18604 34196 18656 34202
rect 18604 34138 18656 34144
rect 18616 33318 18644 34138
rect 18708 34048 18736 34496
rect 19340 34400 19392 34406
rect 19340 34342 19392 34348
rect 18788 34060 18840 34066
rect 18708 34020 18788 34048
rect 18708 33522 18736 34020
rect 18788 34002 18840 34008
rect 19352 33930 19380 34342
rect 19340 33924 19392 33930
rect 19340 33866 19392 33872
rect 19352 33522 19380 33866
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 20180 33658 20208 34546
rect 21824 34536 21876 34542
rect 21824 34478 21876 34484
rect 22008 34536 22060 34542
rect 22008 34478 22060 34484
rect 21836 34202 21864 34478
rect 21824 34196 21876 34202
rect 21824 34138 21876 34144
rect 22020 34134 22048 34478
rect 23124 34202 23152 35566
rect 23112 34196 23164 34202
rect 23112 34138 23164 34144
rect 22008 34128 22060 34134
rect 22008 34070 22060 34076
rect 20168 33652 20220 33658
rect 20168 33594 20220 33600
rect 18696 33516 18748 33522
rect 18696 33458 18748 33464
rect 19340 33516 19392 33522
rect 19340 33458 19392 33464
rect 18420 33312 18472 33318
rect 18420 33254 18472 33260
rect 18604 33312 18656 33318
rect 18604 33254 18656 33260
rect 18328 32972 18380 32978
rect 18328 32914 18380 32920
rect 18236 31952 18288 31958
rect 18236 31894 18288 31900
rect 18432 31822 18460 33254
rect 18708 33114 18736 33458
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 18696 33108 18748 33114
rect 18696 33050 18748 33056
rect 19996 32774 20024 33254
rect 23308 32978 23336 35566
rect 23768 35154 23796 35566
rect 23756 35148 23808 35154
rect 23756 35090 23808 35096
rect 23480 35080 23532 35086
rect 23480 35022 23532 35028
rect 23492 33862 23520 35022
rect 24320 34610 24348 36110
rect 24780 35154 24808 36654
rect 27620 36644 27672 36650
rect 27620 36586 27672 36592
rect 26608 36576 26660 36582
rect 26608 36518 26660 36524
rect 26620 36242 26648 36518
rect 27632 36242 27660 36586
rect 26608 36236 26660 36242
rect 26608 36178 26660 36184
rect 27620 36236 27672 36242
rect 27620 36178 27672 36184
rect 26148 36168 26200 36174
rect 26148 36110 26200 36116
rect 25596 36032 25648 36038
rect 25596 35974 25648 35980
rect 24584 35148 24636 35154
rect 24584 35090 24636 35096
rect 24768 35148 24820 35154
rect 24768 35090 24820 35096
rect 24308 34604 24360 34610
rect 24308 34546 24360 34552
rect 24596 34542 24624 35090
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 24584 34536 24636 34542
rect 24584 34478 24636 34484
rect 23664 34468 23716 34474
rect 23664 34410 23716 34416
rect 23480 33856 23532 33862
rect 23480 33798 23532 33804
rect 23572 33856 23624 33862
rect 23572 33798 23624 33804
rect 23296 32972 23348 32978
rect 23296 32914 23348 32920
rect 22560 32904 22612 32910
rect 22560 32846 22612 32852
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 18788 32428 18840 32434
rect 18788 32370 18840 32376
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 18420 31816 18472 31822
rect 18420 31758 18472 31764
rect 18064 29838 18184 29866
rect 17776 29708 17828 29714
rect 17776 29650 17828 29656
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17040 28484 17092 28490
rect 17040 28426 17092 28432
rect 16856 28416 16908 28422
rect 16856 28358 16908 28364
rect 16868 28082 16896 28358
rect 17052 28150 17080 28426
rect 17040 28144 17092 28150
rect 17040 28086 17092 28092
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 17052 27402 17080 28086
rect 17040 27396 17092 27402
rect 17040 27338 17092 27344
rect 16396 26376 16448 26382
rect 16396 26318 16448 26324
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16408 24274 16436 26318
rect 16684 24818 16712 26318
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16684 24138 16712 24754
rect 17132 24404 17184 24410
rect 17132 24346 17184 24352
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16868 23866 16896 24142
rect 16856 23860 16908 23866
rect 16856 23802 16908 23808
rect 16868 23730 16896 23802
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16960 23662 16988 24210
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 16684 22506 16712 22986
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16868 22642 16896 22918
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16672 22500 16724 22506
rect 16672 22442 16724 22448
rect 15200 22034 15252 22040
rect 16132 22066 16252 22094
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13924 19990 13952 21286
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 13912 19984 13964 19990
rect 13912 19926 13964 19932
rect 14936 19922 14964 20334
rect 14924 19916 14976 19922
rect 14924 19858 14976 19864
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14476 19378 14504 19790
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14660 18970 14688 19722
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 15120 17864 15148 21830
rect 15200 17876 15252 17882
rect 15120 17836 15200 17864
rect 15200 17818 15252 17824
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15120 16522 15148 17070
rect 15108 16516 15160 16522
rect 15108 16458 15160 16464
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13096 12406 13308 12434
rect 13096 11150 13124 12406
rect 13372 12102 13400 15370
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14660 12850 14688 13806
rect 14844 13530 14872 13806
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 15212 13326 15240 17818
rect 15936 16720 15988 16726
rect 15936 16662 15988 16668
rect 15948 16114 15976 16662
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15948 15502 15976 16050
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15212 12986 15240 13262
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 15108 12436 15160 12442
rect 15212 12434 15240 12922
rect 15160 12406 15240 12434
rect 15108 12378 15160 12384
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 11762 13400 12038
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 12084 9586 12112 10406
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6798 9720 7142
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9494 6352 9550 6361
rect 9494 6287 9550 6296
rect 10244 6254 10272 6802
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10244 5710 10272 6190
rect 10980 6186 11008 8366
rect 11164 7954 11192 8774
rect 11808 8566 11836 9454
rect 12728 9042 12756 10406
rect 13096 9926 13124 11086
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13188 10674 13216 10950
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8566 12204 8774
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11440 7546 11468 7890
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11992 6662 12020 8366
rect 12636 7478 12664 8910
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12440 7336 12492 7342
rect 12492 7296 12572 7324
rect 12440 7278 12492 7284
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10980 5914 11008 6122
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10336 5166 10364 5510
rect 12544 5234 12572 7296
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9784 3670 9812 5034
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10506 4856 10562 4865
rect 10506 4791 10562 4800
rect 10520 4622 10548 4791
rect 10704 4622 10732 4966
rect 10796 4690 10824 5170
rect 12438 4856 12494 4865
rect 12438 4791 12494 4800
rect 12452 4758 12480 4791
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10796 4214 10824 4490
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 11532 4146 11560 4422
rect 11900 4282 11928 4558
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11624 4185 11652 4218
rect 11610 4176 11666 4185
rect 11520 4140 11572 4146
rect 11610 4111 11666 4120
rect 11520 4082 11572 4088
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 10888 3534 10916 3878
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 11256 3466 11284 3674
rect 13096 3602 13124 9862
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 11716 3126 11744 3334
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 3974 2952 4030 2961
rect 3974 2887 4030 2896
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 13372 2378 13400 11698
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13832 11150 13860 11630
rect 14016 11218 14044 11766
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13832 10606 13860 11086
rect 14016 10674 14044 11154
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13832 10062 13860 10542
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13740 6458 13768 8502
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 14200 4593 14228 7414
rect 14568 6458 14596 7822
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14292 5710 14320 6054
rect 14384 5710 14412 6326
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14476 5642 14504 6122
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14292 4622 14320 5510
rect 14476 4826 14504 5578
rect 14568 5370 14596 6394
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14568 4622 14596 5306
rect 14660 4690 14688 12106
rect 15108 11280 15160 11286
rect 15108 11222 15160 11228
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 15028 10062 15056 10678
rect 15120 10470 15148 11222
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 10674 15240 10950
rect 15304 10810 15332 15302
rect 16132 14074 16160 22066
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16316 20466 16344 20878
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16960 19922 16988 20878
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16776 19378 16804 19790
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 16316 17678 16344 17818
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16224 15638 16252 16390
rect 16868 15910 16896 17818
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16960 15706 16988 16050
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16224 15366 16252 15574
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16132 13954 16160 14010
rect 16040 13926 16160 13954
rect 16040 13394 16068 13926
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 15396 11354 15424 11562
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15948 11286 15976 11494
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 16040 10810 16068 13330
rect 16776 12918 16804 13466
rect 16868 13190 16896 15302
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 14074 16988 14894
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16868 11762 16896 13126
rect 17052 12986 17080 23598
rect 17144 23526 17172 24346
rect 17236 23866 17264 29106
rect 17684 27532 17736 27538
rect 17684 27474 17736 27480
rect 17696 26926 17724 27474
rect 18064 26994 18092 29838
rect 18144 29776 18196 29782
rect 18144 29718 18196 29724
rect 18156 29306 18184 29718
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18524 26994 18552 27406
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 18512 26988 18564 26994
rect 18512 26930 18564 26936
rect 17684 26920 17736 26926
rect 17684 26862 17736 26868
rect 17316 24132 17368 24138
rect 17316 24074 17368 24080
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 17328 23730 17356 24074
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 17696 23186 17724 26862
rect 18064 26586 18092 26930
rect 18616 26874 18644 31962
rect 18800 30122 18828 32370
rect 19340 32360 19392 32366
rect 19340 32302 19392 32308
rect 18880 32224 18932 32230
rect 18880 32166 18932 32172
rect 18892 31414 18920 32166
rect 18880 31408 18932 31414
rect 18880 31350 18932 31356
rect 19352 31278 19380 32302
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19340 31272 19392 31278
rect 19340 31214 19392 31220
rect 19352 30818 19380 31214
rect 19260 30790 19380 30818
rect 19996 30802 20024 32710
rect 22100 32360 22152 32366
rect 22100 32302 22152 32308
rect 20076 31816 20128 31822
rect 20076 31758 20128 31764
rect 20088 31346 20116 31758
rect 20076 31340 20128 31346
rect 20076 31282 20128 31288
rect 21548 31340 21600 31346
rect 21548 31282 21600 31288
rect 19984 30796 20036 30802
rect 19260 30598 19288 30790
rect 19984 30738 20036 30744
rect 19524 30728 19576 30734
rect 19444 30688 19524 30716
rect 19340 30660 19392 30666
rect 19340 30602 19392 30608
rect 19248 30592 19300 30598
rect 19248 30534 19300 30540
rect 19352 30326 19380 30602
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19340 30184 19392 30190
rect 19444 30172 19472 30688
rect 19524 30670 19576 30676
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19996 30394 20024 30738
rect 20904 30728 20956 30734
rect 20904 30670 20956 30676
rect 20260 30660 20312 30666
rect 20260 30602 20312 30608
rect 20076 30592 20128 30598
rect 20076 30534 20128 30540
rect 19984 30388 20036 30394
rect 19984 30330 20036 30336
rect 19392 30144 19472 30172
rect 19340 30126 19392 30132
rect 18788 30116 18840 30122
rect 18788 30058 18840 30064
rect 19352 29170 19380 30126
rect 20088 30054 20116 30534
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 18880 29096 18932 29102
rect 18880 29038 18932 29044
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 18892 28014 18920 29038
rect 18880 28008 18932 28014
rect 18880 27950 18932 27956
rect 18696 27328 18748 27334
rect 18696 27270 18748 27276
rect 18708 27062 18736 27270
rect 18696 27056 18748 27062
rect 18696 26998 18748 27004
rect 18616 26846 18736 26874
rect 18052 26580 18104 26586
rect 18052 26522 18104 26528
rect 18420 26580 18472 26586
rect 18420 26522 18472 26528
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 18064 22574 18092 23598
rect 18156 23322 18184 24346
rect 18236 23792 18288 23798
rect 18236 23734 18288 23740
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 18052 22568 18104 22574
rect 18052 22510 18104 22516
rect 18156 22438 18184 23258
rect 18248 23118 18276 23734
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 18248 22710 18276 23054
rect 18236 22704 18288 22710
rect 18236 22646 18288 22652
rect 18236 22568 18288 22574
rect 18236 22510 18288 22516
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 18144 22432 18196 22438
rect 18144 22374 18196 22380
rect 17696 21554 17724 22374
rect 18052 22092 18104 22098
rect 18052 22034 18104 22040
rect 18064 21962 18092 22034
rect 18052 21956 18104 21962
rect 18052 21898 18104 21904
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17420 20534 17448 21422
rect 17408 20528 17460 20534
rect 17408 20470 17460 20476
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17604 18290 17632 18702
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17972 18222 18000 19858
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 18064 18068 18092 21898
rect 18248 21894 18276 22510
rect 18432 22098 18460 26522
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18524 23594 18552 24142
rect 18512 23588 18564 23594
rect 18512 23530 18564 23536
rect 18524 23118 18552 23530
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18524 22642 18552 23054
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 18420 22092 18472 22098
rect 18420 22034 18472 22040
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18248 21622 18276 21830
rect 18236 21616 18288 21622
rect 18236 21558 18288 21564
rect 18616 21010 18644 22374
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18156 18834 18184 19110
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 17972 18040 18092 18068
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17328 14074 17356 14282
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17236 13530 17264 13874
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16684 11354 16712 11630
rect 16868 11354 16896 11698
rect 17144 11694 17172 12786
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15212 10554 15240 10610
rect 15212 10526 15332 10554
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15120 10266 15148 10406
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15304 10062 15332 10526
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15488 9586 15516 10406
rect 16040 10266 16068 10746
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15856 9586 15884 9862
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15304 7954 15332 9318
rect 15580 9042 15608 9318
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15396 7426 15424 8910
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15304 7410 15424 7426
rect 15292 7404 15424 7410
rect 15344 7398 15424 7404
rect 15566 7440 15622 7449
rect 15622 7398 15700 7426
rect 15566 7375 15568 7384
rect 15292 7346 15344 7352
rect 15620 7375 15622 7384
rect 15568 7346 15620 7352
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14936 6458 14964 7142
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15212 5098 15240 5510
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 15304 5030 15332 7346
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15580 6866 15608 7210
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15672 6798 15700 7398
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 14280 4616 14332 4622
rect 14186 4584 14242 4593
rect 14280 4558 14332 4564
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14186 4519 14242 4528
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13832 4146 13860 4422
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13464 3058 13492 3878
rect 14568 3194 14596 4558
rect 14660 4282 14688 4626
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 15212 4078 15240 4626
rect 15304 4214 15332 4966
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15396 4146 15424 6598
rect 15672 6458 15700 6734
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15580 5658 15608 6190
rect 15672 5778 15700 6394
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15580 5630 15700 5658
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15488 4282 15516 5306
rect 15672 5166 15700 5630
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15672 4010 15700 5102
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15764 3738 15792 7890
rect 16592 7313 16620 8978
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16578 7304 16634 7313
rect 16578 7239 16634 7248
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16500 6254 16528 6802
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15856 4826 15884 5170
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15948 4690 15976 4966
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 16396 4548 16448 4554
rect 16396 4490 16448 4496
rect 16408 3738 16436 4490
rect 16592 4185 16620 7239
rect 16578 4176 16634 4185
rect 16578 4111 16634 4120
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 16684 3126 16712 8298
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16868 6798 16896 7754
rect 17144 7410 17172 7890
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16868 4554 16896 6734
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 17052 5234 17080 6122
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17144 4758 17172 7346
rect 17236 6798 17264 10474
rect 17420 9518 17448 15846
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17512 13462 17540 13874
rect 17500 13456 17552 13462
rect 17500 13398 17552 13404
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17604 11150 17632 11290
rect 17788 11234 17816 17478
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17880 15366 17908 16050
rect 17972 15978 18000 18040
rect 18156 17814 18184 18770
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18144 17808 18196 17814
rect 18144 17750 18196 17756
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18156 16590 18184 17206
rect 18248 17134 18276 18158
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18432 16998 18460 18702
rect 18708 18358 18736 26846
rect 18892 19446 18920 27950
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19260 24410 19288 25230
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19260 23798 19288 24006
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18984 23594 19012 23666
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 18972 23588 19024 23594
rect 18972 23530 19024 23536
rect 19168 23526 19196 23598
rect 19156 23520 19208 23526
rect 19156 23462 19208 23468
rect 19260 23322 19288 23598
rect 19248 23316 19300 23322
rect 19248 23258 19300 23264
rect 18972 23044 19024 23050
rect 18972 22986 19024 22992
rect 18984 22574 19012 22986
rect 18972 22568 19024 22574
rect 18972 22510 19024 22516
rect 19352 20262 19380 27406
rect 19444 27402 19472 29038
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19432 26920 19484 26926
rect 19432 26862 19484 26868
rect 19444 26450 19472 26862
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19432 26308 19484 26314
rect 19432 26250 19484 26256
rect 19444 25498 19472 26250
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19432 25492 19484 25498
rect 19432 25434 19484 25440
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19996 23254 20024 24142
rect 19984 23248 20036 23254
rect 19984 23190 20036 23196
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19444 22642 19472 22918
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19444 21622 19472 22374
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19432 21616 19484 21622
rect 19432 21558 19484 21564
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 19720 21146 19748 21422
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19628 19854 19656 20266
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18892 18766 18920 19382
rect 19892 19372 19944 19378
rect 19996 19360 20024 20198
rect 19944 19332 20024 19360
rect 19892 19314 19944 19320
rect 19904 18834 19932 19314
rect 20088 18970 20116 29990
rect 20272 29306 20300 30602
rect 20536 30388 20588 30394
rect 20536 30330 20588 30336
rect 20444 30252 20496 30258
rect 20444 30194 20496 30200
rect 20352 30116 20404 30122
rect 20352 30058 20404 30064
rect 20364 29714 20392 30058
rect 20352 29708 20404 29714
rect 20352 29650 20404 29656
rect 20260 29300 20312 29306
rect 20260 29242 20312 29248
rect 20260 27396 20312 27402
rect 20260 27338 20312 27344
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 23730 20208 24754
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 20180 23118 20208 23666
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 20076 18964 20128 18970
rect 20128 18924 20208 18952
rect 20076 18906 20128 18912
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18524 17134 18552 17682
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18340 16658 18368 16934
rect 18432 16726 18460 16934
rect 18420 16720 18472 16726
rect 18420 16662 18472 16668
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18340 16046 18368 16594
rect 18524 16590 18552 17070
rect 18616 16794 18644 17818
rect 18788 17808 18840 17814
rect 18788 17750 18840 17756
rect 18800 17338 18828 17750
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18984 16658 19012 18702
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19352 17626 19380 18566
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 20088 17746 20116 18022
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 19260 17610 19380 17626
rect 19248 17604 19380 17610
rect 19300 17598 19380 17604
rect 19248 17546 19300 17552
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17972 15570 18000 15914
rect 18340 15706 18368 15982
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17880 11898 17908 12718
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17788 11206 17908 11234
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17604 10674 17632 11086
rect 17880 10674 17908 11206
rect 18064 10742 18092 15642
rect 18616 14550 18644 16390
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19444 14958 19472 15438
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19996 15162 20024 16594
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19352 14618 19380 14758
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 18604 14544 18656 14550
rect 18604 14486 18656 14492
rect 19248 14340 19300 14346
rect 19248 14282 19300 14288
rect 19260 14074 19288 14282
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19352 13530 19380 14554
rect 19444 14482 19472 14894
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18248 12306 18276 13262
rect 19352 12986 19380 13466
rect 19444 13394 19472 14418
rect 19536 14346 19564 14826
rect 19628 14414 19656 14962
rect 19812 14618 19840 14962
rect 19800 14612 19852 14618
rect 19800 14554 19852 14560
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19524 14340 19576 14346
rect 19524 14282 19576 14288
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19996 13326 20024 14350
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 20180 12986 20208 18924
rect 20272 17882 20300 27338
rect 20364 24750 20392 29650
rect 20456 29646 20484 30194
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20352 24744 20404 24750
rect 20352 24686 20404 24692
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20364 23730 20392 24142
rect 20352 23724 20404 23730
rect 20352 23666 20404 23672
rect 20364 23322 20392 23666
rect 20352 23316 20404 23322
rect 20352 23258 20404 23264
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20364 22098 20392 22374
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20444 22092 20496 22098
rect 20444 22034 20496 22040
rect 20456 21486 20484 22034
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20272 16658 20300 17546
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20548 14890 20576 30330
rect 20916 29646 20944 30670
rect 21560 30666 21588 31282
rect 21916 31272 21968 31278
rect 21916 31214 21968 31220
rect 21640 31136 21692 31142
rect 21640 31078 21692 31084
rect 21652 30938 21680 31078
rect 21640 30932 21692 30938
rect 21640 30874 21692 30880
rect 21548 30660 21600 30666
rect 21548 30602 21600 30608
rect 21652 30122 21680 30874
rect 21928 30802 21956 31214
rect 22112 30938 22140 32302
rect 22192 31340 22244 31346
rect 22192 31282 22244 31288
rect 22100 30932 22152 30938
rect 22100 30874 22152 30880
rect 21916 30796 21968 30802
rect 21916 30738 21968 30744
rect 22204 30734 22232 31282
rect 22572 30870 22600 32846
rect 22836 31680 22888 31686
rect 22836 31622 22888 31628
rect 22848 31210 22876 31622
rect 23584 31482 23612 33798
rect 23572 31476 23624 31482
rect 23572 31418 23624 31424
rect 23296 31272 23348 31278
rect 23296 31214 23348 31220
rect 22836 31204 22888 31210
rect 22836 31146 22888 31152
rect 22928 31204 22980 31210
rect 22928 31146 22980 31152
rect 22560 30864 22612 30870
rect 22560 30806 22612 30812
rect 22192 30728 22244 30734
rect 22192 30670 22244 30676
rect 22744 30728 22796 30734
rect 22744 30670 22796 30676
rect 21824 30252 21876 30258
rect 21824 30194 21876 30200
rect 21640 30116 21692 30122
rect 21640 30058 21692 30064
rect 21652 29850 21680 30058
rect 21836 29850 21864 30194
rect 22652 30184 22704 30190
rect 22652 30126 22704 30132
rect 21640 29844 21692 29850
rect 21640 29786 21692 29792
rect 21824 29844 21876 29850
rect 21824 29786 21876 29792
rect 22664 29782 22692 30126
rect 22756 29850 22784 30670
rect 22848 30666 22876 31146
rect 22940 30938 22968 31146
rect 23308 30938 23336 31214
rect 22928 30932 22980 30938
rect 22928 30874 22980 30880
rect 23296 30932 23348 30938
rect 23296 30874 23348 30880
rect 22836 30660 22888 30666
rect 22836 30602 22888 30608
rect 23676 30190 23704 34410
rect 24504 34066 24532 34478
rect 24492 34060 24544 34066
rect 24492 34002 24544 34008
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24412 32026 24440 33934
rect 25608 33454 25636 35974
rect 26160 35154 26188 36110
rect 26792 36100 26844 36106
rect 26792 36042 26844 36048
rect 26804 35290 26832 36042
rect 27632 35630 27660 36178
rect 29552 35692 29604 35698
rect 29552 35634 29604 35640
rect 27160 35624 27212 35630
rect 27160 35566 27212 35572
rect 27620 35624 27672 35630
rect 27620 35566 27672 35572
rect 28356 35624 28408 35630
rect 28356 35566 28408 35572
rect 26792 35284 26844 35290
rect 26792 35226 26844 35232
rect 26148 35148 26200 35154
rect 26148 35090 26200 35096
rect 25872 35080 25924 35086
rect 25872 35022 25924 35028
rect 25884 33930 25912 35022
rect 26884 35012 26936 35018
rect 26884 34954 26936 34960
rect 26896 34066 26924 34954
rect 26884 34060 26936 34066
rect 26884 34002 26936 34008
rect 27172 33998 27200 35566
rect 28368 35154 28396 35566
rect 29564 35154 29592 35634
rect 29920 35488 29972 35494
rect 29920 35430 29972 35436
rect 28356 35148 28408 35154
rect 28356 35090 28408 35096
rect 29552 35148 29604 35154
rect 29552 35090 29604 35096
rect 29828 35012 29880 35018
rect 29828 34954 29880 34960
rect 29840 34746 29868 34954
rect 29828 34740 29880 34746
rect 29828 34682 29880 34688
rect 29644 34604 29696 34610
rect 29644 34546 29696 34552
rect 29656 34202 29684 34546
rect 29644 34196 29696 34202
rect 29644 34138 29696 34144
rect 26056 33992 26108 33998
rect 26056 33934 26108 33940
rect 27160 33992 27212 33998
rect 27160 33934 27212 33940
rect 29000 33992 29052 33998
rect 29000 33934 29052 33940
rect 25872 33924 25924 33930
rect 25872 33866 25924 33872
rect 24492 33448 24544 33454
rect 24492 33390 24544 33396
rect 24676 33448 24728 33454
rect 24676 33390 24728 33396
rect 25596 33448 25648 33454
rect 25596 33390 25648 33396
rect 24504 33114 24532 33390
rect 24492 33108 24544 33114
rect 24492 33050 24544 33056
rect 24688 32434 24716 33390
rect 25608 32978 25636 33390
rect 25596 32972 25648 32978
rect 25596 32914 25648 32920
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 24400 32020 24452 32026
rect 24400 31962 24452 31968
rect 24492 32020 24544 32026
rect 24492 31962 24544 31968
rect 24504 31872 24532 31962
rect 24412 31844 24532 31872
rect 23756 31408 23808 31414
rect 23756 31350 23808 31356
rect 23768 31278 23796 31350
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 24412 31142 24440 31844
rect 24584 31816 24636 31822
rect 24584 31758 24636 31764
rect 24492 31748 24544 31754
rect 24492 31690 24544 31696
rect 24504 31414 24532 31690
rect 24492 31408 24544 31414
rect 24492 31350 24544 31356
rect 24400 31136 24452 31142
rect 24400 31078 24452 31084
rect 24412 30938 24440 31078
rect 24400 30932 24452 30938
rect 24400 30874 24452 30880
rect 24216 30728 24268 30734
rect 24216 30670 24268 30676
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 22744 29844 22796 29850
rect 22744 29786 22796 29792
rect 22652 29776 22704 29782
rect 22652 29718 22704 29724
rect 21548 29708 21600 29714
rect 21600 29668 21680 29696
rect 21548 29650 21600 29656
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 21364 29572 21416 29578
rect 21364 29514 21416 29520
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 20732 28966 20760 29106
rect 20720 28960 20772 28966
rect 20720 28902 20772 28908
rect 20732 27878 20760 28902
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20732 27554 20760 27814
rect 20640 27526 20760 27554
rect 20640 27470 20668 27526
rect 21376 27470 21404 29514
rect 21652 28014 21680 29668
rect 23296 29028 23348 29034
rect 23296 28970 23348 28976
rect 22744 28416 22796 28422
rect 22744 28358 22796 28364
rect 21640 28008 21692 28014
rect 21640 27950 21692 27956
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 21364 27464 21416 27470
rect 21364 27406 21416 27412
rect 21376 25294 21404 27406
rect 21652 25362 21680 27950
rect 22468 25764 22520 25770
rect 22468 25706 22520 25712
rect 21824 25492 21876 25498
rect 21824 25434 21876 25440
rect 21640 25356 21692 25362
rect 21640 25298 21692 25304
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21652 24750 21680 25298
rect 21732 25220 21784 25226
rect 21732 25162 21784 25168
rect 21744 24886 21772 25162
rect 21732 24880 21784 24886
rect 21732 24822 21784 24828
rect 21640 24744 21692 24750
rect 21640 24686 21692 24692
rect 21652 24274 21680 24686
rect 21836 24614 21864 25434
rect 21916 25288 21968 25294
rect 21916 25230 21968 25236
rect 21928 24886 21956 25230
rect 22008 25152 22060 25158
rect 22008 25094 22060 25100
rect 21916 24880 21968 24886
rect 21916 24822 21968 24828
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21640 24268 21692 24274
rect 21640 24210 21692 24216
rect 21836 24206 21864 24550
rect 22020 24206 22048 25094
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 22008 24200 22060 24206
rect 22008 24142 22060 24148
rect 22480 24138 22508 25706
rect 22468 24132 22520 24138
rect 22468 24074 22520 24080
rect 22480 23662 22508 24074
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 20824 22642 20852 22918
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 22468 22636 22520 22642
rect 22468 22578 22520 22584
rect 22480 21894 22508 22578
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22480 21690 22508 21830
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22756 21350 22784 28358
rect 23020 25696 23072 25702
rect 23020 25638 23072 25644
rect 22836 25220 22888 25226
rect 22836 25162 22888 25168
rect 22848 24290 22876 25162
rect 23032 24818 23060 25638
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 22928 24744 22980 24750
rect 22928 24686 22980 24692
rect 22940 24410 22968 24686
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 22848 24262 22968 24290
rect 22940 23730 22968 24262
rect 23112 24268 23164 24274
rect 23112 24210 23164 24216
rect 22928 23724 22980 23730
rect 22928 23666 22980 23672
rect 22940 22982 22968 23666
rect 23124 23526 23152 24210
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 22928 22976 22980 22982
rect 22928 22918 22980 22924
rect 22940 22642 22968 22918
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 23124 22438 23152 23462
rect 23112 22432 23164 22438
rect 23112 22374 23164 22380
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 20904 19984 20956 19990
rect 20904 19926 20956 19932
rect 20916 19718 20944 19926
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20640 18630 20668 19178
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20732 17338 20760 18702
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20824 15570 20852 15846
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20536 14884 20588 14890
rect 20536 14826 20588 14832
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18524 11830 18552 12174
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 17880 9994 17908 10610
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 18432 9926 18460 10610
rect 18524 10606 18552 11766
rect 18616 11762 18644 12718
rect 19444 12238 19472 12786
rect 20364 12442 20392 12786
rect 20456 12714 20484 13194
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 20272 11830 20300 12038
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 18616 11082 18644 11698
rect 19444 11558 19472 11698
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 20272 11082 20300 11766
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20364 11354 20392 11494
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 18604 11076 18656 11082
rect 18604 11018 18656 11024
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 18616 10742 18644 11018
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 18604 10736 18656 10742
rect 18604 10678 18656 10684
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 19444 10130 19472 10950
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19720 10062 19748 10406
rect 19708 10056 19760 10062
rect 19338 10024 19394 10033
rect 19708 9998 19760 10004
rect 20272 9994 20300 11018
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 10266 20392 10406
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 19338 9959 19394 9968
rect 20260 9988 20312 9994
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 18616 7886 18644 9862
rect 19352 8090 19380 9959
rect 20260 9930 20312 9936
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19996 8974 20024 9862
rect 20364 9382 20392 10202
rect 20456 9994 20484 12650
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 20456 9654 20484 9930
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20364 9178 20392 9318
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 20456 8906 20484 9590
rect 20548 9568 20576 13330
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20640 11626 20668 11834
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20640 11150 20668 11562
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20628 9580 20680 9586
rect 20548 9540 20628 9568
rect 20628 9522 20680 9528
rect 20640 9042 20668 9522
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19444 8022 19472 8774
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 20732 8294 20760 15370
rect 20916 12238 20944 19654
rect 22112 19174 22140 20198
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21836 18358 21864 18566
rect 21824 18352 21876 18358
rect 21824 18294 21876 18300
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 21008 15162 21036 15370
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21836 14074 21864 14282
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 21008 13530 21036 13874
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 22112 12322 22140 19110
rect 22388 18290 22416 19790
rect 22480 19378 22508 20878
rect 22756 19854 22784 21286
rect 23308 20398 23336 28970
rect 23676 28150 23704 30126
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 24032 28620 24084 28626
rect 24032 28562 24084 28568
rect 23940 28484 23992 28490
rect 23940 28426 23992 28432
rect 23664 28144 23716 28150
rect 23664 28086 23716 28092
rect 23676 26234 23704 28086
rect 23952 27062 23980 28426
rect 24044 27538 24072 28562
rect 24032 27532 24084 27538
rect 24032 27474 24084 27480
rect 23940 27056 23992 27062
rect 23940 26998 23992 27004
rect 23676 26206 23888 26234
rect 23480 24744 23532 24750
rect 23480 24686 23532 24692
rect 23492 24342 23520 24686
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23480 24336 23532 24342
rect 23480 24278 23532 24284
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23400 22710 23428 23666
rect 23388 22704 23440 22710
rect 23388 22646 23440 22652
rect 23492 22522 23520 24278
rect 23676 24206 23704 24550
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23676 23866 23704 24142
rect 23664 23860 23716 23866
rect 23664 23802 23716 23808
rect 23492 22494 23704 22522
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23308 19854 23336 20334
rect 23492 20262 23520 22374
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23584 21622 23612 21966
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23676 21486 23704 22494
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23308 19446 23336 19790
rect 23296 19440 23348 19446
rect 23296 19382 23348 19388
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22664 19174 22692 19314
rect 22652 19168 22704 19174
rect 22652 19110 22704 19116
rect 23308 18970 23336 19382
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23296 18964 23348 18970
rect 23296 18906 23348 18912
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 22296 17066 22324 18022
rect 22756 17542 22784 18702
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22756 17202 22784 17478
rect 23400 17270 23428 19314
rect 23112 17264 23164 17270
rect 23112 17206 23164 17212
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22192 15564 22244 15570
rect 22192 15506 22244 15512
rect 22204 14958 22232 15506
rect 22572 15026 22600 15982
rect 22940 15502 22968 16934
rect 23124 16590 23152 17206
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 23216 16590 23244 17138
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23400 16794 23428 16934
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 23492 16658 23520 17070
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23204 16584 23256 16590
rect 23204 16526 23256 16532
rect 23204 16040 23256 16046
rect 23204 15982 23256 15988
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23216 15706 23244 15982
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 22296 12850 22324 13262
rect 23492 12889 23520 15982
rect 23676 14482 23704 21422
rect 23860 17746 23888 26206
rect 23952 20942 23980 26998
rect 24044 26926 24072 27474
rect 24136 27130 24164 29106
rect 24228 28966 24256 30670
rect 24308 29028 24360 29034
rect 24308 28970 24360 28976
rect 24216 28960 24268 28966
rect 24216 28902 24268 28908
rect 24228 28558 24256 28902
rect 24216 28552 24268 28558
rect 24216 28494 24268 28500
rect 24124 27124 24176 27130
rect 24124 27066 24176 27072
rect 24228 26994 24256 28494
rect 24320 27538 24348 28970
rect 24412 28762 24440 30874
rect 24504 30802 24532 31350
rect 24596 31210 24624 31758
rect 25044 31272 25096 31278
rect 25044 31214 25096 31220
rect 24584 31204 24636 31210
rect 24584 31146 24636 31152
rect 24492 30796 24544 30802
rect 24492 30738 24544 30744
rect 24504 29238 24532 30738
rect 24596 30734 24624 31146
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24492 29232 24544 29238
rect 24492 29174 24544 29180
rect 24400 28756 24452 28762
rect 24400 28698 24452 28704
rect 24308 27532 24360 27538
rect 24308 27474 24360 27480
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24032 26920 24084 26926
rect 24032 26862 24084 26868
rect 24412 26790 24440 28698
rect 24860 28416 24912 28422
rect 24860 28358 24912 28364
rect 24872 27470 24900 28358
rect 24860 27464 24912 27470
rect 24860 27406 24912 27412
rect 25056 27402 25084 31214
rect 25424 30938 25452 32370
rect 25596 31680 25648 31686
rect 25596 31622 25648 31628
rect 25608 31346 25636 31622
rect 26068 31482 26096 33934
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 27172 32978 27200 33254
rect 27160 32972 27212 32978
rect 27160 32914 27212 32920
rect 27252 32836 27304 32842
rect 27252 32778 27304 32784
rect 27264 32570 27292 32778
rect 27252 32564 27304 32570
rect 27252 32506 27304 32512
rect 26056 31476 26108 31482
rect 26056 31418 26108 31424
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 28632 31136 28684 31142
rect 28632 31078 28684 31084
rect 25412 30932 25464 30938
rect 25412 30874 25464 30880
rect 28644 30734 28672 31078
rect 29012 30938 29040 33934
rect 29828 31884 29880 31890
rect 29828 31826 29880 31832
rect 29552 31680 29604 31686
rect 29552 31622 29604 31628
rect 29000 30932 29052 30938
rect 29000 30874 29052 30880
rect 28448 30728 28500 30734
rect 28448 30670 28500 30676
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 27988 30592 28040 30598
rect 27988 30534 28040 30540
rect 25504 28552 25556 28558
rect 25504 28494 25556 28500
rect 25516 28082 25544 28494
rect 25504 28076 25556 28082
rect 25504 28018 25556 28024
rect 25320 28008 25372 28014
rect 25320 27950 25372 27956
rect 26240 28008 26292 28014
rect 26240 27950 26292 27956
rect 25332 27606 25360 27950
rect 26148 27872 26200 27878
rect 26148 27814 26200 27820
rect 26160 27606 26188 27814
rect 25320 27600 25372 27606
rect 25320 27542 25372 27548
rect 26148 27600 26200 27606
rect 26148 27542 26200 27548
rect 24676 27396 24728 27402
rect 24676 27338 24728 27344
rect 25044 27396 25096 27402
rect 25044 27338 25096 27344
rect 24492 26920 24544 26926
rect 24492 26862 24544 26868
rect 24400 26784 24452 26790
rect 24400 26726 24452 26732
rect 24504 25906 24532 26862
rect 24492 25900 24544 25906
rect 24492 25842 24544 25848
rect 24308 24200 24360 24206
rect 24308 24142 24360 24148
rect 24320 21078 24348 24142
rect 24504 23186 24532 25842
rect 24492 23180 24544 23186
rect 24492 23122 24544 23128
rect 24400 21140 24452 21146
rect 24400 21082 24452 21088
rect 24308 21072 24360 21078
rect 24308 21014 24360 21020
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 23952 20534 23980 20878
rect 23940 20528 23992 20534
rect 23940 20470 23992 20476
rect 23952 19854 23980 20470
rect 24308 20392 24360 20398
rect 24308 20334 24360 20340
rect 24320 19922 24348 20334
rect 24412 20262 24440 21082
rect 24504 21010 24532 23122
rect 24492 21004 24544 21010
rect 24492 20946 24544 20952
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24596 20466 24624 20878
rect 24584 20460 24636 20466
rect 24584 20402 24636 20408
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 24412 20058 24440 20198
rect 24400 20052 24452 20058
rect 24400 19994 24452 20000
rect 24308 19916 24360 19922
rect 24308 19858 24360 19864
rect 23940 19848 23992 19854
rect 23940 19790 23992 19796
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 24308 19372 24360 19378
rect 24308 19314 24360 19320
rect 24136 18766 24164 19314
rect 24320 18834 24348 19314
rect 24412 19174 24440 19994
rect 24596 19854 24624 20402
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24596 19718 24624 19790
rect 24584 19712 24636 19718
rect 24584 19654 24636 19660
rect 24596 19378 24624 19654
rect 24584 19372 24636 19378
rect 24584 19314 24636 19320
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24412 18970 24440 19110
rect 24400 18964 24452 18970
rect 24400 18906 24452 18912
rect 24308 18828 24360 18834
rect 24308 18770 24360 18776
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 24320 17134 24348 18770
rect 24596 18766 24624 19314
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23860 15570 23888 16934
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 24412 15094 24440 18158
rect 24688 15638 24716 27338
rect 25688 26308 25740 26314
rect 25688 26250 25740 26256
rect 25412 25696 25464 25702
rect 25412 25638 25464 25644
rect 24952 25356 25004 25362
rect 24952 25298 25004 25304
rect 24964 25158 24992 25298
rect 25424 25226 25452 25638
rect 25700 25378 25728 26250
rect 25872 25832 25924 25838
rect 25872 25774 25924 25780
rect 25884 25498 25912 25774
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 25872 25492 25924 25498
rect 25872 25434 25924 25440
rect 25700 25350 25820 25378
rect 26068 25362 26096 25638
rect 26148 25424 26200 25430
rect 26148 25366 26200 25372
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 24952 25152 25004 25158
rect 24952 25094 25004 25100
rect 24964 24750 24992 25094
rect 25424 24886 25452 25162
rect 25412 24880 25464 24886
rect 25412 24822 25464 24828
rect 25700 24818 25728 25230
rect 25792 25158 25820 25350
rect 26056 25356 26108 25362
rect 26056 25298 26108 25304
rect 25780 25152 25832 25158
rect 25780 25094 25832 25100
rect 26056 25152 26108 25158
rect 26056 25094 26108 25100
rect 26068 24818 26096 25094
rect 25688 24812 25740 24818
rect 25688 24754 25740 24760
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 24952 24744 25004 24750
rect 24952 24686 25004 24692
rect 25596 24744 25648 24750
rect 25596 24686 25648 24692
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24872 23186 24900 23598
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24964 21962 24992 24686
rect 25412 24608 25464 24614
rect 25608 24596 25636 24686
rect 25464 24568 25636 24596
rect 25412 24550 25464 24556
rect 25424 24410 25452 24550
rect 25412 24404 25464 24410
rect 25412 24346 25464 24352
rect 25700 24274 25728 24754
rect 25688 24268 25740 24274
rect 25688 24210 25740 24216
rect 25228 24132 25280 24138
rect 25228 24074 25280 24080
rect 25240 23866 25268 24074
rect 26068 23866 26096 24754
rect 26160 24750 26188 25366
rect 26148 24744 26200 24750
rect 26148 24686 26200 24692
rect 26252 24614 26280 27950
rect 26700 27464 26752 27470
rect 26700 27406 26752 27412
rect 26712 25498 26740 27406
rect 28000 26926 28028 30534
rect 28460 30394 28488 30670
rect 28448 30388 28500 30394
rect 28448 30330 28500 30336
rect 28828 30122 28856 30670
rect 29564 30326 29592 31622
rect 29840 31278 29868 31826
rect 29932 31754 29960 35430
rect 30104 34944 30156 34950
rect 30104 34886 30156 34892
rect 29920 31748 29972 31754
rect 29920 31690 29972 31696
rect 29644 31272 29696 31278
rect 29644 31214 29696 31220
rect 29828 31272 29880 31278
rect 29828 31214 29880 31220
rect 29656 30938 29684 31214
rect 29644 30932 29696 30938
rect 29644 30874 29696 30880
rect 29644 30592 29696 30598
rect 29644 30534 29696 30540
rect 29552 30320 29604 30326
rect 29552 30262 29604 30268
rect 28816 30116 28868 30122
rect 28816 30058 28868 30064
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 28736 29714 28764 29990
rect 28724 29708 28776 29714
rect 28724 29650 28776 29656
rect 27988 26920 28040 26926
rect 27988 26862 28040 26868
rect 28080 26920 28132 26926
rect 28080 26862 28132 26868
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 26884 26308 26936 26314
rect 26884 26250 26936 26256
rect 26700 25492 26752 25498
rect 26700 25434 26752 25440
rect 26896 25378 26924 26250
rect 26896 25350 27108 25378
rect 26976 25288 27028 25294
rect 26976 25230 27028 25236
rect 26608 24676 26660 24682
rect 26608 24618 26660 24624
rect 26240 24608 26292 24614
rect 26240 24550 26292 24556
rect 26620 24206 26648 24618
rect 26988 24410 27016 25230
rect 27080 24750 27108 25350
rect 27068 24744 27120 24750
rect 27068 24686 27120 24692
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 27080 24290 27108 24686
rect 27724 24682 27752 26318
rect 27712 24676 27764 24682
rect 27712 24618 27764 24624
rect 26988 24262 27108 24290
rect 26608 24200 26660 24206
rect 26608 24142 26660 24148
rect 26988 24138 27016 24262
rect 27068 24200 27120 24206
rect 27068 24142 27120 24148
rect 26240 24132 26292 24138
rect 26240 24074 26292 24080
rect 26976 24132 27028 24138
rect 26976 24074 27028 24080
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 26056 23860 26108 23866
rect 26056 23802 26108 23808
rect 25240 22982 25268 23802
rect 26252 23730 26280 24074
rect 26240 23724 26292 23730
rect 26240 23666 26292 23672
rect 27080 23526 27108 24142
rect 27068 23520 27120 23526
rect 27068 23462 27120 23468
rect 25964 23044 26016 23050
rect 25964 22986 26016 22992
rect 25228 22976 25280 22982
rect 25228 22918 25280 22924
rect 25240 22778 25268 22918
rect 25228 22772 25280 22778
rect 25228 22714 25280 22720
rect 25976 21962 26004 22986
rect 27080 22001 27108 23462
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27066 21992 27122 22001
rect 24952 21956 25004 21962
rect 24952 21898 25004 21904
rect 25964 21956 26016 21962
rect 27066 21927 27122 21936
rect 25964 21898 26016 21904
rect 25976 21554 26004 21898
rect 25964 21548 26016 21554
rect 25964 21490 26016 21496
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 25056 21146 25084 21422
rect 25044 21140 25096 21146
rect 25044 21082 25096 21088
rect 25976 20806 26004 21490
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26344 21146 26372 21286
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25964 20800 26016 20806
rect 25964 20742 26016 20748
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24872 16114 24900 16390
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 24676 15632 24728 15638
rect 24676 15574 24728 15580
rect 24400 15088 24452 15094
rect 24400 15030 24452 15036
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23478 12880 23534 12889
rect 22284 12844 22336 12850
rect 23478 12815 23534 12824
rect 22284 12786 22336 12792
rect 23492 12782 23520 12815
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 22480 12442 22508 12718
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22112 12294 22232 12322
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 21916 12164 21968 12170
rect 21916 12106 21968 12112
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 21928 11830 21956 12106
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21652 11082 21680 11222
rect 22020 11218 22048 11698
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 21640 11076 21692 11082
rect 21640 11018 21692 11024
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20824 10674 20852 10950
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20824 9586 20852 9998
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20824 8974 20852 9522
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18328 7744 18380 7750
rect 18380 7704 18460 7732
rect 18328 7686 18380 7692
rect 18432 6798 18460 7704
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19996 7546 20024 7890
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19352 7274 19380 7482
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 17236 6322 17264 6734
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 17880 4622 17908 6598
rect 18432 6390 18460 6734
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18432 5250 18460 6326
rect 19352 5710 19380 7210
rect 20180 6730 20208 7686
rect 20258 6896 20314 6905
rect 20258 6831 20314 6840
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 20088 6390 20116 6598
rect 20076 6384 20128 6390
rect 20076 6326 20128 6332
rect 19708 5908 19760 5914
rect 19708 5850 19760 5856
rect 19720 5794 19748 5850
rect 19720 5778 19932 5794
rect 19432 5772 19484 5778
rect 19720 5772 19944 5778
rect 19720 5766 19892 5772
rect 19432 5714 19484 5720
rect 19892 5714 19944 5720
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19260 5302 19288 5510
rect 19352 5302 19380 5510
rect 19444 5370 19472 5714
rect 19708 5704 19760 5710
rect 19760 5652 19932 5658
rect 19708 5646 19932 5652
rect 19720 5642 19932 5646
rect 19720 5636 19944 5642
rect 19720 5630 19892 5636
rect 19892 5578 19944 5584
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19248 5296 19300 5302
rect 18432 5234 18552 5250
rect 19248 5238 19300 5244
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 18432 5228 18564 5234
rect 18432 5222 18512 5228
rect 18512 5170 18564 5176
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17328 4146 17356 4422
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 18248 4078 18276 4558
rect 19168 4146 19196 4966
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17512 3534 17540 3878
rect 19352 3738 19380 5238
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19720 4826 19748 5170
rect 20088 4865 20116 6326
rect 20272 5302 20300 6831
rect 20456 6662 20484 7754
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20456 5710 20484 6598
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20640 5574 20668 7346
rect 20732 7342 20760 8230
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21284 7546 21312 7754
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21560 7410 21588 9862
rect 21744 7954 21772 9862
rect 22112 9654 22140 12106
rect 22204 11082 22232 12294
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23032 11898 23060 12174
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 22192 11076 22244 11082
rect 22192 11018 22244 11024
rect 22204 10810 22232 11018
rect 22652 11008 22704 11014
rect 22652 10950 22704 10956
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 22112 8566 22140 9590
rect 22664 9586 22692 10950
rect 24412 10130 24440 15030
rect 25228 11756 25280 11762
rect 25228 11698 25280 11704
rect 25240 11218 25268 11698
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 25240 11098 25268 11154
rect 25148 11070 25268 11098
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 24032 8900 24084 8906
rect 24032 8842 24084 8848
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 22100 8560 22152 8566
rect 22100 8502 22152 8508
rect 23768 8498 23796 8774
rect 24044 8498 24072 8842
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 20732 6118 20760 6666
rect 21836 6458 21864 6666
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21088 6180 21140 6186
rect 21008 6140 21088 6168
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20904 6112 20956 6118
rect 21008 6100 21036 6140
rect 21088 6122 21140 6128
rect 20956 6072 21036 6100
rect 20904 6054 20956 6060
rect 22112 6066 22140 7278
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22204 6186 22232 6734
rect 22296 6322 22324 7686
rect 24412 7546 24440 10066
rect 25148 8634 25176 11070
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 25240 8634 25268 8910
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25044 8356 25096 8362
rect 25044 8298 25096 8304
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 23124 7410 23152 7482
rect 23112 7404 23164 7410
rect 23112 7346 23164 7352
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23308 7002 23336 7142
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 23308 6730 23336 6938
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 23938 6352 23994 6361
rect 22284 6316 22336 6322
rect 23938 6287 23940 6296
rect 22284 6258 22336 6264
rect 23992 6287 23994 6296
rect 23940 6258 23992 6264
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 20732 5846 20760 6054
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20732 5370 20760 5578
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20074 4856 20130 4865
rect 19708 4820 19760 4826
rect 20074 4791 20130 4800
rect 19708 4762 19760 4768
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19904 3534 19932 3878
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 17788 3126 17816 3470
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 20916 3126 20944 6054
rect 22112 6038 22232 6066
rect 22204 5642 22232 6038
rect 23756 5772 23808 5778
rect 23756 5714 23808 5720
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 21008 3738 21036 4558
rect 22940 3738 22968 4626
rect 23492 4554 23520 5510
rect 23768 4826 23796 5714
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24780 4826 24808 5578
rect 25056 5166 25084 8298
rect 25332 7954 25360 20742
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 25976 18358 26004 18566
rect 25964 18352 26016 18358
rect 25964 18294 26016 18300
rect 26056 15904 26108 15910
rect 26056 15846 26108 15852
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25424 15162 25452 15438
rect 25412 15156 25464 15162
rect 25412 15098 25464 15104
rect 26068 15094 26096 15846
rect 26056 15088 26108 15094
rect 26056 15030 26108 15036
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 25884 12170 25912 13194
rect 26160 12306 26188 14214
rect 26148 12300 26200 12306
rect 26148 12242 26200 12248
rect 25504 12164 25556 12170
rect 25504 12106 25556 12112
rect 25872 12164 25924 12170
rect 25872 12106 25924 12112
rect 25516 11898 25544 12106
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25412 11620 25464 11626
rect 25412 11562 25464 11568
rect 25424 8498 25452 11562
rect 25884 10826 25912 12106
rect 26160 11762 26188 12242
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 25964 11688 26016 11694
rect 25964 11630 26016 11636
rect 25976 11354 26004 11630
rect 25964 11348 26016 11354
rect 25964 11290 26016 11296
rect 25884 10798 26004 10826
rect 25976 8498 26004 10798
rect 26056 10464 26108 10470
rect 26056 10406 26108 10412
rect 26068 10130 26096 10406
rect 26056 10124 26108 10130
rect 26056 10066 26108 10072
rect 26056 8628 26108 8634
rect 26056 8570 26108 8576
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25872 8492 25924 8498
rect 25872 8434 25924 8440
rect 25964 8492 26016 8498
rect 25964 8434 26016 8440
rect 25320 7948 25372 7954
rect 25320 7890 25372 7896
rect 25332 6905 25360 7890
rect 25424 7342 25452 8434
rect 25596 7880 25648 7886
rect 25596 7822 25648 7828
rect 25412 7336 25464 7342
rect 25412 7278 25464 7284
rect 25318 6896 25374 6905
rect 25318 6831 25374 6840
rect 25608 6390 25636 7822
rect 25884 7546 25912 8434
rect 25976 7818 26004 8434
rect 25964 7812 26016 7818
rect 25964 7754 26016 7760
rect 26068 7546 26096 8570
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 26056 7540 26108 7546
rect 26056 7482 26108 7488
rect 26148 6792 26200 6798
rect 26148 6734 26200 6740
rect 25964 6656 26016 6662
rect 25964 6598 26016 6604
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 25976 5914 26004 6598
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 26160 5778 26188 6734
rect 26148 5772 26200 5778
rect 26148 5714 26200 5720
rect 26344 5370 26372 21082
rect 27448 19990 27476 22578
rect 27528 22432 27580 22438
rect 27580 22392 27660 22420
rect 27528 22374 27580 22380
rect 27632 22098 27660 22392
rect 27620 22092 27672 22098
rect 27620 22034 27672 22040
rect 27528 20868 27580 20874
rect 27528 20810 27580 20816
rect 27540 20602 27568 20810
rect 27528 20596 27580 20602
rect 27528 20538 27580 20544
rect 27436 19984 27488 19990
rect 27436 19926 27488 19932
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26436 18766 26464 19450
rect 28000 19446 28028 26862
rect 28092 25906 28120 26862
rect 28736 26234 28764 29650
rect 28816 29572 28868 29578
rect 28816 29514 28868 29520
rect 28828 28082 28856 29514
rect 29000 29504 29052 29510
rect 29000 29446 29052 29452
rect 28908 29096 28960 29102
rect 28908 29038 28960 29044
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 28920 27538 28948 29038
rect 28908 27532 28960 27538
rect 28908 27474 28960 27480
rect 28736 26206 28856 26234
rect 28080 25900 28132 25906
rect 28080 25842 28132 25848
rect 28172 23656 28224 23662
rect 28172 23598 28224 23604
rect 28184 22438 28212 23598
rect 28172 22432 28224 22438
rect 28172 22374 28224 22380
rect 27068 19440 27120 19446
rect 27068 19382 27120 19388
rect 27988 19440 28040 19446
rect 27988 19382 28040 19388
rect 26424 18760 26476 18766
rect 26424 18702 26476 18708
rect 26884 16992 26936 16998
rect 26884 16934 26936 16940
rect 26896 16590 26924 16934
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26620 13326 26648 14214
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26976 13252 27028 13258
rect 26976 13194 27028 13200
rect 26988 12986 27016 13194
rect 26976 12980 27028 12986
rect 26976 12922 27028 12928
rect 26976 12096 27028 12102
rect 26976 12038 27028 12044
rect 26988 11762 27016 12038
rect 26976 11756 27028 11762
rect 26976 11698 27028 11704
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26620 7954 26648 9454
rect 27080 9042 27108 19382
rect 27620 18896 27672 18902
rect 27620 18838 27672 18844
rect 27632 18222 27660 18838
rect 27804 18352 27856 18358
rect 27804 18294 27856 18300
rect 27620 18216 27672 18222
rect 27672 18176 27752 18204
rect 27620 18158 27672 18164
rect 27160 17808 27212 17814
rect 27160 17750 27212 17756
rect 27172 17066 27200 17750
rect 27252 17196 27304 17202
rect 27252 17138 27304 17144
rect 27160 17060 27212 17066
rect 27160 17002 27212 17008
rect 27172 14482 27200 17002
rect 27264 16250 27292 17138
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27252 16244 27304 16250
rect 27252 16186 27304 16192
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27172 14074 27200 14418
rect 27160 14068 27212 14074
rect 27160 14010 27212 14016
rect 27632 13530 27660 16730
rect 27724 16454 27752 18176
rect 27712 16448 27764 16454
rect 27712 16390 27764 16396
rect 27724 16250 27752 16390
rect 27712 16244 27764 16250
rect 27712 16186 27764 16192
rect 27816 16182 27844 18294
rect 27804 16176 27856 16182
rect 27804 16118 27856 16124
rect 27816 15366 27844 16118
rect 27804 15360 27856 15366
rect 27804 15302 27856 15308
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27160 13184 27212 13190
rect 27160 13126 27212 13132
rect 27172 12850 27200 13126
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27160 11552 27212 11558
rect 27160 11494 27212 11500
rect 27172 11082 27200 11494
rect 27160 11076 27212 11082
rect 27160 11018 27212 11024
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 27068 9036 27120 9042
rect 27068 8978 27120 8984
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 26608 7948 26660 7954
rect 26608 7890 26660 7896
rect 26988 7410 27016 8230
rect 26608 7404 26660 7410
rect 26608 7346 26660 7352
rect 26976 7404 27028 7410
rect 26976 7346 27028 7352
rect 26620 6866 26648 7346
rect 27080 7342 27108 8978
rect 27252 8492 27304 8498
rect 27252 8434 27304 8440
rect 27264 7546 27292 8434
rect 27252 7540 27304 7546
rect 27252 7482 27304 7488
rect 27540 7478 27568 9454
rect 27528 7472 27580 7478
rect 27528 7414 27580 7420
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 27712 6792 27764 6798
rect 27712 6734 27764 6740
rect 26792 5704 26844 5710
rect 26792 5646 26844 5652
rect 26332 5364 26384 5370
rect 26332 5306 26384 5312
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 23480 4548 23532 4554
rect 23480 4490 23532 4496
rect 23492 4146 23520 4490
rect 24780 4486 24808 4762
rect 25056 4690 25084 5102
rect 26344 5098 26372 5306
rect 26332 5092 26384 5098
rect 26332 5034 26384 5040
rect 26804 4690 26832 5646
rect 27724 5166 27752 6734
rect 27816 5642 27844 15302
rect 27896 14952 27948 14958
rect 27896 14894 27948 14900
rect 27908 14278 27936 14894
rect 27896 14272 27948 14278
rect 27896 14214 27948 14220
rect 27908 13802 27936 14214
rect 27896 13796 27948 13802
rect 27896 13738 27948 13744
rect 27908 13462 27936 13738
rect 27896 13456 27948 13462
rect 27896 13398 27948 13404
rect 28184 8090 28212 22374
rect 28828 18358 28856 26206
rect 29012 24750 29040 29446
rect 29656 28558 29684 30534
rect 29736 29504 29788 29510
rect 29736 29446 29788 29452
rect 29748 29238 29776 29446
rect 29736 29232 29788 29238
rect 29736 29174 29788 29180
rect 29840 28626 29868 31214
rect 29932 31210 29960 31690
rect 30012 31680 30064 31686
rect 30012 31622 30064 31628
rect 29920 31204 29972 31210
rect 29920 31146 29972 31152
rect 29932 30734 29960 31146
rect 30024 30938 30052 31622
rect 30116 31346 30144 34886
rect 30104 31340 30156 31346
rect 30104 31282 30156 31288
rect 30012 30932 30064 30938
rect 30012 30874 30064 30880
rect 30116 30734 30144 31282
rect 29920 30728 29972 30734
rect 29920 30670 29972 30676
rect 30104 30728 30156 30734
rect 30104 30670 30156 30676
rect 29932 29714 29960 30670
rect 30116 30410 30144 30670
rect 30024 30382 30144 30410
rect 29920 29708 29972 29714
rect 29920 29650 29972 29656
rect 29828 28620 29880 28626
rect 29828 28562 29880 28568
rect 29644 28552 29696 28558
rect 29644 28494 29696 28500
rect 29920 28552 29972 28558
rect 29920 28494 29972 28500
rect 29644 28416 29696 28422
rect 29644 28358 29696 28364
rect 29656 28218 29684 28358
rect 29644 28212 29696 28218
rect 29644 28154 29696 28160
rect 29736 28008 29788 28014
rect 29736 27950 29788 27956
rect 29748 27674 29776 27950
rect 29736 27668 29788 27674
rect 29736 27610 29788 27616
rect 29552 26512 29604 26518
rect 29552 26454 29604 26460
rect 29564 26382 29592 26454
rect 29552 26376 29604 26382
rect 29552 26318 29604 26324
rect 29276 25832 29328 25838
rect 29276 25774 29328 25780
rect 29000 24744 29052 24750
rect 29000 24686 29052 24692
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28920 19446 28948 19790
rect 28908 19440 28960 19446
rect 28908 19382 28960 19388
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 28816 18352 28868 18358
rect 28816 18294 28868 18300
rect 29012 17270 29040 18702
rect 29000 17264 29052 17270
rect 29000 17206 29052 17212
rect 29092 16448 29144 16454
rect 29092 16390 29144 16396
rect 29104 15910 29132 16390
rect 29092 15904 29144 15910
rect 29092 15846 29144 15852
rect 29104 15366 29132 15846
rect 29092 15360 29144 15366
rect 29092 15302 29144 15308
rect 29104 14006 29132 15302
rect 29288 15094 29316 25774
rect 29552 25152 29604 25158
rect 29552 25094 29604 25100
rect 29564 21146 29592 25094
rect 29644 24744 29696 24750
rect 29644 24686 29696 24692
rect 29656 21894 29684 24686
rect 29748 23186 29776 27610
rect 29932 24886 29960 28494
rect 30024 28218 30052 30382
rect 30104 29164 30156 29170
rect 30104 29106 30156 29112
rect 30116 28762 30144 29106
rect 30104 28756 30156 28762
rect 30104 28698 30156 28704
rect 30012 28212 30064 28218
rect 30012 28154 30064 28160
rect 30024 26994 30052 28154
rect 30012 26988 30064 26994
rect 30012 26930 30064 26936
rect 30012 26308 30064 26314
rect 30012 26250 30064 26256
rect 30024 25362 30052 26250
rect 30012 25356 30064 25362
rect 30012 25298 30064 25304
rect 29920 24880 29972 24886
rect 29920 24822 29972 24828
rect 29920 24744 29972 24750
rect 29920 24686 29972 24692
rect 29932 24274 29960 24686
rect 29920 24268 29972 24274
rect 29920 24210 29972 24216
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 29840 23798 29868 24006
rect 29828 23792 29880 23798
rect 29828 23734 29880 23740
rect 29736 23180 29788 23186
rect 29736 23122 29788 23128
rect 29920 23112 29972 23118
rect 29920 23054 29972 23060
rect 29932 22778 29960 23054
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 29920 22772 29972 22778
rect 29920 22714 29972 22720
rect 29736 22636 29788 22642
rect 29736 22578 29788 22584
rect 30012 22636 30064 22642
rect 30012 22578 30064 22584
rect 29748 22234 29776 22578
rect 30024 22438 30052 22578
rect 30012 22432 30064 22438
rect 30012 22374 30064 22380
rect 29736 22228 29788 22234
rect 29736 22170 29788 22176
rect 29644 21888 29696 21894
rect 29644 21830 29696 21836
rect 29552 21140 29604 21146
rect 29552 21082 29604 21088
rect 29656 21010 29684 21830
rect 30116 21622 30144 22918
rect 30104 21616 30156 21622
rect 30104 21558 30156 21564
rect 30208 21434 30236 37062
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 37844 35894 37872 37198
rect 37660 35866 37872 35894
rect 30288 35692 30340 35698
rect 30288 35634 30340 35640
rect 32220 35692 32272 35698
rect 32220 35634 32272 35640
rect 30300 34746 30328 35634
rect 32128 35624 32180 35630
rect 32128 35566 32180 35572
rect 31944 35080 31996 35086
rect 31944 35022 31996 35028
rect 30288 34740 30340 34746
rect 30288 34682 30340 34688
rect 30472 34604 30524 34610
rect 30472 34546 30524 34552
rect 30484 34202 30512 34546
rect 31956 34202 31984 35022
rect 32140 34678 32168 35566
rect 32232 35290 32260 35634
rect 33508 35488 33560 35494
rect 33508 35430 33560 35436
rect 32220 35284 32272 35290
rect 32220 35226 32272 35232
rect 32128 34672 32180 34678
rect 32128 34614 32180 34620
rect 33232 34604 33284 34610
rect 33232 34546 33284 34552
rect 33244 34202 33272 34546
rect 30472 34196 30524 34202
rect 30472 34138 30524 34144
rect 31944 34196 31996 34202
rect 31944 34138 31996 34144
rect 33232 34196 33284 34202
rect 33232 34138 33284 34144
rect 31576 34060 31628 34066
rect 31576 34002 31628 34008
rect 30748 33992 30800 33998
rect 30748 33934 30800 33940
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30472 30252 30524 30258
rect 30472 30194 30524 30200
rect 30300 29170 30328 30194
rect 30380 30116 30432 30122
rect 30380 30058 30432 30064
rect 30288 29164 30340 29170
rect 30288 29106 30340 29112
rect 30288 26512 30340 26518
rect 30288 26454 30340 26460
rect 30300 22642 30328 26454
rect 30392 25294 30420 30058
rect 30484 29306 30512 30194
rect 30760 30054 30788 33934
rect 31588 33454 31616 34002
rect 31668 33992 31720 33998
rect 31668 33934 31720 33940
rect 32496 33992 32548 33998
rect 32496 33934 32548 33940
rect 31576 33448 31628 33454
rect 31576 33390 31628 33396
rect 31392 31680 31444 31686
rect 31392 31622 31444 31628
rect 31404 31346 31432 31622
rect 31300 31340 31352 31346
rect 31300 31282 31352 31288
rect 31392 31340 31444 31346
rect 31392 31282 31444 31288
rect 30840 30796 30892 30802
rect 30840 30738 30892 30744
rect 30748 30048 30800 30054
rect 30748 29990 30800 29996
rect 30748 29572 30800 29578
rect 30748 29514 30800 29520
rect 30472 29300 30524 29306
rect 30472 29242 30524 29248
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 30564 24608 30616 24614
rect 30564 24550 30616 24556
rect 30472 23520 30524 23526
rect 30472 23462 30524 23468
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 30484 22574 30512 23462
rect 30576 22778 30604 24550
rect 30668 24410 30696 24754
rect 30656 24404 30708 24410
rect 30656 24346 30708 24352
rect 30668 23730 30696 24346
rect 30656 23724 30708 23730
rect 30656 23666 30708 23672
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30472 22568 30524 22574
rect 30472 22510 30524 22516
rect 30116 21406 30236 21434
rect 29920 21140 29972 21146
rect 29920 21082 29972 21088
rect 29644 21004 29696 21010
rect 29644 20946 29696 20952
rect 29552 18828 29604 18834
rect 29552 18770 29604 18776
rect 29564 17338 29592 18770
rect 29552 17332 29604 17338
rect 29552 17274 29604 17280
rect 29276 15088 29328 15094
rect 29276 15030 29328 15036
rect 29288 14414 29316 15030
rect 29276 14408 29328 14414
rect 29276 14350 29328 14356
rect 29552 14340 29604 14346
rect 29552 14282 29604 14288
rect 29184 14272 29236 14278
rect 29184 14214 29236 14220
rect 29092 14000 29144 14006
rect 29092 13942 29144 13948
rect 29000 13184 29052 13190
rect 29000 13126 29052 13132
rect 29012 11150 29040 13126
rect 29104 11830 29132 13942
rect 29196 13938 29224 14214
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 29368 13728 29420 13734
rect 29368 13670 29420 13676
rect 29380 12850 29408 13670
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 29092 11824 29144 11830
rect 29092 11766 29144 11772
rect 29000 11144 29052 11150
rect 29000 11086 29052 11092
rect 28632 9580 28684 9586
rect 28632 9522 28684 9528
rect 28644 8634 28672 9522
rect 29368 9512 29420 9518
rect 29368 9454 29420 9460
rect 29092 9036 29144 9042
rect 29092 8978 29144 8984
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28816 8356 28868 8362
rect 28816 8298 28868 8304
rect 28172 8084 28224 8090
rect 28172 8026 28224 8032
rect 28724 7880 28776 7886
rect 28724 7822 28776 7828
rect 28080 7336 28132 7342
rect 28080 7278 28132 7284
rect 28092 6934 28120 7278
rect 28632 7200 28684 7206
rect 28632 7142 28684 7148
rect 28446 7032 28502 7041
rect 28644 7002 28672 7142
rect 28446 6967 28502 6976
rect 28632 6996 28684 7002
rect 28080 6928 28132 6934
rect 28080 6870 28132 6876
rect 27804 5636 27856 5642
rect 27804 5578 27856 5584
rect 27712 5160 27764 5166
rect 27712 5102 27764 5108
rect 26976 5024 27028 5030
rect 26976 4966 27028 4972
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 26792 4684 26844 4690
rect 26792 4626 26844 4632
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24688 4146 24716 4422
rect 26804 4146 26832 4626
rect 26988 4622 27016 4966
rect 26976 4616 27028 4622
rect 26976 4558 27028 4564
rect 27620 4480 27672 4486
rect 27620 4422 27672 4428
rect 27632 4146 27660 4422
rect 27724 4282 27752 5102
rect 28092 4690 28120 6870
rect 28460 5370 28488 6967
rect 28632 6938 28684 6944
rect 28736 6798 28764 7822
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28448 5364 28500 5370
rect 28448 5306 28500 5312
rect 28080 4684 28132 4690
rect 28080 4626 28132 4632
rect 27712 4276 27764 4282
rect 27712 4218 27764 4224
rect 28828 4146 28856 8298
rect 29104 5778 29132 8978
rect 29380 8362 29408 9454
rect 29564 9178 29592 14282
rect 29552 9172 29604 9178
rect 29552 9114 29604 9120
rect 29564 8906 29592 9114
rect 29552 8900 29604 8906
rect 29552 8842 29604 8848
rect 29368 8356 29420 8362
rect 29368 8298 29420 8304
rect 29184 7472 29236 7478
rect 29184 7414 29236 7420
rect 29196 7041 29224 7414
rect 29276 7404 29328 7410
rect 29276 7346 29328 7352
rect 29182 7032 29238 7041
rect 29182 6967 29238 6976
rect 29092 5772 29144 5778
rect 29092 5714 29144 5720
rect 29104 5166 29132 5714
rect 29092 5160 29144 5166
rect 29092 5102 29144 5108
rect 29104 4690 29132 5102
rect 29092 4684 29144 4690
rect 29092 4626 29144 4632
rect 29196 4554 29224 6967
rect 29288 6934 29316 7346
rect 29564 7206 29592 8842
rect 29656 7478 29684 20946
rect 29932 20806 29960 21082
rect 29920 20800 29972 20806
rect 29920 20742 29972 20748
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29736 18964 29788 18970
rect 29736 18906 29788 18912
rect 29748 18222 29776 18906
rect 29840 18630 29868 19246
rect 29828 18624 29880 18630
rect 29828 18566 29880 18572
rect 29840 18426 29868 18566
rect 29932 18426 29960 19450
rect 29828 18420 29880 18426
rect 29828 18362 29880 18368
rect 29920 18420 29972 18426
rect 29920 18362 29972 18368
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 29748 17066 29776 18158
rect 29932 17882 29960 18362
rect 29920 17876 29972 17882
rect 29920 17818 29972 17824
rect 29736 17060 29788 17066
rect 29736 17002 29788 17008
rect 29748 15502 29776 17002
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29748 15162 29776 15438
rect 29736 15156 29788 15162
rect 29736 15098 29788 15104
rect 29828 13252 29880 13258
rect 29828 13194 29880 13200
rect 29840 12986 29868 13194
rect 29828 12980 29880 12986
rect 29828 12922 29880 12928
rect 30116 11286 30144 21406
rect 30484 18970 30512 22510
rect 30760 22506 30788 29514
rect 30852 28014 30880 30738
rect 31116 30592 31168 30598
rect 31116 30534 31168 30540
rect 30932 30184 30984 30190
rect 30932 30126 30984 30132
rect 30944 30054 30972 30126
rect 30932 30048 30984 30054
rect 30932 29990 30984 29996
rect 31128 29238 31156 30534
rect 31116 29232 31168 29238
rect 31116 29174 31168 29180
rect 31312 29034 31340 31282
rect 31404 30734 31432 31282
rect 31392 30728 31444 30734
rect 31392 30670 31444 30676
rect 31404 29782 31432 30670
rect 31588 30054 31616 33390
rect 31680 31482 31708 33934
rect 32508 33658 32536 33934
rect 32496 33652 32548 33658
rect 32496 33594 32548 33600
rect 32312 33516 32364 33522
rect 32312 33458 32364 33464
rect 31760 31680 31812 31686
rect 31760 31622 31812 31628
rect 32220 31680 32272 31686
rect 32220 31622 32272 31628
rect 31668 31476 31720 31482
rect 31668 31418 31720 31424
rect 31772 31414 31800 31622
rect 32232 31482 32260 31622
rect 32220 31476 32272 31482
rect 32220 31418 32272 31424
rect 31760 31408 31812 31414
rect 31760 31350 31812 31356
rect 32324 30938 32352 33458
rect 33520 31906 33548 35430
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34796 34672 34848 34678
rect 34796 34614 34848 34620
rect 34336 34400 34388 34406
rect 34336 34342 34388 34348
rect 33152 31878 33548 31906
rect 33152 31754 33180 31878
rect 33140 31748 33192 31754
rect 33140 31690 33192 31696
rect 33324 31748 33376 31754
rect 33324 31690 33376 31696
rect 32404 31680 32456 31686
rect 32404 31622 32456 31628
rect 32312 30932 32364 30938
rect 32312 30874 32364 30880
rect 32416 30734 32444 31622
rect 33336 31482 33364 31690
rect 33416 31680 33468 31686
rect 33416 31622 33468 31628
rect 33324 31476 33376 31482
rect 33324 31418 33376 31424
rect 32496 31272 32548 31278
rect 32496 31214 32548 31220
rect 33140 31272 33192 31278
rect 33140 31214 33192 31220
rect 32508 30734 32536 31214
rect 33152 30802 33180 31214
rect 33428 30938 33456 31622
rect 33416 30932 33468 30938
rect 33416 30874 33468 30880
rect 33140 30796 33192 30802
rect 33140 30738 33192 30744
rect 33520 30734 33548 31878
rect 33600 31884 33652 31890
rect 33600 31826 33652 31832
rect 32404 30728 32456 30734
rect 32404 30670 32456 30676
rect 32496 30728 32548 30734
rect 32496 30670 32548 30676
rect 33508 30728 33560 30734
rect 33508 30670 33560 30676
rect 31852 30660 31904 30666
rect 31852 30602 31904 30608
rect 31576 30048 31628 30054
rect 31576 29990 31628 29996
rect 31392 29776 31444 29782
rect 31392 29718 31444 29724
rect 31404 29238 31432 29718
rect 31864 29714 31892 30602
rect 32508 30410 32536 30670
rect 33416 30592 33468 30598
rect 33416 30534 33468 30540
rect 32416 30394 32536 30410
rect 32404 30388 32536 30394
rect 32456 30382 32536 30388
rect 32404 30330 32456 30336
rect 31852 29708 31904 29714
rect 31852 29650 31904 29656
rect 31392 29232 31444 29238
rect 31392 29174 31444 29180
rect 31300 29028 31352 29034
rect 31300 28970 31352 28976
rect 30840 28008 30892 28014
rect 30840 27950 30892 27956
rect 30852 25362 30880 27950
rect 30932 26444 30984 26450
rect 30932 26386 30984 26392
rect 30944 25974 30972 26386
rect 31312 26234 31340 28970
rect 31404 28762 31432 29174
rect 31392 28756 31444 28762
rect 31392 28698 31444 28704
rect 31404 27130 31432 28698
rect 31392 27124 31444 27130
rect 31392 27066 31444 27072
rect 31668 27124 31720 27130
rect 31668 27066 31720 27072
rect 31392 26852 31444 26858
rect 31392 26794 31444 26800
rect 31404 26450 31432 26794
rect 31392 26444 31444 26450
rect 31392 26386 31444 26392
rect 31312 26206 31432 26234
rect 30932 25968 30984 25974
rect 30932 25910 30984 25916
rect 30840 25356 30892 25362
rect 30840 25298 30892 25304
rect 30852 24614 30880 25298
rect 30932 25288 30984 25294
rect 30932 25230 30984 25236
rect 30944 24818 30972 25230
rect 31116 25220 31168 25226
rect 31116 25162 31168 25168
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 30944 23186 30972 24754
rect 31128 24614 31156 25162
rect 31116 24608 31168 24614
rect 31116 24550 31168 24556
rect 30932 23180 30984 23186
rect 30932 23122 30984 23128
rect 30840 23112 30892 23118
rect 30840 23054 30892 23060
rect 30748 22500 30800 22506
rect 30748 22442 30800 22448
rect 30852 21146 30880 23054
rect 30944 22710 30972 23122
rect 30932 22704 30984 22710
rect 30932 22646 30984 22652
rect 31024 22092 31076 22098
rect 31024 22034 31076 22040
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 30944 21690 30972 21966
rect 30932 21684 30984 21690
rect 30932 21626 30984 21632
rect 30840 21140 30892 21146
rect 30840 21082 30892 21088
rect 30944 20874 30972 21626
rect 31036 21010 31064 22034
rect 31024 21004 31076 21010
rect 31024 20946 31076 20952
rect 30932 20868 30984 20874
rect 30932 20810 30984 20816
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30840 18692 30892 18698
rect 30840 18634 30892 18640
rect 30564 18080 30616 18086
rect 30564 18022 30616 18028
rect 30576 17678 30604 18022
rect 30852 17882 30880 18634
rect 30840 17876 30892 17882
rect 30840 17818 30892 17824
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30564 17536 30616 17542
rect 30564 17478 30616 17484
rect 30576 17338 30604 17478
rect 30564 17332 30616 17338
rect 30564 17274 30616 17280
rect 30196 17196 30248 17202
rect 30196 17138 30248 17144
rect 30208 16046 30236 17138
rect 30288 16992 30340 16998
rect 30288 16934 30340 16940
rect 30300 16590 30328 16934
rect 30288 16584 30340 16590
rect 30576 16574 30604 17274
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30668 16726 30696 17138
rect 31036 17134 31064 20946
rect 31024 17128 31076 17134
rect 31024 17070 31076 17076
rect 30656 16720 30708 16726
rect 30656 16662 30708 16668
rect 30576 16546 30696 16574
rect 30288 16526 30340 16532
rect 30196 16040 30248 16046
rect 30196 15982 30248 15988
rect 30208 15434 30236 15982
rect 30196 15428 30248 15434
rect 30196 15370 30248 15376
rect 30208 14482 30236 15370
rect 30380 14884 30432 14890
rect 30380 14826 30432 14832
rect 30196 14476 30248 14482
rect 30196 14418 30248 14424
rect 30392 14346 30420 14826
rect 30380 14340 30432 14346
rect 30380 14282 30432 14288
rect 30392 14074 30420 14282
rect 30380 14068 30432 14074
rect 30380 14010 30432 14016
rect 30392 13802 30420 14010
rect 30380 13796 30432 13802
rect 30380 13738 30432 13744
rect 30380 12164 30432 12170
rect 30380 12106 30432 12112
rect 30288 11348 30340 11354
rect 30288 11290 30340 11296
rect 30104 11280 30156 11286
rect 30104 11222 30156 11228
rect 29920 11008 29972 11014
rect 29920 10950 29972 10956
rect 29932 9926 29960 10950
rect 30116 10742 30144 11222
rect 30104 10736 30156 10742
rect 30104 10678 30156 10684
rect 30300 10130 30328 11290
rect 30392 11150 30420 12106
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 30380 11144 30432 11150
rect 30380 11086 30432 11092
rect 30392 10810 30420 11086
rect 30380 10804 30432 10810
rect 30380 10746 30432 10752
rect 30288 10124 30340 10130
rect 30288 10066 30340 10072
rect 29920 9920 29972 9926
rect 29920 9862 29972 9868
rect 29932 9518 29960 9862
rect 29920 9512 29972 9518
rect 29920 9454 29972 9460
rect 29932 9178 29960 9454
rect 29920 9172 29972 9178
rect 29920 9114 29972 9120
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30392 8498 30420 8774
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30484 8430 30512 11698
rect 30472 8424 30524 8430
rect 30472 8366 30524 8372
rect 30484 8090 30512 8366
rect 30472 8084 30524 8090
rect 30472 8026 30524 8032
rect 30484 7970 30512 8026
rect 30484 7942 30604 7970
rect 29644 7472 29696 7478
rect 29644 7414 29696 7420
rect 30380 7404 30432 7410
rect 30380 7346 30432 7352
rect 30472 7404 30524 7410
rect 30472 7346 30524 7352
rect 29552 7200 29604 7206
rect 29552 7142 29604 7148
rect 30392 6934 30420 7346
rect 30484 7002 30512 7346
rect 30576 7002 30604 7942
rect 30472 6996 30524 7002
rect 30472 6938 30524 6944
rect 30564 6996 30616 7002
rect 30564 6938 30616 6944
rect 29276 6928 29328 6934
rect 29276 6870 29328 6876
rect 30380 6928 30432 6934
rect 30380 6870 30432 6876
rect 29184 4548 29236 4554
rect 29184 4490 29236 4496
rect 29092 4480 29144 4486
rect 29092 4422 29144 4428
rect 29104 4146 29132 4422
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23664 4140 23716 4146
rect 23664 4082 23716 4088
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 26792 4140 26844 4146
rect 26792 4082 26844 4088
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 28816 4140 28868 4146
rect 28816 4082 28868 4088
rect 29092 4140 29144 4146
rect 29092 4082 29144 4088
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 23492 3602 23520 4082
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 23492 3194 23520 3538
rect 23676 3466 23704 4082
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23768 3670 23796 4014
rect 24584 3936 24636 3942
rect 24584 3878 24636 3884
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 23756 3664 23808 3670
rect 23756 3606 23808 3612
rect 24596 3534 24624 3878
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 23664 3460 23716 3466
rect 23664 3402 23716 3408
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 24412 3126 24440 3334
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 20904 3120 20956 3126
rect 20904 3062 20956 3068
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 27632 3058 27660 3878
rect 29288 3670 29316 6870
rect 30380 6792 30432 6798
rect 30380 6734 30432 6740
rect 30288 6248 30340 6254
rect 30288 6190 30340 6196
rect 29828 6180 29880 6186
rect 29828 6122 29880 6128
rect 29840 5642 29868 6122
rect 30300 5778 30328 6190
rect 30288 5772 30340 5778
rect 30288 5714 30340 5720
rect 30392 5710 30420 6734
rect 30576 5778 30604 6938
rect 30564 5772 30616 5778
rect 30564 5714 30616 5720
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 29828 5636 29880 5642
rect 29828 5578 29880 5584
rect 29840 5370 29868 5578
rect 30576 5370 30604 5714
rect 30668 5642 30696 16546
rect 30932 13796 30984 13802
rect 30932 13738 30984 13744
rect 30944 13530 30972 13738
rect 30932 13524 30984 13530
rect 30932 13466 30984 13472
rect 31128 11898 31156 24550
rect 31208 19236 31260 19242
rect 31208 19178 31260 19184
rect 31220 18698 31248 19178
rect 31208 18692 31260 18698
rect 31208 18634 31260 18640
rect 31220 17678 31248 18634
rect 31208 17672 31260 17678
rect 31208 17614 31260 17620
rect 31220 16794 31248 17614
rect 31404 17542 31432 26206
rect 31680 24682 31708 27066
rect 31864 26518 31892 29650
rect 32036 29028 32088 29034
rect 32036 28970 32088 28976
rect 31944 27328 31996 27334
rect 31944 27270 31996 27276
rect 31956 27062 31984 27270
rect 31944 27056 31996 27062
rect 31944 26998 31996 27004
rect 31852 26512 31904 26518
rect 31852 26454 31904 26460
rect 31956 25770 31984 26998
rect 32048 26382 32076 28970
rect 32508 28966 32536 30382
rect 33428 30054 33456 30534
rect 33416 30048 33468 30054
rect 33416 29990 33468 29996
rect 32496 28960 32548 28966
rect 32496 28902 32548 28908
rect 32508 28150 32536 28902
rect 32496 28144 32548 28150
rect 32496 28086 32548 28092
rect 32220 28076 32272 28082
rect 32220 28018 32272 28024
rect 33324 28076 33376 28082
rect 33324 28018 33376 28024
rect 32232 26994 32260 28018
rect 33232 27328 33284 27334
rect 33232 27270 33284 27276
rect 32220 26988 32272 26994
rect 32220 26930 32272 26936
rect 32404 26988 32456 26994
rect 32404 26930 32456 26936
rect 32232 26450 32260 26930
rect 32416 26586 32444 26930
rect 32404 26580 32456 26586
rect 32404 26522 32456 26528
rect 33140 26512 33192 26518
rect 33140 26454 33192 26460
rect 32220 26444 32272 26450
rect 32220 26386 32272 26392
rect 32036 26376 32088 26382
rect 32036 26318 32088 26324
rect 32048 25974 32076 26318
rect 32220 26308 32272 26314
rect 32220 26250 32272 26256
rect 32680 26308 32732 26314
rect 32680 26250 32732 26256
rect 32036 25968 32088 25974
rect 32036 25910 32088 25916
rect 32128 25900 32180 25906
rect 32128 25842 32180 25848
rect 32140 25770 32168 25842
rect 31944 25764 31996 25770
rect 31944 25706 31996 25712
rect 32128 25764 32180 25770
rect 32128 25706 32180 25712
rect 32140 25294 32168 25706
rect 32232 25498 32260 26250
rect 32692 25906 32720 26250
rect 32680 25900 32732 25906
rect 32680 25842 32732 25848
rect 32220 25492 32272 25498
rect 32220 25434 32272 25440
rect 32692 25294 32720 25842
rect 32956 25696 33008 25702
rect 32956 25638 33008 25644
rect 32128 25288 32180 25294
rect 32128 25230 32180 25236
rect 32312 25288 32364 25294
rect 32312 25230 32364 25236
rect 32680 25288 32732 25294
rect 32680 25230 32732 25236
rect 31852 25152 31904 25158
rect 31852 25094 31904 25100
rect 31668 24676 31720 24682
rect 31668 24618 31720 24624
rect 31484 22976 31536 22982
rect 31484 22918 31536 22924
rect 31496 21962 31524 22918
rect 31484 21956 31536 21962
rect 31484 21898 31536 21904
rect 31680 19310 31708 24618
rect 31864 24614 31892 25094
rect 31852 24608 31904 24614
rect 31852 24550 31904 24556
rect 31760 21888 31812 21894
rect 31760 21830 31812 21836
rect 31772 21350 31800 21830
rect 31760 21344 31812 21350
rect 31760 21286 31812 21292
rect 31772 20942 31800 21286
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31668 19304 31720 19310
rect 31668 19246 31720 19252
rect 31668 18216 31720 18222
rect 31668 18158 31720 18164
rect 31484 17604 31536 17610
rect 31484 17546 31536 17552
rect 31392 17536 31444 17542
rect 31392 17478 31444 17484
rect 31496 17338 31524 17546
rect 31484 17332 31536 17338
rect 31484 17274 31536 17280
rect 31208 16788 31260 16794
rect 31208 16730 31260 16736
rect 31484 13864 31536 13870
rect 31484 13806 31536 13812
rect 31116 11892 31168 11898
rect 31116 11834 31168 11840
rect 30932 10668 30984 10674
rect 30932 10610 30984 10616
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 30748 9920 30800 9926
rect 30748 9862 30800 9868
rect 30760 9042 30788 9862
rect 30852 9722 30880 9998
rect 30840 9716 30892 9722
rect 30840 9658 30892 9664
rect 30748 9036 30800 9042
rect 30748 8978 30800 8984
rect 30852 8974 30880 9658
rect 30840 8968 30892 8974
rect 30840 8910 30892 8916
rect 30944 8498 30972 10610
rect 31300 10124 31352 10130
rect 31300 10066 31352 10072
rect 31312 9110 31340 10066
rect 31496 10062 31524 13806
rect 31680 13258 31708 18158
rect 31864 14414 31892 24550
rect 32324 24274 32352 25230
rect 32312 24268 32364 24274
rect 32312 24210 32364 24216
rect 32680 24200 32732 24206
rect 32680 24142 32732 24148
rect 32692 23526 32720 24142
rect 32680 23520 32732 23526
rect 32680 23462 32732 23468
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 31944 21888 31996 21894
rect 31944 21830 31996 21836
rect 31956 21690 31984 21830
rect 32140 21690 32168 21966
rect 32312 21888 32364 21894
rect 32312 21830 32364 21836
rect 31944 21684 31996 21690
rect 31944 21626 31996 21632
rect 32128 21684 32180 21690
rect 32128 21626 32180 21632
rect 32324 19378 32352 21830
rect 32588 20936 32640 20942
rect 32588 20878 32640 20884
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32496 19372 32548 19378
rect 32496 19314 32548 19320
rect 32324 18358 32352 19314
rect 32508 18358 32536 19314
rect 32600 18766 32628 20878
rect 32588 18760 32640 18766
rect 32588 18702 32640 18708
rect 32312 18352 32364 18358
rect 32312 18294 32364 18300
rect 32496 18352 32548 18358
rect 32496 18294 32548 18300
rect 32508 16114 32536 18294
rect 32588 18148 32640 18154
rect 32588 18090 32640 18096
rect 32600 17882 32628 18090
rect 32588 17876 32640 17882
rect 32588 17818 32640 17824
rect 32600 17270 32628 17818
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32692 16998 32720 23462
rect 32968 22642 32996 25638
rect 33152 25362 33180 26454
rect 33244 25906 33272 27270
rect 33336 26450 33364 28018
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 33428 26314 33456 29990
rect 33612 28762 33640 31826
rect 34348 31754 34376 34342
rect 34060 31748 34112 31754
rect 34060 31690 34112 31696
rect 34336 31748 34388 31754
rect 34336 31690 34388 31696
rect 33600 28756 33652 28762
rect 33600 28698 33652 28704
rect 33784 28484 33836 28490
rect 33784 28426 33836 28432
rect 33600 28008 33652 28014
rect 33600 27950 33652 27956
rect 33612 27538 33640 27950
rect 33600 27532 33652 27538
rect 33600 27474 33652 27480
rect 33508 26784 33560 26790
rect 33508 26726 33560 26732
rect 33520 26450 33548 26726
rect 33508 26444 33560 26450
rect 33508 26386 33560 26392
rect 33416 26308 33468 26314
rect 33416 26250 33468 26256
rect 33428 25974 33456 26250
rect 33416 25968 33468 25974
rect 33416 25910 33468 25916
rect 33232 25900 33284 25906
rect 33232 25842 33284 25848
rect 33428 25838 33456 25910
rect 33416 25832 33468 25838
rect 33416 25774 33468 25780
rect 33140 25356 33192 25362
rect 33140 25298 33192 25304
rect 33232 25288 33284 25294
rect 33232 25230 33284 25236
rect 33244 24682 33272 25230
rect 33508 25152 33560 25158
rect 33508 25094 33560 25100
rect 33232 24676 33284 24682
rect 33232 24618 33284 24624
rect 33520 24206 33548 25094
rect 33612 24818 33640 27474
rect 33692 27464 33744 27470
rect 33692 27406 33744 27412
rect 33704 27130 33732 27406
rect 33692 27124 33744 27130
rect 33692 27066 33744 27072
rect 33796 26450 33824 28426
rect 34072 27130 34100 31690
rect 34336 31340 34388 31346
rect 34336 31282 34388 31288
rect 34348 30326 34376 31282
rect 34808 31278 34836 34614
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 37660 31958 37688 35866
rect 38108 33992 38160 33998
rect 38106 33960 38108 33969
rect 38160 33960 38162 33969
rect 38106 33895 38162 33904
rect 37740 33856 37792 33862
rect 37740 33798 37792 33804
rect 37648 31952 37700 31958
rect 37648 31894 37700 31900
rect 35256 31816 35308 31822
rect 35256 31758 35308 31764
rect 35268 31278 35296 31758
rect 36176 31748 36228 31754
rect 36176 31690 36228 31696
rect 34796 31272 34848 31278
rect 34796 31214 34848 31220
rect 35256 31272 35308 31278
rect 35256 31214 35308 31220
rect 34336 30320 34388 30326
rect 34336 30262 34388 30268
rect 34808 30190 34836 31214
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 36188 30938 36216 31690
rect 36544 31136 36596 31142
rect 36544 31078 36596 31084
rect 36176 30932 36228 30938
rect 36176 30874 36228 30880
rect 35440 30728 35492 30734
rect 35440 30670 35492 30676
rect 35348 30252 35400 30258
rect 35348 30194 35400 30200
rect 34796 30184 34848 30190
rect 34796 30126 34848 30132
rect 34808 29850 34836 30126
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 35360 29850 35388 30194
rect 34796 29844 34848 29850
rect 34796 29786 34848 29792
rect 35348 29844 35400 29850
rect 35348 29786 35400 29792
rect 34520 29640 34572 29646
rect 34520 29582 34572 29588
rect 34532 27606 34560 29582
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 35452 28218 35480 30670
rect 36556 29646 36584 31078
rect 36728 30796 36780 30802
rect 36728 30738 36780 30744
rect 36740 29714 36768 30738
rect 37188 29776 37240 29782
rect 37188 29718 37240 29724
rect 36728 29708 36780 29714
rect 36728 29650 36780 29656
rect 35900 29640 35952 29646
rect 35900 29582 35952 29588
rect 36544 29640 36596 29646
rect 36544 29582 36596 29588
rect 35912 28558 35940 29582
rect 36176 29504 36228 29510
rect 36176 29446 36228 29452
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35440 28212 35492 28218
rect 35440 28154 35492 28160
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34520 27600 34572 27606
rect 34520 27542 34572 27548
rect 35992 27532 36044 27538
rect 35992 27474 36044 27480
rect 35624 27328 35676 27334
rect 35624 27270 35676 27276
rect 34060 27124 34112 27130
rect 34060 27066 34112 27072
rect 34072 26858 34100 27066
rect 34060 26852 34112 26858
rect 34060 26794 34112 26800
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 33784 26444 33836 26450
rect 33784 26386 33836 26392
rect 35636 26382 35664 27270
rect 36004 26926 36032 27474
rect 36188 27470 36216 29446
rect 36360 28552 36412 28558
rect 36360 28494 36412 28500
rect 36176 27464 36228 27470
rect 36176 27406 36228 27412
rect 36084 27396 36136 27402
rect 36084 27338 36136 27344
rect 35992 26920 36044 26926
rect 35992 26862 36044 26868
rect 35900 26784 35952 26790
rect 35900 26726 35952 26732
rect 35624 26376 35676 26382
rect 35624 26318 35676 26324
rect 35912 26246 35940 26726
rect 36004 26450 36032 26862
rect 35992 26444 36044 26450
rect 35992 26386 36044 26392
rect 35900 26240 35952 26246
rect 35900 26182 35952 26188
rect 35912 25702 35940 26182
rect 35900 25696 35952 25702
rect 35900 25638 35952 25644
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 33600 24812 33652 24818
rect 33600 24754 33652 24760
rect 33612 24274 33640 24754
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 33600 24268 33652 24274
rect 33600 24210 33652 24216
rect 33508 24200 33560 24206
rect 33508 24142 33560 24148
rect 34336 24064 34388 24070
rect 34336 24006 34388 24012
rect 34348 23730 34376 24006
rect 34336 23724 34388 23730
rect 34336 23666 34388 23672
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34796 23520 34848 23526
rect 34796 23462 34848 23468
rect 33876 23112 33928 23118
rect 33876 23054 33928 23060
rect 33888 22778 33916 23054
rect 33692 22772 33744 22778
rect 33692 22714 33744 22720
rect 33876 22772 33928 22778
rect 33876 22714 33928 22720
rect 32956 22636 33008 22642
rect 32956 22578 33008 22584
rect 33704 22030 33732 22714
rect 34532 22710 34560 23462
rect 34808 23118 34836 23462
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34796 23112 34848 23118
rect 34796 23054 34848 23060
rect 34520 22704 34572 22710
rect 34520 22646 34572 22652
rect 34612 22636 34664 22642
rect 34612 22578 34664 22584
rect 33784 22500 33836 22506
rect 33784 22442 33836 22448
rect 33692 22024 33744 22030
rect 33692 21966 33744 21972
rect 32956 19168 33008 19174
rect 32956 19110 33008 19116
rect 32968 18766 32996 19110
rect 33796 18766 33824 22442
rect 34520 22432 34572 22438
rect 34520 22374 34572 22380
rect 34532 22098 34560 22374
rect 34520 22092 34572 22098
rect 34624 22094 34652 22578
rect 34808 22574 34836 23054
rect 34796 22568 34848 22574
rect 34796 22510 34848 22516
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34624 22066 34744 22094
rect 34520 22034 34572 22040
rect 33968 21956 34020 21962
rect 33968 21898 34020 21904
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32956 18760 33008 18766
rect 32956 18702 33008 18708
rect 33784 18760 33836 18766
rect 33784 18702 33836 18708
rect 32784 18426 32812 18702
rect 32772 18420 32824 18426
rect 32772 18362 32824 18368
rect 33980 18222 34008 21898
rect 34532 19310 34560 22034
rect 34520 19304 34572 19310
rect 34520 19246 34572 19252
rect 34532 18902 34560 19246
rect 34520 18896 34572 18902
rect 34520 18838 34572 18844
rect 34612 18760 34664 18766
rect 34612 18702 34664 18708
rect 34624 18290 34652 18702
rect 34612 18284 34664 18290
rect 34612 18226 34664 18232
rect 33968 18216 34020 18222
rect 33968 18158 34020 18164
rect 32680 16992 32732 16998
rect 32680 16934 32732 16940
rect 32496 16108 32548 16114
rect 32496 16050 32548 16056
rect 32692 15706 32720 16934
rect 32680 15700 32732 15706
rect 32680 15642 32732 15648
rect 32220 15496 32272 15502
rect 32220 15438 32272 15444
rect 32232 14414 32260 15438
rect 34336 14612 34388 14618
rect 34336 14554 34388 14560
rect 31852 14408 31904 14414
rect 31852 14350 31904 14356
rect 32220 14408 32272 14414
rect 32220 14350 32272 14356
rect 32232 14074 32260 14350
rect 33140 14272 33192 14278
rect 33140 14214 33192 14220
rect 32220 14068 32272 14074
rect 32220 14010 32272 14016
rect 33152 13326 33180 14214
rect 34348 13938 34376 14554
rect 34428 14272 34480 14278
rect 34428 14214 34480 14220
rect 33324 13932 33376 13938
rect 33324 13874 33376 13880
rect 34336 13932 34388 13938
rect 34336 13874 34388 13880
rect 33336 13530 33364 13874
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33324 13524 33376 13530
rect 33324 13466 33376 13472
rect 33612 13326 33640 13806
rect 33140 13320 33192 13326
rect 33140 13262 33192 13268
rect 33600 13320 33652 13326
rect 33600 13262 33652 13268
rect 31668 13252 31720 13258
rect 31668 13194 31720 13200
rect 31680 10810 31708 13194
rect 34440 13190 34468 14214
rect 34520 13864 34572 13870
rect 34520 13806 34572 13812
rect 34532 13258 34560 13806
rect 34520 13252 34572 13258
rect 34520 13194 34572 13200
rect 34428 13184 34480 13190
rect 34428 13126 34480 13132
rect 34440 12850 34468 13126
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 34532 12434 34560 13194
rect 34624 12866 34652 18226
rect 34716 16794 34744 22066
rect 35808 22024 35860 22030
rect 35808 21966 35860 21972
rect 35820 21690 35848 21966
rect 35808 21684 35860 21690
rect 35808 21626 35860 21632
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 36004 20058 36032 26386
rect 36096 26246 36124 27338
rect 36176 26920 36228 26926
rect 36176 26862 36228 26868
rect 36084 26240 36136 26246
rect 36084 26182 36136 26188
rect 36096 23322 36124 26182
rect 36188 26042 36216 26862
rect 36372 26042 36400 28494
rect 37004 27532 37056 27538
rect 37004 27474 37056 27480
rect 36820 27328 36872 27334
rect 36820 27270 36872 27276
rect 36832 27130 36860 27270
rect 36820 27124 36872 27130
rect 36820 27066 36872 27072
rect 36452 26988 36504 26994
rect 36452 26930 36504 26936
rect 36464 26586 36492 26930
rect 36452 26580 36504 26586
rect 36452 26522 36504 26528
rect 36636 26444 36688 26450
rect 36636 26386 36688 26392
rect 36176 26036 36228 26042
rect 36176 25978 36228 25984
rect 36360 26036 36412 26042
rect 36360 25978 36412 25984
rect 36648 25838 36676 26386
rect 36636 25832 36688 25838
rect 36636 25774 36688 25780
rect 36268 25696 36320 25702
rect 36268 25638 36320 25644
rect 36280 25158 36308 25638
rect 36268 25152 36320 25158
rect 36268 25094 36320 25100
rect 36084 23316 36136 23322
rect 36084 23258 36136 23264
rect 36280 22438 36308 25094
rect 36648 24410 36676 25774
rect 36636 24404 36688 24410
rect 36636 24346 36688 24352
rect 36268 22432 36320 22438
rect 36268 22374 36320 22380
rect 35992 20052 36044 20058
rect 35992 19994 36044 20000
rect 35992 19780 36044 19786
rect 35992 19722 36044 19728
rect 35440 19372 35492 19378
rect 35440 19314 35492 19320
rect 34796 19168 34848 19174
rect 34796 19110 34848 19116
rect 34808 18970 34836 19110
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 35452 18970 35480 19314
rect 36004 19174 36032 19722
rect 35992 19168 36044 19174
rect 35992 19110 36044 19116
rect 36084 19168 36136 19174
rect 36084 19110 36136 19116
rect 34796 18964 34848 18970
rect 34796 18906 34848 18912
rect 35440 18964 35492 18970
rect 35440 18906 35492 18912
rect 35532 18760 35584 18766
rect 35532 18702 35584 18708
rect 35348 18692 35400 18698
rect 35348 18634 35400 18640
rect 35360 18426 35388 18634
rect 35440 18624 35492 18630
rect 35440 18566 35492 18572
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34704 16788 34756 16794
rect 34704 16730 34756 16736
rect 35348 15904 35400 15910
rect 35348 15846 35400 15852
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34796 15020 34848 15026
rect 34796 14962 34848 14968
rect 34808 14498 34836 14962
rect 35360 14890 35388 15846
rect 35452 15502 35480 18566
rect 35544 18426 35572 18702
rect 35808 18692 35860 18698
rect 35808 18634 35860 18640
rect 35532 18420 35584 18426
rect 35532 18362 35584 18368
rect 35820 18290 35848 18634
rect 36096 18426 36124 19110
rect 36084 18420 36136 18426
rect 36084 18362 36136 18368
rect 35808 18284 35860 18290
rect 35808 18226 35860 18232
rect 35624 17672 35676 17678
rect 35624 17614 35676 17620
rect 35636 17338 35664 17614
rect 35624 17332 35676 17338
rect 35624 17274 35676 17280
rect 35532 16788 35584 16794
rect 35532 16730 35584 16736
rect 35544 16114 35572 16730
rect 35636 16658 35664 17274
rect 35624 16652 35676 16658
rect 35624 16594 35676 16600
rect 35532 16108 35584 16114
rect 35532 16050 35584 16056
rect 35544 15994 35572 16050
rect 35544 15966 35664 15994
rect 35440 15496 35492 15502
rect 35492 15444 35572 15450
rect 35440 15438 35572 15444
rect 35452 15422 35572 15438
rect 35544 15026 35572 15422
rect 35532 15020 35584 15026
rect 35532 14962 35584 14968
rect 35348 14884 35400 14890
rect 35348 14826 35400 14832
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 35544 14618 35572 14962
rect 35532 14612 35584 14618
rect 35532 14554 35584 14560
rect 34808 14470 35020 14498
rect 34992 14414 35020 14470
rect 34980 14408 35032 14414
rect 34980 14350 35032 14356
rect 34704 14272 34756 14278
rect 34704 14214 34756 14220
rect 34716 12986 34744 14214
rect 34992 14074 35020 14350
rect 34980 14068 35032 14074
rect 34980 14010 35032 14016
rect 35544 13938 35572 14554
rect 35256 13932 35308 13938
rect 35256 13874 35308 13880
rect 35532 13932 35584 13938
rect 35532 13874 35584 13880
rect 35268 13818 35296 13874
rect 35268 13790 35388 13818
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34796 13252 34848 13258
rect 34796 13194 34848 13200
rect 34704 12980 34756 12986
rect 34704 12922 34756 12928
rect 34624 12850 34744 12866
rect 34624 12844 34756 12850
rect 34624 12838 34704 12844
rect 34704 12786 34756 12792
rect 34440 12406 34560 12434
rect 33876 11348 33928 11354
rect 33876 11290 33928 11296
rect 31668 10804 31720 10810
rect 31668 10746 31720 10752
rect 31484 10056 31536 10062
rect 31484 9998 31536 10004
rect 31392 9988 31444 9994
rect 31392 9930 31444 9936
rect 31300 9104 31352 9110
rect 31300 9046 31352 9052
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 30748 8288 30800 8294
rect 30748 8230 30800 8236
rect 30760 7410 30788 8230
rect 30748 7404 30800 7410
rect 30748 7346 30800 7352
rect 30760 6798 30788 7346
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30656 5636 30708 5642
rect 30656 5578 30708 5584
rect 31024 5568 31076 5574
rect 31024 5510 31076 5516
rect 29828 5364 29880 5370
rect 29828 5306 29880 5312
rect 30564 5364 30616 5370
rect 30564 5306 30616 5312
rect 31036 4622 31064 5510
rect 31024 4616 31076 4622
rect 31024 4558 31076 4564
rect 31208 4480 31260 4486
rect 31208 4422 31260 4428
rect 29644 4140 29696 4146
rect 29644 4082 29696 4088
rect 29656 3738 29684 4082
rect 31116 4072 31168 4078
rect 31116 4014 31168 4020
rect 29644 3732 29696 3738
rect 29644 3674 29696 3680
rect 29276 3664 29328 3670
rect 29276 3606 29328 3612
rect 31128 3602 31156 4014
rect 31116 3596 31168 3602
rect 31116 3538 31168 3544
rect 27896 3460 27948 3466
rect 27896 3402 27948 3408
rect 27908 3194 27936 3402
rect 31128 3194 31156 3538
rect 31220 3466 31248 4422
rect 31208 3460 31260 3466
rect 31208 3402 31260 3408
rect 27896 3188 27948 3194
rect 27896 3130 27948 3136
rect 31116 3188 31168 3194
rect 31116 3130 31168 3136
rect 31404 3126 31432 9930
rect 33508 9376 33560 9382
rect 33508 9318 33560 9324
rect 31668 8832 31720 8838
rect 31668 8774 31720 8780
rect 31680 8401 31708 8774
rect 33520 8430 33548 9318
rect 33508 8424 33560 8430
rect 31666 8392 31722 8401
rect 33508 8366 33560 8372
rect 31666 8327 31722 8336
rect 33600 8356 33652 8362
rect 33600 8298 33652 8304
rect 33612 7478 33640 8298
rect 33600 7472 33652 7478
rect 33600 7414 33652 7420
rect 33612 7274 33640 7414
rect 33600 7268 33652 7274
rect 33600 7210 33652 7216
rect 33324 6860 33376 6866
rect 33324 6802 33376 6808
rect 31760 6792 31812 6798
rect 33336 6746 33364 6802
rect 33612 6798 33640 7210
rect 31760 6734 31812 6740
rect 31772 4078 31800 6734
rect 32876 6730 33364 6746
rect 33600 6792 33652 6798
rect 33600 6734 33652 6740
rect 32864 6724 33364 6730
rect 32916 6718 33364 6724
rect 32864 6666 32916 6672
rect 32220 6656 32272 6662
rect 32220 6598 32272 6604
rect 32232 6322 32260 6598
rect 32220 6316 32272 6322
rect 32220 6258 32272 6264
rect 33612 6254 33640 6734
rect 32496 6248 32548 6254
rect 32496 6190 32548 6196
rect 33600 6248 33652 6254
rect 33600 6190 33652 6196
rect 32220 6112 32272 6118
rect 32220 6054 32272 6060
rect 32232 5846 32260 6054
rect 32220 5840 32272 5846
rect 32220 5782 32272 5788
rect 31760 4072 31812 4078
rect 31760 4014 31812 4020
rect 32508 3738 32536 6190
rect 33888 4146 33916 11290
rect 34336 10532 34388 10538
rect 34336 10474 34388 10480
rect 34348 10062 34376 10474
rect 34336 10056 34388 10062
rect 34336 9998 34388 10004
rect 34244 9580 34296 9586
rect 34244 9522 34296 9528
rect 34256 9110 34284 9522
rect 34348 9518 34376 9998
rect 34440 9586 34468 12406
rect 34716 11354 34744 12786
rect 34808 12714 34836 13194
rect 34796 12708 34848 12714
rect 34796 12650 34848 12656
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 35360 12238 35388 13790
rect 35440 13252 35492 13258
rect 35440 13194 35492 13200
rect 35452 12646 35480 13194
rect 35440 12640 35492 12646
rect 35440 12582 35492 12588
rect 35452 12442 35480 12582
rect 35440 12436 35492 12442
rect 35636 12434 35664 15966
rect 35820 15570 35848 18226
rect 36280 18222 36308 22374
rect 36648 21894 36676 24346
rect 36636 21888 36688 21894
rect 36636 21830 36688 21836
rect 37016 20058 37044 27474
rect 37200 27062 37228 29718
rect 37372 29504 37424 29510
rect 37372 29446 37424 29452
rect 37188 27056 37240 27062
rect 37188 26998 37240 27004
rect 37096 26988 37148 26994
rect 37096 26930 37148 26936
rect 37108 26450 37136 26930
rect 37200 26858 37228 26998
rect 37188 26852 37240 26858
rect 37188 26794 37240 26800
rect 37096 26444 37148 26450
rect 37096 26386 37148 26392
rect 37384 26382 37412 29446
rect 37660 27470 37688 31894
rect 37752 29646 37780 33798
rect 37832 30048 37884 30054
rect 37832 29990 37884 29996
rect 38108 30048 38160 30054
rect 38108 29990 38160 29996
rect 37844 29714 37872 29990
rect 38120 29889 38148 29990
rect 38106 29880 38162 29889
rect 38106 29815 38162 29824
rect 37832 29708 37884 29714
rect 37832 29650 37884 29656
rect 37740 29640 37792 29646
rect 37740 29582 37792 29588
rect 37648 27464 37700 27470
rect 37648 27406 37700 27412
rect 38016 26512 38068 26518
rect 38016 26454 38068 26460
rect 37372 26376 37424 26382
rect 37372 26318 37424 26324
rect 37648 26376 37700 26382
rect 37648 26318 37700 26324
rect 37660 25702 37688 26318
rect 38028 25945 38056 26454
rect 38014 25936 38070 25945
rect 38014 25871 38070 25880
rect 37648 25696 37700 25702
rect 37648 25638 37700 25644
rect 37004 20052 37056 20058
rect 37004 19994 37056 20000
rect 36820 19916 36872 19922
rect 36820 19858 36872 19864
rect 36452 19712 36504 19718
rect 36452 19654 36504 19660
rect 36464 19174 36492 19654
rect 36452 19168 36504 19174
rect 36452 19110 36504 19116
rect 36832 18970 36860 19858
rect 36820 18964 36872 18970
rect 36820 18906 36872 18912
rect 36452 18828 36504 18834
rect 36452 18770 36504 18776
rect 36464 18290 36492 18770
rect 36832 18698 36860 18906
rect 36820 18692 36872 18698
rect 36820 18634 36872 18640
rect 36912 18624 36964 18630
rect 36912 18566 36964 18572
rect 36924 18358 36952 18566
rect 36912 18352 36964 18358
rect 36912 18294 36964 18300
rect 36452 18284 36504 18290
rect 36452 18226 36504 18232
rect 36268 18216 36320 18222
rect 36268 18158 36320 18164
rect 36268 16516 36320 16522
rect 36268 16458 36320 16464
rect 36280 16250 36308 16458
rect 36268 16244 36320 16250
rect 36268 16186 36320 16192
rect 36464 16182 36492 18226
rect 37188 16448 37240 16454
rect 37188 16390 37240 16396
rect 36084 16176 36136 16182
rect 36084 16118 36136 16124
rect 36452 16176 36504 16182
rect 36452 16118 36504 16124
rect 36096 15706 36124 16118
rect 37200 16114 37228 16390
rect 37188 16108 37240 16114
rect 37188 16050 37240 16056
rect 35900 15700 35952 15706
rect 35900 15642 35952 15648
rect 36084 15700 36136 15706
rect 36084 15642 36136 15648
rect 35808 15564 35860 15570
rect 35808 15506 35860 15512
rect 35820 14074 35848 15506
rect 35912 15094 35940 15642
rect 35900 15088 35952 15094
rect 35900 15030 35952 15036
rect 36452 15088 36504 15094
rect 36452 15030 36504 15036
rect 36464 14482 36492 15030
rect 36452 14476 36504 14482
rect 36452 14418 36504 14424
rect 35808 14068 35860 14074
rect 35808 14010 35860 14016
rect 36464 13530 36492 14418
rect 37280 13932 37332 13938
rect 37280 13874 37332 13880
rect 36452 13524 36504 13530
rect 36452 13466 36504 13472
rect 37292 12442 37320 13874
rect 37660 13734 37688 25638
rect 38014 21992 38070 22001
rect 38014 21927 38070 21936
rect 38028 21690 38056 21927
rect 38016 21684 38068 21690
rect 38016 21626 38068 21632
rect 37832 21548 37884 21554
rect 37832 21490 37884 21496
rect 37844 18290 37872 21490
rect 37924 18760 37976 18766
rect 37924 18702 37976 18708
rect 37936 18426 37964 18702
rect 37924 18420 37976 18426
rect 37924 18362 37976 18368
rect 37832 18284 37884 18290
rect 37832 18226 37884 18232
rect 38014 17912 38070 17921
rect 38014 17847 38016 17856
rect 38068 17847 38070 17856
rect 38016 17818 38068 17824
rect 37740 17672 37792 17678
rect 37740 17614 37792 17620
rect 37648 13728 37700 13734
rect 37648 13670 37700 13676
rect 35440 12378 35492 12384
rect 35544 12406 35664 12434
rect 37280 12436 37332 12442
rect 35348 12232 35400 12238
rect 35348 12174 35400 12180
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34704 11348 34756 11354
rect 34704 11290 34756 11296
rect 34704 10668 34756 10674
rect 34704 10610 34756 10616
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34520 9920 34572 9926
rect 34520 9862 34572 9868
rect 34428 9580 34480 9586
rect 34428 9522 34480 9528
rect 34532 9518 34560 9862
rect 34336 9512 34388 9518
rect 34336 9454 34388 9460
rect 34520 9512 34572 9518
rect 34520 9454 34572 9460
rect 34532 9178 34560 9454
rect 34612 9444 34664 9450
rect 34612 9386 34664 9392
rect 34520 9172 34572 9178
rect 34520 9114 34572 9120
rect 34244 9104 34296 9110
rect 34244 9046 34296 9052
rect 34624 8906 34652 9386
rect 34716 9382 34744 10610
rect 34808 9722 34836 10610
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 35072 9988 35124 9994
rect 35072 9930 35124 9936
rect 34796 9716 34848 9722
rect 34796 9658 34848 9664
rect 34704 9376 34756 9382
rect 34704 9318 34756 9324
rect 34716 8974 34744 9318
rect 34808 9042 34836 9658
rect 35084 9654 35112 9930
rect 35072 9648 35124 9654
rect 35072 9590 35124 9596
rect 35348 9648 35400 9654
rect 35348 9590 35400 9596
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34796 9036 34848 9042
rect 34796 8978 34848 8984
rect 34704 8968 34756 8974
rect 34704 8910 34756 8916
rect 35164 8968 35216 8974
rect 35164 8910 35216 8916
rect 35256 8968 35308 8974
rect 35256 8910 35308 8916
rect 34612 8900 34664 8906
rect 34612 8842 34664 8848
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34532 8498 34560 8774
rect 35176 8566 35204 8910
rect 35164 8560 35216 8566
rect 35164 8502 35216 8508
rect 35268 8514 35296 8910
rect 35360 8634 35388 9590
rect 35544 8650 35572 12406
rect 37280 12378 37332 12384
rect 36360 9920 36412 9926
rect 36360 9862 36412 9868
rect 35624 9104 35676 9110
rect 35624 9046 35676 9052
rect 35348 8628 35400 8634
rect 35348 8570 35400 8576
rect 35452 8622 35572 8650
rect 35268 8498 35388 8514
rect 34520 8492 34572 8498
rect 35268 8492 35400 8498
rect 35268 8486 35348 8492
rect 34520 8434 34572 8440
rect 35348 8434 35400 8440
rect 34152 8424 34204 8430
rect 34152 8366 34204 8372
rect 34164 6866 34192 8366
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 35360 7970 35388 8434
rect 35452 8362 35480 8622
rect 35532 8560 35584 8566
rect 35532 8502 35584 8508
rect 35440 8356 35492 8362
rect 35440 8298 35492 8304
rect 35544 8090 35572 8502
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35176 7942 35388 7970
rect 35176 7886 35204 7942
rect 35636 7886 35664 9046
rect 36372 9042 36400 9862
rect 35900 9036 35952 9042
rect 35900 8978 35952 8984
rect 36360 9036 36412 9042
rect 36360 8978 36412 8984
rect 35912 8566 35940 8978
rect 35900 8560 35952 8566
rect 35900 8502 35952 8508
rect 35716 8356 35768 8362
rect 35716 8298 35768 8304
rect 35164 7880 35216 7886
rect 35164 7822 35216 7828
rect 35348 7880 35400 7886
rect 35348 7822 35400 7828
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 35176 7546 35204 7822
rect 35164 7540 35216 7546
rect 35164 7482 35216 7488
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34152 6860 34204 6866
rect 34152 6802 34204 6808
rect 34060 6792 34112 6798
rect 34060 6734 34112 6740
rect 34072 6458 34100 6734
rect 34060 6452 34112 6458
rect 34060 6394 34112 6400
rect 35360 6322 35388 7822
rect 35728 6866 35756 8298
rect 35900 7744 35952 7750
rect 35900 7686 35952 7692
rect 35912 6866 35940 7686
rect 36176 7200 36228 7206
rect 36176 7142 36228 7148
rect 35716 6860 35768 6866
rect 35716 6802 35768 6808
rect 35900 6860 35952 6866
rect 35900 6802 35952 6808
rect 35624 6792 35676 6798
rect 35624 6734 35676 6740
rect 35636 6458 35664 6734
rect 35624 6452 35676 6458
rect 35624 6394 35676 6400
rect 35912 6390 35940 6802
rect 36188 6730 36216 7142
rect 36176 6724 36228 6730
rect 36176 6666 36228 6672
rect 36452 6724 36504 6730
rect 36452 6666 36504 6672
rect 35992 6656 36044 6662
rect 35992 6598 36044 6604
rect 35900 6384 35952 6390
rect 35900 6326 35952 6332
rect 34796 6316 34848 6322
rect 34796 6258 34848 6264
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 34704 5024 34756 5030
rect 34704 4966 34756 4972
rect 34612 4684 34664 4690
rect 34612 4626 34664 4632
rect 34520 4480 34572 4486
rect 34520 4422 34572 4428
rect 34532 4146 34560 4422
rect 33876 4140 33928 4146
rect 33876 4082 33928 4088
rect 34520 4140 34572 4146
rect 34520 4082 34572 4088
rect 32496 3732 32548 3738
rect 32496 3674 32548 3680
rect 33888 3398 33916 4082
rect 34060 3936 34112 3942
rect 34060 3878 34112 3884
rect 33876 3392 33928 3398
rect 33876 3334 33928 3340
rect 34072 3126 34100 3878
rect 34624 3738 34652 4626
rect 34716 4078 34744 4966
rect 34808 4622 34836 6258
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35912 4826 35940 6326
rect 36004 6322 36032 6598
rect 36464 6458 36492 6666
rect 36452 6452 36504 6458
rect 36452 6394 36504 6400
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 35900 4820 35952 4826
rect 35900 4762 35952 4768
rect 37752 4758 37780 17614
rect 38016 14340 38068 14346
rect 38016 14282 38068 14288
rect 37924 14272 37976 14278
rect 37924 14214 37976 14220
rect 37830 8392 37886 8401
rect 37830 8327 37886 8336
rect 37844 6322 37872 8327
rect 37936 7449 37964 14214
rect 38028 13977 38056 14282
rect 38014 13968 38070 13977
rect 38014 13903 38070 13912
rect 38108 10056 38160 10062
rect 38108 9998 38160 10004
rect 38120 9897 38148 9998
rect 38106 9888 38162 9897
rect 38106 9823 38162 9832
rect 37922 7440 37978 7449
rect 37922 7375 37978 7384
rect 37832 6316 37884 6322
rect 37832 6258 37884 6264
rect 38016 6112 38068 6118
rect 38016 6054 38068 6060
rect 38028 5953 38056 6054
rect 38014 5944 38070 5953
rect 38014 5879 38070 5888
rect 37740 4752 37792 4758
rect 37740 4694 37792 4700
rect 34796 4616 34848 4622
rect 34796 4558 34848 4564
rect 34796 4480 34848 4486
rect 34796 4422 34848 4428
rect 35808 4480 35860 4486
rect 35808 4422 35860 4428
rect 36268 4480 36320 4486
rect 36268 4422 36320 4428
rect 34704 4072 34756 4078
rect 34704 4014 34756 4020
rect 34808 3890 34836 4422
rect 35440 4140 35492 4146
rect 35440 4082 35492 4088
rect 34716 3862 34836 3890
rect 34612 3732 34664 3738
rect 34612 3674 34664 3680
rect 31392 3120 31444 3126
rect 31392 3062 31444 3068
rect 34060 3120 34112 3126
rect 34060 3062 34112 3068
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 34624 2446 34652 3674
rect 34716 3466 34744 3862
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35452 3738 35480 4082
rect 35440 3732 35492 3738
rect 35440 3674 35492 3680
rect 35820 3534 35848 4422
rect 36280 3942 36308 4422
rect 36268 3936 36320 3942
rect 36268 3878 36320 3884
rect 36280 3602 36308 3878
rect 36268 3596 36320 3602
rect 36268 3538 36320 3544
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 34704 3460 34756 3466
rect 34704 3402 34756 3408
rect 34716 3194 34744 3402
rect 34704 3188 34756 3194
rect 34704 3130 34756 3136
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 38028 2009 38056 2246
rect 38014 2000 38070 2009
rect 38014 1935 38070 1944
rect 2778 368 2834 377
rect 2778 303 2834 312
<< via2 >>
rect 3422 39616 3478 39672
rect 1398 33496 1454 33552
rect 1398 32136 1454 32192
rect 1398 30812 1400 30832
rect 1400 30812 1452 30832
rect 1452 30812 1454 30832
rect 1398 30776 1454 30812
rect 1398 29416 1454 29472
rect 3238 28736 3294 28792
rect 1398 28092 1400 28112
rect 1400 28092 1452 28112
rect 1452 28092 1454 28112
rect 1398 28056 1454 28092
rect 1398 26696 1454 26752
rect 1398 25372 1400 25392
rect 1400 25372 1452 25392
rect 1452 25372 1454 25392
rect 1398 25336 1454 25372
rect 1398 23976 1454 24032
rect 3054 24692 3056 24712
rect 3056 24692 3108 24712
rect 3108 24692 3110 24712
rect 3054 24656 3110 24692
rect 3606 38936 3662 38992
rect 3698 38256 3754 38312
rect 3974 37576 4030 37632
rect 3790 36896 3846 36952
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4066 36216 4122 36272
rect 4066 35556 4122 35592
rect 4066 35536 4068 35556
rect 4068 35536 4120 35556
rect 4120 35536 4122 35556
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4066 34892 4068 34912
rect 4068 34892 4120 34912
rect 4120 34892 4122 34912
rect 4066 34856 4122 34892
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4066 34176 4122 34232
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 3238 23296 3294 23352
rect 1398 22652 1400 22672
rect 1400 22652 1452 22672
rect 1452 22652 1454 22672
rect 1398 22616 1454 22652
rect 1398 21256 1454 21312
rect 1398 19896 1454 19952
rect 1398 18536 1454 18592
rect 1398 17212 1400 17232
rect 1400 17212 1452 17232
rect 1452 17212 1454 17232
rect 1398 17176 1454 17212
rect 2870 19252 2872 19272
rect 2872 19252 2924 19272
rect 2924 19252 2926 19272
rect 2870 19216 2926 19252
rect 1398 15816 1454 15872
rect 1398 14456 1454 14512
rect 1398 13096 1454 13152
rect 4066 32816 4122 32872
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4158 31456 4214 31512
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 3882 30096 3938 30152
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 3974 27376 4030 27432
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4526 21936 4582 21992
rect 4526 21548 4582 21584
rect 4526 21528 4528 21548
rect 4528 21528 4580 21548
rect 4580 21528 4582 21548
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4066 20576 4122 20632
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4066 16496 4122 16552
rect 3974 15136 4030 15192
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 3882 13776 3938 13832
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 1398 11772 1400 11792
rect 1400 11772 1452 11792
rect 1452 11772 1454 11792
rect 1398 11736 1454 11772
rect 1398 10376 1454 10432
rect 1398 9052 1400 9072
rect 1400 9052 1452 9072
rect 1452 9052 1454 9072
rect 1398 9016 1454 9052
rect 3514 12416 3570 12472
rect 1398 7656 1454 7712
rect 1398 6296 1454 6352
rect 1398 4936 1454 4992
rect 1398 3576 1454 3632
rect 2686 2216 2742 2272
rect 1858 1536 1914 1592
rect 1398 856 1454 912
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4066 11076 4122 11112
rect 4066 11056 4068 11076
rect 4068 11056 4120 11076
rect 4120 11056 4122 11076
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4066 9716 4122 9752
rect 4066 9696 4068 9716
rect 4068 9696 4120 9716
rect 4120 9696 4122 9716
rect 5630 26016 5686 26072
rect 7102 21800 7158 21856
rect 5538 17740 5594 17776
rect 5538 17720 5540 17740
rect 5540 17720 5592 17740
rect 5592 17720 5594 17740
rect 38014 37848 38070 37904
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 14462 34468 14518 34504
rect 14462 34448 14464 34468
rect 14464 34448 14516 34468
rect 14516 34448 14518 34468
rect 14646 33224 14702 33280
rect 10598 21936 10654 21992
rect 12898 21800 12954 21856
rect 12622 21528 12678 21584
rect 9770 12824 9826 12880
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4066 8356 4122 8392
rect 4066 8336 4068 8356
rect 4068 8336 4120 8356
rect 4120 8336 4122 8356
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4066 6976 4122 7032
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4066 5616 4122 5672
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 5722 4564 5724 4584
rect 5724 4564 5776 4584
rect 5776 4564 5778 4584
rect 5722 4528 5778 4564
rect 4066 4256 4122 4312
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 11058 9968 11114 10024
rect 17682 34584 17738 34640
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 17958 33224 18014 33280
rect 18602 34584 18658 34640
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 18418 34468 18474 34504
rect 18418 34448 18420 34468
rect 18420 34448 18472 34468
rect 18472 34448 18474 34468
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 9494 6296 9550 6352
rect 10506 4800 10562 4856
rect 12438 4800 12494 4856
rect 11610 4120 11666 4176
rect 3974 2896 4030 2952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 15566 7404 15622 7440
rect 15566 7384 15568 7404
rect 15568 7384 15620 7404
rect 15620 7384 15622 7404
rect 14186 4528 14242 4584
rect 16578 7248 16634 7304
rect 16578 4120 16634 4176
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19338 9968 19394 10024
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 27066 21936 27122 21992
rect 23478 12824 23534 12880
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 20258 6840 20314 6896
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 23938 6316 23994 6352
rect 23938 6296 23940 6316
rect 23940 6296 23992 6316
rect 23992 6296 23994 6316
rect 20074 4800 20130 4856
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 25318 6840 25374 6896
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 28446 6976 28502 7032
rect 29182 6976 29238 7032
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 38106 33940 38108 33960
rect 38108 33940 38160 33960
rect 38160 33940 38162 33960
rect 38106 33904 38162 33940
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 31666 8336 31722 8392
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 38106 29824 38162 29880
rect 38014 25880 38070 25936
rect 38014 21936 38070 21992
rect 38014 17876 38070 17912
rect 38014 17856 38016 17876
rect 38016 17856 38068 17876
rect 38068 17856 38070 17876
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 37830 8336 37886 8392
rect 38014 13912 38070 13968
rect 38106 9832 38162 9888
rect 37922 7384 37978 7440
rect 38014 5888 38070 5944
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 38014 1944 38070 2000
rect 2778 312 2834 368
<< metal3 >>
rect 0 39674 800 39704
rect 3417 39674 3483 39677
rect 0 39672 3483 39674
rect 0 39616 3422 39672
rect 3478 39616 3483 39672
rect 0 39614 3483 39616
rect 0 39584 800 39614
rect 3417 39611 3483 39614
rect 0 38994 800 39024
rect 3601 38994 3667 38997
rect 0 38992 3667 38994
rect 0 38936 3606 38992
rect 3662 38936 3667 38992
rect 0 38934 3667 38936
rect 0 38904 800 38934
rect 3601 38931 3667 38934
rect 0 38314 800 38344
rect 3693 38314 3759 38317
rect 0 38312 3759 38314
rect 0 38256 3698 38312
rect 3754 38256 3759 38312
rect 0 38254 3759 38256
rect 0 38224 800 38254
rect 3693 38251 3759 38254
rect 38009 37906 38075 37909
rect 39200 37906 40000 37936
rect 38009 37904 40000 37906
rect 38009 37848 38014 37904
rect 38070 37848 40000 37904
rect 38009 37846 40000 37848
rect 38009 37843 38075 37846
rect 39200 37816 40000 37846
rect 0 37634 800 37664
rect 3969 37634 4035 37637
rect 0 37632 4035 37634
rect 0 37576 3974 37632
rect 4030 37576 4035 37632
rect 0 37574 4035 37576
rect 0 37544 800 37574
rect 3969 37571 4035 37574
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 19568 37024 19888 37025
rect 0 36954 800 36984
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 3785 36954 3851 36957
rect 0 36952 3851 36954
rect 0 36896 3790 36952
rect 3846 36896 3851 36952
rect 0 36894 3851 36896
rect 0 36864 800 36894
rect 3785 36891 3851 36894
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36274 800 36304
rect 4061 36274 4127 36277
rect 0 36272 4127 36274
rect 0 36216 4066 36272
rect 4122 36216 4127 36272
rect 0 36214 4127 36216
rect 0 36184 800 36214
rect 4061 36211 4127 36214
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35594 800 35624
rect 4061 35594 4127 35597
rect 0 35592 4127 35594
rect 0 35536 4066 35592
rect 4122 35536 4127 35592
rect 0 35534 4127 35536
rect 0 35504 800 35534
rect 4061 35531 4127 35534
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34914 800 34944
rect 4061 34914 4127 34917
rect 0 34912 4127 34914
rect 0 34856 4066 34912
rect 4122 34856 4127 34912
rect 0 34854 4127 34856
rect 0 34824 800 34854
rect 4061 34851 4127 34854
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 17677 34642 17743 34645
rect 18597 34642 18663 34645
rect 17677 34640 18663 34642
rect 17677 34584 17682 34640
rect 17738 34584 18602 34640
rect 18658 34584 18663 34640
rect 17677 34582 18663 34584
rect 17677 34579 17743 34582
rect 18597 34579 18663 34582
rect 14457 34506 14523 34509
rect 18413 34506 18479 34509
rect 14457 34504 18479 34506
rect 14457 34448 14462 34504
rect 14518 34448 18418 34504
rect 18474 34448 18479 34504
rect 14457 34446 18479 34448
rect 14457 34443 14523 34446
rect 18413 34443 18479 34446
rect 4208 34304 4528 34305
rect 0 34234 800 34264
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 4061 34234 4127 34237
rect 0 34232 4127 34234
rect 0 34176 4066 34232
rect 4122 34176 4127 34232
rect 0 34174 4127 34176
rect 0 34144 800 34174
rect 4061 34171 4127 34174
rect 38101 33962 38167 33965
rect 39200 33962 40000 33992
rect 38101 33960 40000 33962
rect 38101 33904 38106 33960
rect 38162 33904 40000 33960
rect 38101 33902 40000 33904
rect 38101 33899 38167 33902
rect 39200 33872 40000 33902
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33554 800 33584
rect 1393 33554 1459 33557
rect 0 33552 1459 33554
rect 0 33496 1398 33552
rect 1454 33496 1459 33552
rect 0 33494 1459 33496
rect 0 33464 800 33494
rect 1393 33491 1459 33494
rect 14641 33282 14707 33285
rect 17953 33282 18019 33285
rect 14641 33280 18019 33282
rect 14641 33224 14646 33280
rect 14702 33224 17958 33280
rect 18014 33224 18019 33280
rect 14641 33222 18019 33224
rect 14641 33219 14707 33222
rect 17953 33219 18019 33222
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32874 800 32904
rect 4061 32874 4127 32877
rect 0 32872 4127 32874
rect 0 32816 4066 32872
rect 4122 32816 4127 32872
rect 0 32814 4127 32816
rect 0 32784 800 32814
rect 4061 32811 4127 32814
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 0 32194 800 32224
rect 1393 32194 1459 32197
rect 0 32192 1459 32194
rect 0 32136 1398 32192
rect 1454 32136 1459 32192
rect 0 32134 1459 32136
rect 0 32104 800 32134
rect 1393 32131 1459 32134
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 0 31514 800 31544
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 4153 31514 4219 31517
rect 0 31512 4219 31514
rect 0 31456 4158 31512
rect 4214 31456 4219 31512
rect 0 31454 4219 31456
rect 0 31424 800 31454
rect 4153 31451 4219 31454
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30834 800 30864
rect 1393 30834 1459 30837
rect 0 30832 1459 30834
rect 0 30776 1398 30832
rect 1454 30776 1459 30832
rect 0 30774 1459 30776
rect 0 30744 800 30774
rect 1393 30771 1459 30774
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 30154 800 30184
rect 3877 30154 3943 30157
rect 0 30152 3943 30154
rect 0 30096 3882 30152
rect 3938 30096 3943 30152
rect 0 30094 3943 30096
rect 0 30064 800 30094
rect 3877 30091 3943 30094
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 38101 29882 38167 29885
rect 39200 29882 40000 29912
rect 38101 29880 40000 29882
rect 38101 29824 38106 29880
rect 38162 29824 40000 29880
rect 38101 29822 40000 29824
rect 38101 29819 38167 29822
rect 39200 29792 40000 29822
rect 0 29474 800 29504
rect 1393 29474 1459 29477
rect 0 29472 1459 29474
rect 0 29416 1398 29472
rect 1454 29416 1459 29472
rect 0 29414 1459 29416
rect 0 29384 800 29414
rect 1393 29411 1459 29414
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 4208 28864 4528 28865
rect 0 28794 800 28824
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 3233 28794 3299 28797
rect 0 28792 3299 28794
rect 0 28736 3238 28792
rect 3294 28736 3299 28792
rect 0 28734 3299 28736
rect 0 28704 800 28734
rect 3233 28731 3299 28734
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 28114 800 28144
rect 1393 28114 1459 28117
rect 0 28112 1459 28114
rect 0 28056 1398 28112
rect 1454 28056 1459 28112
rect 0 28054 1459 28056
rect 0 28024 800 28054
rect 1393 28051 1459 28054
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27434 800 27464
rect 3969 27434 4035 27437
rect 0 27432 4035 27434
rect 0 27376 3974 27432
rect 4030 27376 4035 27432
rect 0 27374 4035 27376
rect 0 27344 800 27374
rect 3969 27371 4035 27374
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 0 26754 800 26784
rect 1393 26754 1459 26757
rect 0 26752 1459 26754
rect 0 26696 1398 26752
rect 1454 26696 1459 26752
rect 0 26694 1459 26696
rect 0 26664 800 26694
rect 1393 26691 1459 26694
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 19568 26144 19888 26145
rect 0 26074 800 26104
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 5625 26074 5691 26077
rect 0 26072 5691 26074
rect 0 26016 5630 26072
rect 5686 26016 5691 26072
rect 0 26014 5691 26016
rect 0 25984 800 26014
rect 5625 26011 5691 26014
rect 38009 25938 38075 25941
rect 39200 25938 40000 25968
rect 38009 25936 40000 25938
rect 38009 25880 38014 25936
rect 38070 25880 40000 25936
rect 38009 25878 40000 25880
rect 38009 25875 38075 25878
rect 39200 25848 40000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25394 800 25424
rect 1393 25394 1459 25397
rect 0 25392 1459 25394
rect 0 25336 1398 25392
rect 1454 25336 1459 25392
rect 0 25334 1459 25336
rect 0 25304 800 25334
rect 1393 25331 1459 25334
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24714 800 24744
rect 3049 24714 3115 24717
rect 0 24712 3115 24714
rect 0 24656 3054 24712
rect 3110 24656 3115 24712
rect 0 24654 3115 24656
rect 0 24624 800 24654
rect 3049 24651 3115 24654
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 0 24034 800 24064
rect 1393 24034 1459 24037
rect 0 24032 1459 24034
rect 0 23976 1398 24032
rect 1454 23976 1459 24032
rect 0 23974 1459 23976
rect 0 23944 800 23974
rect 1393 23971 1459 23974
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 4208 23424 4528 23425
rect 0 23354 800 23384
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 3233 23354 3299 23357
rect 0 23352 3299 23354
rect 0 23296 3238 23352
rect 3294 23296 3299 23352
rect 0 23294 3299 23296
rect 0 23264 800 23294
rect 3233 23291 3299 23294
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22674 800 22704
rect 1393 22674 1459 22677
rect 0 22672 1459 22674
rect 0 22616 1398 22672
rect 1454 22616 1459 22672
rect 0 22614 1459 22616
rect 0 22584 800 22614
rect 1393 22611 1459 22614
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21994 800 22024
rect 4521 21994 4587 21997
rect 0 21992 4587 21994
rect 0 21936 4526 21992
rect 4582 21936 4587 21992
rect 0 21934 4587 21936
rect 0 21904 800 21934
rect 4521 21931 4587 21934
rect 10593 21994 10659 21997
rect 27061 21994 27127 21997
rect 10593 21992 27127 21994
rect 10593 21936 10598 21992
rect 10654 21936 27066 21992
rect 27122 21936 27127 21992
rect 10593 21934 27127 21936
rect 10593 21931 10659 21934
rect 27061 21931 27127 21934
rect 38009 21994 38075 21997
rect 39200 21994 40000 22024
rect 38009 21992 40000 21994
rect 38009 21936 38014 21992
rect 38070 21936 40000 21992
rect 38009 21934 40000 21936
rect 38009 21931 38075 21934
rect 39200 21904 40000 21934
rect 7097 21858 7163 21861
rect 12893 21858 12959 21861
rect 7097 21856 12959 21858
rect 7097 21800 7102 21856
rect 7158 21800 12898 21856
rect 12954 21800 12959 21856
rect 7097 21798 12959 21800
rect 7097 21795 7163 21798
rect 12893 21795 12959 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 4521 21586 4587 21589
rect 12617 21586 12683 21589
rect 4521 21584 12683 21586
rect 4521 21528 4526 21584
rect 4582 21528 12622 21584
rect 12678 21528 12683 21584
rect 4521 21526 12683 21528
rect 4521 21523 4587 21526
rect 12617 21523 12683 21526
rect 0 21314 800 21344
rect 1393 21314 1459 21317
rect 0 21312 1459 21314
rect 0 21256 1398 21312
rect 1454 21256 1459 21312
rect 0 21254 1459 21256
rect 0 21224 800 21254
rect 1393 21251 1459 21254
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 19568 20704 19888 20705
rect 0 20634 800 20664
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 4061 20634 4127 20637
rect 0 20632 4127 20634
rect 0 20576 4066 20632
rect 4122 20576 4127 20632
rect 0 20574 4127 20576
rect 0 20544 800 20574
rect 4061 20571 4127 20574
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19954 800 19984
rect 1393 19954 1459 19957
rect 0 19952 1459 19954
rect 0 19896 1398 19952
rect 1454 19896 1459 19952
rect 0 19894 1459 19896
rect 0 19864 800 19894
rect 1393 19891 1459 19894
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19274 800 19304
rect 2865 19274 2931 19277
rect 0 19272 2931 19274
rect 0 19216 2870 19272
rect 2926 19216 2931 19272
rect 0 19214 2931 19216
rect 0 19184 800 19214
rect 2865 19211 2931 19214
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 0 18594 800 18624
rect 1393 18594 1459 18597
rect 0 18592 1459 18594
rect 0 18536 1398 18592
rect 1454 18536 1459 18592
rect 0 18534 1459 18536
rect 0 18504 800 18534
rect 1393 18531 1459 18534
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 4208 17984 4528 17985
rect 0 17914 800 17944
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 38009 17914 38075 17917
rect 39200 17914 40000 17944
rect 0 17854 4124 17914
rect 0 17824 800 17854
rect 4064 17778 4124 17854
rect 38009 17912 40000 17914
rect 38009 17856 38014 17912
rect 38070 17856 40000 17912
rect 38009 17854 40000 17856
rect 38009 17851 38075 17854
rect 39200 17824 40000 17854
rect 5533 17778 5599 17781
rect 4064 17776 5599 17778
rect 4064 17720 5538 17776
rect 5594 17720 5599 17776
rect 4064 17718 5599 17720
rect 5533 17715 5599 17718
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17234 800 17264
rect 1393 17234 1459 17237
rect 0 17232 1459 17234
rect 0 17176 1398 17232
rect 1454 17176 1459 17232
rect 0 17174 1459 17176
rect 0 17144 800 17174
rect 1393 17171 1459 17174
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16554 800 16584
rect 4061 16554 4127 16557
rect 0 16552 4127 16554
rect 0 16496 4066 16552
rect 4122 16496 4127 16552
rect 0 16494 4127 16496
rect 0 16464 800 16494
rect 4061 16491 4127 16494
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 0 15874 800 15904
rect 1393 15874 1459 15877
rect 0 15872 1459 15874
rect 0 15816 1398 15872
rect 1454 15816 1459 15872
rect 0 15814 1459 15816
rect 0 15784 800 15814
rect 1393 15811 1459 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 19568 15264 19888 15265
rect 0 15194 800 15224
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 3969 15194 4035 15197
rect 0 15192 4035 15194
rect 0 15136 3974 15192
rect 4030 15136 4035 15192
rect 0 15134 4035 15136
rect 0 15104 800 15134
rect 3969 15131 4035 15134
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14514 800 14544
rect 1393 14514 1459 14517
rect 0 14512 1459 14514
rect 0 14456 1398 14512
rect 1454 14456 1459 14512
rect 0 14454 1459 14456
rect 0 14424 800 14454
rect 1393 14451 1459 14454
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 38009 13970 38075 13973
rect 39200 13970 40000 14000
rect 38009 13968 40000 13970
rect 38009 13912 38014 13968
rect 38070 13912 40000 13968
rect 38009 13910 40000 13912
rect 38009 13907 38075 13910
rect 39200 13880 40000 13910
rect 0 13834 800 13864
rect 3877 13834 3943 13837
rect 0 13832 3943 13834
rect 0 13776 3882 13832
rect 3938 13776 3943 13832
rect 0 13774 3943 13776
rect 0 13744 800 13774
rect 3877 13771 3943 13774
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 0 13154 800 13184
rect 1393 13154 1459 13157
rect 0 13152 1459 13154
rect 0 13096 1398 13152
rect 1454 13096 1459 13152
rect 0 13094 1459 13096
rect 0 13064 800 13094
rect 1393 13091 1459 13094
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 9765 12882 9831 12885
rect 23473 12882 23539 12885
rect 9765 12880 23539 12882
rect 9765 12824 9770 12880
rect 9826 12824 23478 12880
rect 23534 12824 23539 12880
rect 9765 12822 23539 12824
rect 9765 12819 9831 12822
rect 23473 12819 23539 12822
rect 4208 12544 4528 12545
rect 0 12474 800 12504
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 3509 12474 3575 12477
rect 0 12472 3575 12474
rect 0 12416 3514 12472
rect 3570 12416 3575 12472
rect 0 12414 3575 12416
rect 0 12384 800 12414
rect 3509 12411 3575 12414
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11794 800 11824
rect 1393 11794 1459 11797
rect 0 11792 1459 11794
rect 0 11736 1398 11792
rect 1454 11736 1459 11792
rect 0 11734 1459 11736
rect 0 11704 800 11734
rect 1393 11731 1459 11734
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 11114 800 11144
rect 4061 11114 4127 11117
rect 0 11112 4127 11114
rect 0 11056 4066 11112
rect 4122 11056 4127 11112
rect 0 11054 4127 11056
rect 0 11024 800 11054
rect 4061 11051 4127 11054
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 11053 10026 11119 10029
rect 19333 10026 19399 10029
rect 11053 10024 19399 10026
rect 11053 9968 11058 10024
rect 11114 9968 19338 10024
rect 19394 9968 19399 10024
rect 11053 9966 19399 9968
rect 11053 9963 11119 9966
rect 19333 9963 19399 9966
rect 38101 9890 38167 9893
rect 39200 9890 40000 9920
rect 38101 9888 40000 9890
rect 38101 9832 38106 9888
rect 38162 9832 40000 9888
rect 38101 9830 40000 9832
rect 38101 9827 38167 9830
rect 19568 9824 19888 9825
rect 0 9754 800 9784
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 39200 9800 40000 9830
rect 19568 9759 19888 9760
rect 4061 9754 4127 9757
rect 0 9752 4127 9754
rect 0 9696 4066 9752
rect 4122 9696 4127 9752
rect 0 9694 4127 9696
rect 0 9664 800 9694
rect 4061 9691 4127 9694
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 9074 800 9104
rect 1393 9074 1459 9077
rect 0 9072 1459 9074
rect 0 9016 1398 9072
rect 1454 9016 1459 9072
rect 0 9014 1459 9016
rect 0 8984 800 9014
rect 1393 9011 1459 9014
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8394 800 8424
rect 4061 8394 4127 8397
rect 0 8392 4127 8394
rect 0 8336 4066 8392
rect 4122 8336 4127 8392
rect 0 8334 4127 8336
rect 0 8304 800 8334
rect 4061 8331 4127 8334
rect 31661 8394 31727 8397
rect 37825 8394 37891 8397
rect 31661 8392 37891 8394
rect 31661 8336 31666 8392
rect 31722 8336 37830 8392
rect 37886 8336 37891 8392
rect 31661 8334 37891 8336
rect 31661 8331 31727 8334
rect 37825 8331 37891 8334
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 0 7714 800 7744
rect 1393 7714 1459 7717
rect 0 7712 1459 7714
rect 0 7656 1398 7712
rect 1454 7656 1459 7712
rect 0 7654 1459 7656
rect 0 7624 800 7654
rect 1393 7651 1459 7654
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 15561 7442 15627 7445
rect 37917 7442 37983 7445
rect 15561 7440 37983 7442
rect 15561 7384 15566 7440
rect 15622 7384 37922 7440
rect 37978 7384 37983 7440
rect 15561 7382 37983 7384
rect 15561 7379 15627 7382
rect 37917 7379 37983 7382
rect 16573 7306 16639 7309
rect 16573 7304 26250 7306
rect 16573 7248 16578 7304
rect 16634 7248 26250 7304
rect 16573 7246 26250 7248
rect 16573 7243 16639 7246
rect 4208 7104 4528 7105
rect 0 7034 800 7064
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 4061 7034 4127 7037
rect 0 7032 4127 7034
rect 0 6976 4066 7032
rect 4122 6976 4127 7032
rect 0 6974 4127 6976
rect 26190 7034 26250 7246
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 28441 7034 28507 7037
rect 29177 7034 29243 7037
rect 26190 7032 29243 7034
rect 26190 6976 28446 7032
rect 28502 6976 29182 7032
rect 29238 6976 29243 7032
rect 26190 6974 29243 6976
rect 0 6944 800 6974
rect 4061 6971 4127 6974
rect 28441 6971 28507 6974
rect 29177 6971 29243 6974
rect 20253 6898 20319 6901
rect 25313 6898 25379 6901
rect 20253 6896 25379 6898
rect 20253 6840 20258 6896
rect 20314 6840 25318 6896
rect 25374 6840 25379 6896
rect 20253 6838 25379 6840
rect 20253 6835 20319 6838
rect 25313 6835 25379 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6354 800 6384
rect 1393 6354 1459 6357
rect 0 6352 1459 6354
rect 0 6296 1398 6352
rect 1454 6296 1459 6352
rect 0 6294 1459 6296
rect 0 6264 800 6294
rect 1393 6291 1459 6294
rect 9489 6354 9555 6357
rect 23933 6354 23999 6357
rect 9489 6352 23999 6354
rect 9489 6296 9494 6352
rect 9550 6296 23938 6352
rect 23994 6296 23999 6352
rect 9489 6294 23999 6296
rect 9489 6291 9555 6294
rect 23933 6291 23999 6294
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 38009 5946 38075 5949
rect 39200 5946 40000 5976
rect 38009 5944 40000 5946
rect 38009 5888 38014 5944
rect 38070 5888 40000 5944
rect 38009 5886 40000 5888
rect 38009 5883 38075 5886
rect 39200 5856 40000 5886
rect 0 5674 800 5704
rect 4061 5674 4127 5677
rect 0 5672 4127 5674
rect 0 5616 4066 5672
rect 4122 5616 4127 5672
rect 0 5614 4127 5616
rect 0 5584 800 5614
rect 4061 5611 4127 5614
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4994 800 5024
rect 1393 4994 1459 4997
rect 0 4992 1459 4994
rect 0 4936 1398 4992
rect 1454 4936 1459 4992
rect 0 4934 1459 4936
rect 0 4904 800 4934
rect 1393 4931 1459 4934
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 10501 4858 10567 4861
rect 12433 4858 12499 4861
rect 20069 4858 20135 4861
rect 10501 4856 20135 4858
rect 10501 4800 10506 4856
rect 10562 4800 12438 4856
rect 12494 4800 20074 4856
rect 20130 4800 20135 4856
rect 10501 4798 20135 4800
rect 10501 4795 10567 4798
rect 12433 4795 12499 4798
rect 20069 4795 20135 4798
rect 5717 4586 5783 4589
rect 14181 4586 14247 4589
rect 5717 4584 14247 4586
rect 5717 4528 5722 4584
rect 5778 4528 14186 4584
rect 14242 4528 14247 4584
rect 5717 4526 14247 4528
rect 5717 4523 5783 4526
rect 14181 4523 14247 4526
rect 19568 4384 19888 4385
rect 0 4314 800 4344
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 4061 4314 4127 4317
rect 0 4312 4127 4314
rect 0 4256 4066 4312
rect 4122 4256 4127 4312
rect 0 4254 4127 4256
rect 0 4224 800 4254
rect 4061 4251 4127 4254
rect 11605 4178 11671 4181
rect 16573 4178 16639 4181
rect 11605 4176 16639 4178
rect 11605 4120 11610 4176
rect 11666 4120 16578 4176
rect 16634 4120 16639 4176
rect 11605 4118 16639 4120
rect 11605 4115 11671 4118
rect 16573 4115 16639 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3634 800 3664
rect 1393 3634 1459 3637
rect 0 3632 1459 3634
rect 0 3576 1398 3632
rect 1454 3576 1459 3632
rect 0 3574 1459 3576
rect 0 3544 800 3574
rect 1393 3571 1459 3574
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 0 2954 800 2984
rect 3969 2954 4035 2957
rect 0 2952 4035 2954
rect 0 2896 3974 2952
rect 4030 2896 4035 2952
rect 0 2894 4035 2896
rect 0 2864 800 2894
rect 3969 2891 4035 2894
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 0 2274 800 2304
rect 2681 2274 2747 2277
rect 0 2272 2747 2274
rect 0 2216 2686 2272
rect 2742 2216 2747 2272
rect 0 2214 2747 2216
rect 0 2184 800 2214
rect 2681 2211 2747 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 38009 2002 38075 2005
rect 39200 2002 40000 2032
rect 38009 2000 40000 2002
rect 38009 1944 38014 2000
rect 38070 1944 40000 2000
rect 38009 1942 40000 1944
rect 38009 1939 38075 1942
rect 39200 1912 40000 1942
rect 0 1594 800 1624
rect 1853 1594 1919 1597
rect 0 1592 1919 1594
rect 0 1536 1858 1592
rect 1914 1536 1919 1592
rect 0 1534 1919 1536
rect 0 1504 800 1534
rect 1853 1531 1919 1534
rect 0 914 800 944
rect 1393 914 1459 917
rect 0 912 1459 914
rect 0 856 1398 912
rect 1454 856 1459 912
rect 0 854 1459 856
rect 0 824 800 854
rect 1393 851 1459 854
rect 0 370 800 400
rect 2773 370 2839 373
rect 0 368 2839 370
rect 0 312 2778 368
rect 2834 312 2839 368
rect 0 310 2839 312
rect 0 280 800 310
rect 2773 307 2839 310
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12420 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A
timestamp 1644511149
transform 1 0 12972 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1644511149
transform 1 0 17480 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A
timestamp 1644511149
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__D
timestamp 1644511149
transform 1 0 17204 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1644511149
transform 1 0 17848 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1644511149
transform 1 0 17480 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1644511149
transform -1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__D
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A
timestamp 1644511149
transform 1 0 17940 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__D
timestamp 1644511149
transform -1 0 18492 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__D
timestamp 1644511149
transform 1 0 17020 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A
timestamp 1644511149
transform -1 0 16744 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__D
timestamp 1644511149
transform -1 0 15272 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1644511149
transform -1 0 16928 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A
timestamp 1644511149
transform 1 0 10856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1644511149
transform 1 0 10856 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A
timestamp 1644511149
transform -1 0 15548 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A
timestamp 1644511149
transform 1 0 11592 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1644511149
transform 1 0 19320 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1644511149
transform -1 0 20884 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__C
timestamp 1644511149
transform 1 0 22264 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__D
timestamp 1644511149
transform 1 0 22448 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A
timestamp 1644511149
transform -1 0 19412 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__D
timestamp 1644511149
transform 1 0 22908 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A
timestamp 1644511149
transform 1 0 19688 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__D
timestamp 1644511149
transform -1 0 20424 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A
timestamp 1644511149
transform 1 0 15456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__C
timestamp 1644511149
transform 1 0 16008 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__D
timestamp 1644511149
transform -1 0 19596 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__D
timestamp 1644511149
transform 1 0 19780 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A
timestamp 1644511149
transform 1 0 13064 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1644511149
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__D
timestamp 1644511149
transform 1 0 18584 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A
timestamp 1644511149
transform 1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__C
timestamp 1644511149
transform -1 0 17848 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__D
timestamp 1644511149
transform -1 0 19320 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__C
timestamp 1644511149
transform 1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1644511149
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1644511149
transform -1 0 20240 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__D
timestamp 1644511149
transform -1 0 22172 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__C
timestamp 1644511149
transform 1 0 15824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__D
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__C
timestamp 1644511149
transform 1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1644511149
transform -1 0 11868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1644511149
transform 1 0 12420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1644511149
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1644511149
transform 1 0 6992 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A
timestamp 1644511149
transform 1 0 8832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A
timestamp 1644511149
transform 1 0 7544 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A
timestamp 1644511149
transform 1 0 8280 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1644511149
transform 1 0 4048 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__C
timestamp 1644511149
transform -1 0 8464 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__C
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__D
timestamp 1644511149
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1644511149
transform 1 0 27048 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A
timestamp 1644511149
transform -1 0 25208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1644511149
transform -1 0 24196 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__C
timestamp 1644511149
transform 1 0 24840 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__D
timestamp 1644511149
transform -1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__C
timestamp 1644511149
transform 1 0 26312 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__D
timestamp 1644511149
transform -1 0 25944 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__C
timestamp 1644511149
transform -1 0 26496 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__D
timestamp 1644511149
transform -1 0 26128 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__C
timestamp 1644511149
transform 1 0 25852 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__D
timestamp 1644511149
transform 1 0 25208 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__C
timestamp 1644511149
transform -1 0 26772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__D
timestamp 1644511149
transform -1 0 27784 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1644511149
transform -1 0 7636 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1644511149
transform 1 0 8004 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__C
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__D
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__C
timestamp 1644511149
transform -1 0 8372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__D
timestamp 1644511149
transform -1 0 7912 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__C
timestamp 1644511149
transform 1 0 6532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1644511149
transform 1 0 6624 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A
timestamp 1644511149
transform 1 0 5704 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A
timestamp 1644511149
transform -1 0 6256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1644511149
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1644511149
transform 1 0 13340 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A
timestamp 1644511149
transform -1 0 14720 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A
timestamp 1644511149
transform -1 0 14260 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__D
timestamp 1644511149
transform 1 0 11684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__D
timestamp 1644511149
transform 1 0 10856 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__D
timestamp 1644511149
transform 1 0 25300 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__D
timestamp 1644511149
transform -1 0 23920 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__D
timestamp 1644511149
transform -1 0 25576 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1644511149
transform 1 0 19504 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A
timestamp 1644511149
transform 1 0 23184 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1644511149
transform 1 0 22172 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__C
timestamp 1644511149
transform 1 0 23644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__C
timestamp 1644511149
transform -1 0 25484 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A
timestamp 1644511149
transform -1 0 21344 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1644511149
transform 1 0 13892 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1644511149
transform -1 0 12144 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__A
timestamp 1644511149
transform -1 0 20884 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A
timestamp 1644511149
transform -1 0 31464 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A
timestamp 1644511149
transform -1 0 32844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1644511149
transform 1 0 12052 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__B
timestamp 1644511149
transform 1 0 13340 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1644511149
transform 1 0 20792 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__B
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__C
timestamp 1644511149
transform 1 0 18124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1644511149
transform 1 0 31004 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A
timestamp 1644511149
transform 1 0 25944 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__B2
timestamp 1644511149
transform -1 0 33580 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A
timestamp 1644511149
transform 1 0 32936 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1644511149
transform -1 0 31648 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__A1
timestamp 1644511149
transform -1 0 29900 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A1
timestamp 1644511149
transform -1 0 28060 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__A1
timestamp 1644511149
transform 1 0 28520 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A1
timestamp 1644511149
transform 1 0 30452 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A2
timestamp 1644511149
transform -1 0 30912 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A1
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A2
timestamp 1644511149
transform 1 0 32292 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A
timestamp 1644511149
transform 1 0 31280 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A0
timestamp 1644511149
transform 1 0 34776 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A1
timestamp 1644511149
transform -1 0 32200 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A2
timestamp 1644511149
transform 1 0 31464 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__A
timestamp 1644511149
transform 1 0 23828 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A0
timestamp 1644511149
transform 1 0 36064 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1
timestamp 1644511149
transform 1 0 32476 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A2
timestamp 1644511149
transform 1 0 33028 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A1
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A0
timestamp 1644511149
transform 1 0 29808 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A1
timestamp 1644511149
transform -1 0 34040 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A
timestamp 1644511149
transform 1 0 29716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A0
timestamp 1644511149
transform 1 0 29900 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A0
timestamp 1644511149
transform 1 0 28888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A
timestamp 1644511149
transform 1 0 30728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A0
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__S
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A
timestamp 1644511149
transform 1 0 30452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A0
timestamp 1644511149
transform 1 0 27784 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A
timestamp 1644511149
transform 1 0 28336 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A0
timestamp 1644511149
transform 1 0 29440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__A
timestamp 1644511149
transform -1 0 29716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__A0
timestamp 1644511149
transform 1 0 28980 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__S
timestamp 1644511149
transform -1 0 30636 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__A
timestamp 1644511149
transform -1 0 29808 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A0
timestamp 1644511149
transform 1 0 26036 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__S
timestamp 1644511149
transform -1 0 26404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A0
timestamp 1644511149
transform 1 0 28888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A
timestamp 1644511149
transform 1 0 28428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__C1
timestamp 1644511149
transform 1 0 35236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A
timestamp 1644511149
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A1
timestamp 1644511149
transform 1 0 15732 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A
timestamp 1644511149
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__B
timestamp 1644511149
transform -1 0 17112 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__C
timestamp 1644511149
transform 1 0 17296 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B2
timestamp 1644511149
transform 1 0 15088 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A
timestamp 1644511149
transform -1 0 14720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A
timestamp 1644511149
transform -1 0 20516 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A1
timestamp 1644511149
transform -1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B2
timestamp 1644511149
transform 1 0 12328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A
timestamp 1644511149
transform -1 0 12236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A1
timestamp 1644511149
transform -1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B2
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A1
timestamp 1644511149
transform 1 0 5428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__B2
timestamp 1644511149
transform 1 0 6532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A
timestamp 1644511149
transform 1 0 4600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A1
timestamp 1644511149
transform 1 0 5152 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__B2
timestamp 1644511149
transform 1 0 5704 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A
timestamp 1644511149
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__A1
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A
timestamp 1644511149
transform -1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A1
timestamp 1644511149
transform -1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__A0
timestamp 1644511149
transform -1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A1
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__A0
timestamp 1644511149
transform 1 0 20884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A0
timestamp 1644511149
transform 1 0 20056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A1
timestamp 1644511149
transform -1 0 20792 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__B
timestamp 1644511149
transform 1 0 15364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A0
timestamp 1644511149
transform -1 0 26496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A0
timestamp 1644511149
transform 1 0 28428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__A0
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A0
timestamp 1644511149
transform 1 0 23736 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A0
timestamp 1644511149
transform -1 0 29992 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__A
timestamp 1644511149
transform -1 0 31188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A0
timestamp 1644511149
transform -1 0 20148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A0
timestamp 1644511149
transform 1 0 26496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A0
timestamp 1644511149
transform 1 0 28888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__A
timestamp 1644511149
transform 1 0 30268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__C1
timestamp 1644511149
transform -1 0 35420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__C
timestamp 1644511149
transform -1 0 32936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__B1
timestamp 1644511149
transform 1 0 33948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__A
timestamp 1644511149
transform -1 0 34132 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__B1
timestamp 1644511149
transform 1 0 33488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__CLK
timestamp 1644511149
transform -1 0 35144 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1366__CLK
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__CLK
timestamp 1644511149
transform 1 0 32936 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__CLK
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__CLK
timestamp 1644511149
transform 1 0 32936 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__CLK
timestamp 1644511149
transform 1 0 28520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__CLK
timestamp 1644511149
transform 1 0 33120 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__CLK
timestamp 1644511149
transform 1 0 35880 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__CLK
timestamp 1644511149
transform 1 0 28336 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__CLK
timestamp 1644511149
transform 1 0 28888 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__CLK
timestamp 1644511149
transform 1 0 34776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__CLK
timestamp 1644511149
transform 1 0 35236 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__CLK
timestamp 1644511149
transform 1 0 35604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__CLK
timestamp 1644511149
transform 1 0 35144 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__CLK
timestamp 1644511149
transform 1 0 35420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__CLK
timestamp 1644511149
transform 1 0 32016 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__CLK
timestamp 1644511149
transform -1 0 15180 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__CLK
timestamp 1644511149
transform 1 0 11592 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__CLK
timestamp 1644511149
transform 1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__CLK
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__CLK
timestamp 1644511149
transform 1 0 5336 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__CLK
timestamp 1644511149
transform -1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__CLK
timestamp 1644511149
transform -1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__CLK
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__CLK
timestamp 1644511149
transform -1 0 19596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__CLK
timestamp 1644511149
transform 1 0 29808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__CLK
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__CLK
timestamp 1644511149
transform 1 0 28796 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__CLK
timestamp 1644511149
transform -1 0 23000 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__CLK
timestamp 1644511149
transform 1 0 30544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__CLK
timestamp 1644511149
transform 1 0 20884 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__CLK
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__CLK
timestamp 1644511149
transform 1 0 29808 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__CLK
timestamp 1644511149
transform -1 0 32936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__CLK
timestamp 1644511149
transform 1 0 34684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__CLK
timestamp 1644511149
transform 1 0 36156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__CLK
timestamp 1644511149
transform 1 0 34040 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__CLK
timestamp 1644511149
transform 1 0 34040 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__CLK
timestamp 1644511149
transform 1 0 31280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__A
timestamp 1644511149
transform -1 0 25484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1644511149
transform -1 0 20240 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 2208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 1564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 2208 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 2208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 1564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 2208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 1564 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 2208 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 1564 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 2208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 2208 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 1564 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 2208 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 2208 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 2208 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 2208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 2208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 2208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1644511149
transform -1 0 1564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1644511149
transform -1 0 2208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1644511149
transform -1 0 2208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1644511149
transform -1 0 2208 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1644511149
transform -1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1644511149
transform -1 0 29992 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1644511149
transform -1 0 37444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1644511149
transform -1 0 37536 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output30_A
timestamp 1644511149
transform -1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output34_A
timestamp 1644511149
transform 1 0 37628 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output35_A
timestamp 1644511149
transform -1 0 37444 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1644511149
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1644511149
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_17
timestamp 1644511149
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1644511149
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_29
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1644511149
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_92
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_104
timestamp 1644511149
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_147
timestamp 1644511149
transform 1 0 14628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_153
timestamp 1644511149
transform 1 0 15180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1644511149
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_201
timestamp 1644511149
transform 1 0 19596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_213
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1644511149
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_233
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_238
timestamp 1644511149
transform 1 0 23000 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_258
timestamp 1644511149
transform 1 0 24840 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_270
timestamp 1644511149
transform 1 0 25944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_287 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_291
timestamp 1644511149
transform 1 0 27876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_303
timestamp 1644511149
transform 1 0 28980 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_315
timestamp 1644511149
transform 1 0 30084 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_327
timestamp 1644511149
transform 1 0 31188 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_343
timestamp 1644511149
transform 1 0 32660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_346
timestamp 1644511149
transform 1 0 32936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_366
timestamp 1644511149
transform 1 0 34776 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1644511149
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_6
timestamp 1644511149
transform 1 0 1656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_12
timestamp 1644511149
transform 1 0 2208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_16
timestamp 1644511149
transform 1 0 2576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_51
timestamp 1644511149
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_63
timestamp 1644511149
transform 1 0 6900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1644511149
transform 1 0 9660 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_110
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_116
timestamp 1644511149
transform 1 0 11776 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_128
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_182
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1644511149
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_218
timestamp 1644511149
transform 1 0 21160 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_230
timestamp 1644511149
transform 1 0 22264 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_236
timestamp 1644511149
transform 1 0 22816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_246
timestamp 1644511149
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_256
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_268
timestamp 1644511149
transform 1 0 25760 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_280
timestamp 1644511149
transform 1 0 26864 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_311
timestamp 1644511149
transform 1 0 29716 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_319
timestamp 1644511149
transform 1 0 30452 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp 1644511149
transform 1 0 30728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_343
timestamp 1644511149
transform 1 0 32660 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_355
timestamp 1644511149
transform 1 0 33764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_371
timestamp 1644511149
transform 1 0 35236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_383
timestamp 1644511149
transform 1 0 36340 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_395
timestamp 1644511149
transform 1 0 37444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_12
timestamp 1644511149
transform 1 0 2208 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_18
timestamp 1644511149
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_35
timestamp 1644511149
transform 1 0 4324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_42
timestamp 1644511149
transform 1 0 4968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1644511149
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_75
timestamp 1644511149
transform 1 0 8004 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_87
timestamp 1644511149
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_99
timestamp 1644511149
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1644511149
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_121
timestamp 1644511149
transform 1 0 12236 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_133
timestamp 1644511149
transform 1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_139
timestamp 1644511149
transform 1 0 13892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_145
timestamp 1644511149
transform 1 0 14444 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_148
timestamp 1644511149
transform 1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_175
timestamp 1644511149
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_179
timestamp 1644511149
transform 1 0 17572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_191
timestamp 1644511149
transform 1 0 18676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_199
timestamp 1644511149
transform 1 0 19412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_206
timestamp 1644511149
transform 1 0 20056 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1644511149
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_250
timestamp 1644511149
transform 1 0 24104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_259
timestamp 1644511149
transform 1 0 24932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_271
timestamp 1644511149
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_288
timestamp 1644511149
transform 1 0 27600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_308
timestamp 1644511149
transform 1 0 29440 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_314
timestamp 1644511149
transform 1 0 29992 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_326
timestamp 1644511149
transform 1 0 31096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1644511149
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_355
timestamp 1644511149
transform 1 0 33764 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_359
timestamp 1644511149
transform 1 0 34132 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_383
timestamp 1644511149
transform 1 0 36340 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 1644511149
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_43
timestamp 1644511149
transform 1 0 5060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_57
timestamp 1644511149
transform 1 0 6348 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_61
timestamp 1644511149
transform 1 0 6716 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_71
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_101
timestamp 1644511149
transform 1 0 10396 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1644511149
transform 1 0 11960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_124
timestamp 1644511149
transform 1 0 12512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_146
timestamp 1644511149
transform 1 0 14536 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_161
timestamp 1644511149
transform 1 0 15916 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_173
timestamp 1644511149
transform 1 0 17020 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_181
timestamp 1644511149
transform 1 0 17756 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_201
timestamp 1644511149
transform 1 0 19596 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_211
timestamp 1644511149
transform 1 0 20516 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_217
timestamp 1644511149
transform 1 0 21068 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_229
timestamp 1644511149
transform 1 0 22172 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_241
timestamp 1644511149
transform 1 0 23276 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_262
timestamp 1644511149
transform 1 0 25208 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_274
timestamp 1644511149
transform 1 0 26312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_278
timestamp 1644511149
transform 1 0 26680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_284
timestamp 1644511149
transform 1 0 27232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_297
timestamp 1644511149
transform 1 0 28428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_328
timestamp 1644511149
transform 1 0 31280 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_340
timestamp 1644511149
transform 1 0 32384 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_352
timestamp 1644511149
transform 1 0 33488 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_373
timestamp 1644511149
transform 1 0 35420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_385
timestamp 1644511149
transform 1 0 36524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_393
timestamp 1644511149
transform 1 0 37260 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1644511149
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1644511149
transform 1 0 1656 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_12
timestamp 1644511149
transform 1 0 2208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp 1644511149
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1644511149
transform 1 0 4048 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1644511149
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_67
timestamp 1644511149
transform 1 0 7268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_88
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_96
timestamp 1644511149
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1644511149
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_126
timestamp 1644511149
transform 1 0 12696 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_138
timestamp 1644511149
transform 1 0 13800 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_150
timestamp 1644511149
transform 1 0 14904 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1644511149
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1644511149
transform 1 0 18124 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_208
timestamp 1644511149
transform 1 0 20240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_214
timestamp 1644511149
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1644511149
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1644511149
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_299
timestamp 1644511149
transform 1 0 28612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_311
timestamp 1644511149
transform 1 0 29716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_314
timestamp 1644511149
transform 1 0 29992 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_322
timestamp 1644511149
transform 1 0 30728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_327
timestamp 1644511149
transform 1 0 31188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1644511149
transform 1 0 34868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_379
timestamp 1644511149
transform 1 0 35972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1644511149
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_31
timestamp 1644511149
transform 1 0 3956 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1644511149
transform 1 0 4968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_55
timestamp 1644511149
transform 1 0 6164 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_61
timestamp 1644511149
transform 1 0 6716 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_69
timestamp 1644511149
transform 1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_87
timestamp 1644511149
transform 1 0 9108 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_95
timestamp 1644511149
transform 1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_102
timestamp 1644511149
transform 1 0 10488 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_114
timestamp 1644511149
transform 1 0 11592 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_126
timestamp 1644511149
transform 1 0 12696 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1644511149
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1644511149
transform 1 0 14720 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_154
timestamp 1644511149
transform 1 0 15272 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_162
timestamp 1644511149
transform 1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_167
timestamp 1644511149
transform 1 0 16468 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_179
timestamp 1644511149
transform 1 0 17572 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1644511149
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_206
timestamp 1644511149
transform 1 0 20056 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_214
timestamp 1644511149
transform 1 0 20792 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_226
timestamp 1644511149
transform 1 0 21896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1644511149
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_288
timestamp 1644511149
transform 1 0 27600 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_300
timestamp 1644511149
transform 1 0 28704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_313
timestamp 1644511149
transform 1 0 29900 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_323
timestamp 1644511149
transform 1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_332
timestamp 1644511149
transform 1 0 31648 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_344
timestamp 1644511149
transform 1 0 32752 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_356
timestamp 1644511149
transform 1 0 33856 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_11
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_28
timestamp 1644511149
transform 1 0 3680 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_43
timestamp 1644511149
transform 1 0 5060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 1644511149
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_77
timestamp 1644511149
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_141
timestamp 1644511149
transform 1 0 14076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_151
timestamp 1644511149
transform 1 0 14996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_177
timestamp 1644511149
transform 1 0 17388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_189
timestamp 1644511149
transform 1 0 18492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_201
timestamp 1644511149
transform 1 0 19596 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1644511149
transform 1 0 20516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_228
timestamp 1644511149
transform 1 0 22080 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_240
timestamp 1644511149
transform 1 0 23184 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1644511149
transform 1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1644511149
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_341
timestamp 1644511149
transform 1 0 32476 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_353
timestamp 1644511149
transform 1 0 33580 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_359
timestamp 1644511149
transform 1 0 34132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1644511149
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp 1644511149
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_12
timestamp 1644511149
transform 1 0 2208 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1644511149
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_40
timestamp 1644511149
transform 1 0 4784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1644511149
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_52
timestamp 1644511149
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_64
timestamp 1644511149
transform 1 0 6992 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1644511149
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_94
timestamp 1644511149
transform 1 0 9752 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_106
timestamp 1644511149
transform 1 0 10856 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_118
timestamp 1644511149
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1644511149
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1644511149
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1644511149
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_199
timestamp 1644511149
transform 1 0 19412 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_230
timestamp 1644511149
transform 1 0 22264 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_242
timestamp 1644511149
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1644511149
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_273
timestamp 1644511149
transform 1 0 26220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_279
timestamp 1644511149
transform 1 0 26772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_291
timestamp 1644511149
transform 1 0 27876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_299
timestamp 1644511149
transform 1 0 28612 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1644511149
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_314
timestamp 1644511149
transform 1 0 29992 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_322
timestamp 1644511149
transform 1 0 30728 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_330
timestamp 1644511149
transform 1 0 31464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_350
timestamp 1644511149
transform 1 0 33304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1644511149
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_373
timestamp 1644511149
transform 1 0 35420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_379
timestamp 1644511149
transform 1 0 35972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_399
timestamp 1644511149
transform 1 0 37812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_102
timestamp 1644511149
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1644511149
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_121
timestamp 1644511149
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_144
timestamp 1644511149
transform 1 0 14352 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_159
timestamp 1644511149
transform 1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_177
timestamp 1644511149
transform 1 0 17388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_189
timestamp 1644511149
transform 1 0 18492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_201
timestamp 1644511149
transform 1 0 19596 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_207
timestamp 1644511149
transform 1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1644511149
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_235
timestamp 1644511149
transform 1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_243
timestamp 1644511149
transform 1 0 23460 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_265
timestamp 1644511149
transform 1 0 25484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1644511149
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_284
timestamp 1644511149
transform 1 0 27232 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_311
timestamp 1644511149
transform 1 0 29716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_322
timestamp 1644511149
transform 1 0 30728 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1644511149
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_341
timestamp 1644511149
transform 1 0 32476 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_354
timestamp 1644511149
transform 1 0 33672 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_366
timestamp 1644511149
transform 1 0 34776 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_378
timestamp 1644511149
transform 1 0 35880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_383
timestamp 1644511149
transform 1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_6
timestamp 1644511149
transform 1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_12
timestamp 1644511149
transform 1 0 2208 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_64
timestamp 1644511149
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1644511149
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_105
timestamp 1644511149
transform 1 0 10764 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_128
timestamp 1644511149
transform 1 0 12880 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_149
timestamp 1644511149
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_173
timestamp 1644511149
transform 1 0 17020 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_179
timestamp 1644511149
transform 1 0 17572 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_184
timestamp 1644511149
transform 1 0 18032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_190
timestamp 1644511149
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_219
timestamp 1644511149
transform 1 0 21252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1644511149
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1644511149
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_261
timestamp 1644511149
transform 1 0 25116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_284
timestamp 1644511149
transform 1 0 27232 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_296
timestamp 1644511149
transform 1 0 28336 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_319
timestamp 1644511149
transform 1 0 30452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_331
timestamp 1644511149
transform 1 0 31556 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_343
timestamp 1644511149
transform 1 0 32660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_355
timestamp 1644511149
transform 1 0 33764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_369
timestamp 1644511149
transform 1 0 35052 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_375
timestamp 1644511149
transform 1 0 35604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_387
timestamp 1644511149
transform 1 0 36708 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_399
timestamp 1644511149
transform 1 0 37812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_59
timestamp 1644511149
transform 1 0 6532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_72
timestamp 1644511149
transform 1 0 7728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_84
timestamp 1644511149
transform 1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1644511149
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_117
timestamp 1644511149
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1644511149
transform 1 0 13892 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_151
timestamp 1644511149
transform 1 0 14996 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp 1644511149
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_173
timestamp 1644511149
transform 1 0 17020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_185
timestamp 1644511149
transform 1 0 18124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_197
timestamp 1644511149
transform 1 0 19228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_209
timestamp 1644511149
transform 1 0 20332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1644511149
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_245
timestamp 1644511149
transform 1 0 23644 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_256
timestamp 1644511149
transform 1 0 24656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_260
timestamp 1644511149
transform 1 0 25024 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_265
timestamp 1644511149
transform 1 0 25484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1644511149
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_297
timestamp 1644511149
transform 1 0 28428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_303
timestamp 1644511149
transform 1 0 28980 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_311
timestamp 1644511149
transform 1 0 29716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_324
timestamp 1644511149
transform 1 0 30912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1644511149
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_359
timestamp 1644511149
transform 1 0 34132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_369
timestamp 1644511149
transform 1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_377
timestamp 1644511149
transform 1 0 35788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp 1644511149
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_5
timestamp 1644511149
transform 1 0 1564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1644511149
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_49
timestamp 1644511149
transform 1 0 5612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1644511149
transform 1 0 6808 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_74
timestamp 1644511149
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1644511149
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1644511149
transform 1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_110
timestamp 1644511149
transform 1 0 11224 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1644511149
transform 1 0 11776 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_120
timestamp 1644511149
transform 1 0 12144 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1644511149
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_176
timestamp 1644511149
transform 1 0 17296 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_188
timestamp 1644511149
transform 1 0 18400 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_201
timestamp 1644511149
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_205
timestamp 1644511149
transform 1 0 19964 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_211
timestamp 1644511149
transform 1 0 20516 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_218
timestamp 1644511149
transform 1 0 21160 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_230
timestamp 1644511149
transform 1 0 22264 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_242
timestamp 1644511149
transform 1 0 23368 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1644511149
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_261
timestamp 1644511149
transform 1 0 25116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_283
timestamp 1644511149
transform 1 0 27140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_295
timestamp 1644511149
transform 1 0 28244 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1644511149
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_319
timestamp 1644511149
transform 1 0 30452 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1644511149
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_374
timestamp 1644511149
transform 1 0 35512 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_381
timestamp 1644511149
transform 1 0 36156 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_393
timestamp 1644511149
transform 1 0 37260 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1644511149
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_6
timestamp 1644511149
transform 1 0 1656 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_14
timestamp 1644511149
transform 1 0 2392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1644511149
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_30
timestamp 1644511149
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_42
timestamp 1644511149
transform 1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_46
timestamp 1644511149
transform 1 0 5336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1644511149
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_59
timestamp 1644511149
transform 1 0 6532 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_92
timestamp 1644511149
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1644511149
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1644511149
transform 1 0 12420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1644511149
transform 1 0 13524 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_147
timestamp 1644511149
transform 1 0 14628 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_153
timestamp 1644511149
transform 1 0 15180 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_157
timestamp 1644511149
transform 1 0 15548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_245
timestamp 1644511149
transform 1 0 23644 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_258
timestamp 1644511149
transform 1 0 24840 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_270
timestamp 1644511149
transform 1 0 25944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1644511149
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_291
timestamp 1644511149
transform 1 0 27876 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_302
timestamp 1644511149
transform 1 0 28888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_310
timestamp 1644511149
transform 1 0 29624 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_330
timestamp 1644511149
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_343
timestamp 1644511149
transform 1 0 32660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_346
timestamp 1644511149
transform 1 0 32936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_354
timestamp 1644511149
transform 1 0 33672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_364
timestamp 1644511149
transform 1 0 34592 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_384
timestamp 1644511149
transform 1 0 36432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1644511149
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1644511149
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1644511149
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 1644511149
transform 1 0 6716 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_67
timestamp 1644511149
transform 1 0 7268 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1644511149
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_119
timestamp 1644511149
transform 1 0 12052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_126
timestamp 1644511149
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1644511149
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1644511149
transform 1 0 14812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_157
timestamp 1644511149
transform 1 0 15548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1644511149
transform 1 0 16100 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_171
timestamp 1644511149
transform 1 0 16836 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_174
timestamp 1644511149
transform 1 0 17112 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_186
timestamp 1644511149
transform 1 0 18216 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1644511149
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_205
timestamp 1644511149
transform 1 0 19964 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1644511149
transform 1 0 20884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_225
timestamp 1644511149
transform 1 0 21804 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_237
timestamp 1644511149
transform 1 0 22908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1644511149
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_274
timestamp 1644511149
transform 1 0 26312 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_286
timestamp 1644511149
transform 1 0 27416 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_298
timestamp 1644511149
transform 1 0 28520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1644511149
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1644511149
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_318
timestamp 1644511149
transform 1 0 30360 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_325
timestamp 1644511149
transform 1 0 31004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_334
timestamp 1644511149
transform 1 0 31832 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_346
timestamp 1644511149
transform 1 0 32936 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1644511149
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_384
timestamp 1644511149
transform 1 0 36432 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_396
timestamp 1644511149
transform 1 0 37536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_403
timestamp 1644511149
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_12
timestamp 1644511149
transform 1 0 2208 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_18
timestamp 1644511149
transform 1 0 2760 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_28
timestamp 1644511149
transform 1 0 3680 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_99
timestamp 1644511149
transform 1 0 10212 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1644511149
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1644511149
transform 1 0 13524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_139
timestamp 1644511149
transform 1 0 13892 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_143
timestamp 1644511149
transform 1 0 14260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_156
timestamp 1644511149
transform 1 0 15456 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1644511149
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 1644511149
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_191
timestamp 1644511149
transform 1 0 18676 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp 1644511149
transform 1 0 19412 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_203
timestamp 1644511149
transform 1 0 19780 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_210
timestamp 1644511149
transform 1 0 20424 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1644511149
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_229
timestamp 1644511149
transform 1 0 22172 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_241
timestamp 1644511149
transform 1 0 23276 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_253
timestamp 1644511149
transform 1 0 24380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_265
timestamp 1644511149
transform 1 0 25484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1644511149
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_309
timestamp 1644511149
transform 1 0 29532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_312
timestamp 1644511149
transform 1 0 29808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_320
timestamp 1644511149
transform 1 0 30544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_328
timestamp 1644511149
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_369
timestamp 1644511149
transform 1 0 35052 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_381
timestamp 1644511149
transform 1 0 36156 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1644511149
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1644511149
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_111
timestamp 1644511149
transform 1 0 11316 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_127
timestamp 1644511149
transform 1 0 12788 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_132
timestamp 1644511149
transform 1 0 13248 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1644511149
transform 1 0 14444 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_161
timestamp 1644511149
transform 1 0 15916 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_169
timestamp 1644511149
transform 1 0 16652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_172
timestamp 1644511149
transform 1 0 16928 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1644511149
transform 1 0 17480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_200
timestamp 1644511149
transform 1 0 19504 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_208
timestamp 1644511149
transform 1 0 20240 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1644511149
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_225
timestamp 1644511149
transform 1 0 21804 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_235
timestamp 1644511149
transform 1 0 22724 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_243
timestamp 1644511149
transform 1 0 23460 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1644511149
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_280
timestamp 1644511149
transform 1 0 26864 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_300
timestamp 1644511149
transform 1 0 28704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_311
timestamp 1644511149
transform 1 0 29716 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_319
timestamp 1644511149
transform 1 0 30452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_324
timestamp 1644511149
transform 1 0 30912 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_336
timestamp 1644511149
transform 1 0 32016 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_342
timestamp 1644511149
transform 1 0 32568 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_347
timestamp 1644511149
transform 1 0 33028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_359
timestamp 1644511149
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_5
timestamp 1644511149
transform 1 0 1564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_17
timestamp 1644511149
transform 1 0 2668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_29
timestamp 1644511149
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_41
timestamp 1644511149
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1644511149
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_60
timestamp 1644511149
transform 1 0 6624 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_72
timestamp 1644511149
transform 1 0 7728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_84
timestamp 1644511149
transform 1 0 8832 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_96
timestamp 1644511149
transform 1 0 9936 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1644511149
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1644511149
transform 1 0 11868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1644511149
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1644511149
transform 1 0 13892 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_151
timestamp 1644511149
transform 1 0 14996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_159
timestamp 1644511149
transform 1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1644511149
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_182
timestamp 1644511149
transform 1 0 17848 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_200
timestamp 1644511149
transform 1 0 19504 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_210
timestamp 1644511149
transform 1 0 20424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_231
timestamp 1644511149
transform 1 0 22356 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_243
timestamp 1644511149
transform 1 0 23460 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_255
timestamp 1644511149
transform 1 0 24564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_263
timestamp 1644511149
transform 1 0 25300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1644511149
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_284
timestamp 1644511149
transform 1 0 27232 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_296
timestamp 1644511149
transform 1 0 28336 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_308
timestamp 1644511149
transform 1 0 29440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_315
timestamp 1644511149
transform 1 0 30084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_321
timestamp 1644511149
transform 1 0 30636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1644511149
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_6
timestamp 1644511149
transform 1 0 1656 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_14
timestamp 1644511149
transform 1 0 2392 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1644511149
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1644511149
transform 1 0 7176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1644511149
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1644511149
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1644511149
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_115
timestamp 1644511149
transform 1 0 11684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_125
timestamp 1644511149
transform 1 0 12604 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1644511149
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_143
timestamp 1644511149
transform 1 0 14260 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_155
timestamp 1644511149
transform 1 0 15364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_167
timestamp 1644511149
transform 1 0 16468 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_179
timestamp 1644511149
transform 1 0 17572 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1644511149
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1644511149
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_208
timestamp 1644511149
transform 1 0 20240 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_220
timestamp 1644511149
transform 1 0 21344 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_232
timestamp 1644511149
transform 1 0 22448 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1644511149
transform 1 0 23092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_272
timestamp 1644511149
transform 1 0 26128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_278
timestamp 1644511149
transform 1 0 26680 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_290
timestamp 1644511149
transform 1 0 27784 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_302
timestamp 1644511149
transform 1 0 28888 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_375
timestamp 1644511149
transform 1 0 35604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_395
timestamp 1644511149
transform 1 0 37444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_21
timestamp 1644511149
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_33
timestamp 1644511149
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_37
timestamp 1644511149
transform 1 0 4508 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_41
timestamp 1644511149
transform 1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1644511149
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1644511149
transform 1 0 8188 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_100
timestamp 1644511149
transform 1 0 10304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1644511149
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_121
timestamp 1644511149
transform 1 0 12236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_135
timestamp 1644511149
transform 1 0 13524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 1644511149
transform 1 0 14996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_155
timestamp 1644511149
transform 1 0 15364 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_158
timestamp 1644511149
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1644511149
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_176
timestamp 1644511149
transform 1 0 17296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_190
timestamp 1644511149
transform 1 0 18584 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1644511149
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_207
timestamp 1644511149
transform 1 0 20148 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1644511149
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_229
timestamp 1644511149
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_251
timestamp 1644511149
transform 1 0 24196 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_263
timestamp 1644511149
transform 1 0 25300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1644511149
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_284
timestamp 1644511149
transform 1 0 27232 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_296
timestamp 1644511149
transform 1 0 28336 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_308
timestamp 1644511149
transform 1 0 29440 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_315
timestamp 1644511149
transform 1 0 30084 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_327
timestamp 1644511149
transform 1 0 31188 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_366
timestamp 1644511149
transform 1 0 34776 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_372
timestamp 1644511149
transform 1 0 35328 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1644511149
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_6
timestamp 1644511149
transform 1 0 1656 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_12
timestamp 1644511149
transform 1 0 2208 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1644511149
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_89
timestamp 1644511149
transform 1 0 9292 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_100
timestamp 1644511149
transform 1 0 10304 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 1644511149
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_116
timestamp 1644511149
transform 1 0 11776 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_122
timestamp 1644511149
transform 1 0 12328 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_125
timestamp 1644511149
transform 1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_129
timestamp 1644511149
transform 1 0 12972 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_149
timestamp 1644511149
transform 1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_156
timestamp 1644511149
transform 1 0 15456 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1644511149
transform 1 0 16376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_176
timestamp 1644511149
transform 1 0 17296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_182
timestamp 1644511149
transform 1 0 17848 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1644511149
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1644511149
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_208
timestamp 1644511149
transform 1 0 20240 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_220
timestamp 1644511149
transform 1 0 21344 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_228
timestamp 1644511149
transform 1 0 22080 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_234
timestamp 1644511149
transform 1 0 22632 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 1644511149
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_272
timestamp 1644511149
transform 1 0 26128 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_292
timestamp 1644511149
transform 1 0 27968 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_298
timestamp 1644511149
transform 1 0 28520 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1644511149
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_325
timestamp 1644511149
transform 1 0 31004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_338
timestamp 1644511149
transform 1 0 32200 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_346
timestamp 1644511149
transform 1 0 32936 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_352
timestamp 1644511149
transform 1 0 33488 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_385
timestamp 1644511149
transform 1 0 36524 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_397
timestamp 1644511149
transform 1 0 37628 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1644511149
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_23
timestamp 1644511149
transform 1 0 3220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1644511149
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_68
timestamp 1644511149
transform 1 0 7360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_80
timestamp 1644511149
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_103
timestamp 1644511149
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1644511149
transform 1 0 12420 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_150
timestamp 1644511149
transform 1 0 14904 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1644511149
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_172
timestamp 1644511149
transform 1 0 16928 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_179
timestamp 1644511149
transform 1 0 17572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1644511149
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_195
timestamp 1644511149
transform 1 0 19044 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_198
timestamp 1644511149
transform 1 0 19320 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_210
timestamp 1644511149
transform 1 0 20424 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1644511149
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1644511149
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_299
timestamp 1644511149
transform 1 0 28612 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_308
timestamp 1644511149
transform 1 0 29440 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_318
timestamp 1644511149
transform 1 0 30360 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_328
timestamp 1644511149
transform 1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_354
timestamp 1644511149
transform 1 0 33672 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_358
timestamp 1644511149
transform 1 0 34040 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_364
timestamp 1644511149
transform 1 0 34592 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_374
timestamp 1644511149
transform 1 0 35512 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_386
timestamp 1644511149
transform 1 0 36616 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_396
timestamp 1644511149
transform 1 0 37536 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_404
timestamp 1644511149
transform 1 0 38272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1644511149
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1644511149
transform 1 0 4048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_36
timestamp 1644511149
transform 1 0 4416 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_47
timestamp 1644511149
transform 1 0 5428 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_74
timestamp 1644511149
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1644511149
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_94
timestamp 1644511149
transform 1 0 9752 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_104
timestamp 1644511149
transform 1 0 10672 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_116
timestamp 1644511149
transform 1 0 11776 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_128
timestamp 1644511149
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_160
timestamp 1644511149
transform 1 0 15824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_185
timestamp 1644511149
transform 1 0 18124 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_204
timestamp 1644511149
transform 1 0 19872 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1644511149
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_244
timestamp 1644511149
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_273
timestamp 1644511149
transform 1 0 26220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_286
timestamp 1644511149
transform 1 0 27416 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_298
timestamp 1644511149
transform 1 0 28520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1644511149
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_320
timestamp 1644511149
transform 1 0 30544 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_332
timestamp 1644511149
transform 1 0 31648 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_344
timestamp 1644511149
transform 1 0 32752 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_351
timestamp 1644511149
transform 1 0 33396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1644511149
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_369
timestamp 1644511149
transform 1 0 35052 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_381
timestamp 1644511149
transform 1 0 36156 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_395
timestamp 1644511149
transform 1 0 37444 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1644511149
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_6
timestamp 1644511149
transform 1 0 1656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_12
timestamp 1644511149
transform 1 0 2208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_24
timestamp 1644511149
transform 1 0 3312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_30
timestamp 1644511149
transform 1 0 3864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_65
timestamp 1644511149
transform 1 0 7084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_89
timestamp 1644511149
transform 1 0 9292 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_99
timestamp 1644511149
transform 1 0 10212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_121
timestamp 1644511149
transform 1 0 12236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_145
timestamp 1644511149
transform 1 0 14444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_157
timestamp 1644511149
transform 1 0 15548 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_191
timestamp 1644511149
transform 1 0 18676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_203
timestamp 1644511149
transform 1 0 19780 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_212
timestamp 1644511149
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_233
timestamp 1644511149
transform 1 0 22540 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1644511149
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_302
timestamp 1644511149
transform 1 0 28888 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_310
timestamp 1644511149
transform 1 0 29624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_313
timestamp 1644511149
transform 1 0 29900 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_325
timestamp 1644511149
transform 1 0 31004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1644511149
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_369
timestamp 1644511149
transform 1 0 35052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_375
timestamp 1644511149
transform 1 0 35604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_387
timestamp 1644511149
transform 1 0 36708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_51
timestamp 1644511149
transform 1 0 5796 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_58
timestamp 1644511149
transform 1 0 6440 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_66
timestamp 1644511149
transform 1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_72
timestamp 1644511149
transform 1 0 7728 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_88
timestamp 1644511149
transform 1 0 9200 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_100
timestamp 1644511149
transform 1 0 10304 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_112
timestamp 1644511149
transform 1 0 11408 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_118
timestamp 1644511149
transform 1 0 11960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 1644511149
transform 1 0 12880 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1644511149
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_157
timestamp 1644511149
transform 1 0 15548 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_170
timestamp 1644511149
transform 1 0 16744 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1644511149
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_184
timestamp 1644511149
transform 1 0 18032 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_207
timestamp 1644511149
transform 1 0 20148 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1644511149
transform 1 0 20700 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_235
timestamp 1644511149
transform 1 0 22724 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_239
timestamp 1644511149
transform 1 0 23092 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1644511149
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_271
timestamp 1644511149
transform 1 0 26036 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_283
timestamp 1644511149
transform 1 0 27140 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_292
timestamp 1644511149
transform 1 0 27968 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_298
timestamp 1644511149
transform 1 0 28520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1644511149
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_317
timestamp 1644511149
transform 1 0 30268 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_329
timestamp 1644511149
transform 1 0 31372 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_337
timestamp 1644511149
transform 1 0 32108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_344
timestamp 1644511149
transform 1 0 32752 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1644511149
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_373
timestamp 1644511149
transform 1 0 35420 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_381
timestamp 1644511149
transform 1 0 36156 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_393
timestamp 1644511149
transform 1 0 37260 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1644511149
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_12
timestamp 1644511149
transform 1 0 2208 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_20
timestamp 1644511149
transform 1 0 2944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_60
timestamp 1644511149
transform 1 0 6624 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_72
timestamp 1644511149
transform 1 0 7728 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_84
timestamp 1644511149
transform 1 0 8832 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_129
timestamp 1644511149
transform 1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1644511149
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1644511149
transform 1 0 14628 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_159
timestamp 1644511149
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1644511149
transform 1 0 17296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1644511149
transform 1 0 18032 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1644511149
transform 1 0 19136 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_208
timestamp 1644511149
transform 1 0 20240 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_254
timestamp 1644511149
transform 1 0 24472 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_288
timestamp 1644511149
transform 1 0 27600 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_301
timestamp 1644511149
transform 1 0 28796 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_313
timestamp 1644511149
transform 1 0 29900 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_325
timestamp 1644511149
transform 1 0 31004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1644511149
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_371
timestamp 1644511149
transform 1 0 35236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_383
timestamp 1644511149
transform 1 0 36340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1644511149
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_38
timestamp 1644511149
transform 1 0 4600 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_50
timestamp 1644511149
transform 1 0 5704 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_62
timestamp 1644511149
transform 1 0 6808 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_73
timestamp 1644511149
transform 1 0 7820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1644511149
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_108
timestamp 1644511149
transform 1 0 11040 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_120
timestamp 1644511149
transform 1 0 12144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_124
timestamp 1644511149
transform 1 0 12512 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_131
timestamp 1644511149
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_168
timestamp 1644511149
transform 1 0 16560 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_176
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_184
timestamp 1644511149
transform 1 0 18032 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1644511149
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_214
timestamp 1644511149
transform 1 0 20792 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_226
timestamp 1644511149
transform 1 0 21896 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_238
timestamp 1644511149
transform 1 0 23000 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_294
timestamp 1644511149
transform 1 0 28152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_300
timestamp 1644511149
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_311
timestamp 1644511149
transform 1 0 29716 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_320
timestamp 1644511149
transform 1 0 30544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_332
timestamp 1644511149
transform 1 0 31648 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_344
timestamp 1644511149
transform 1 0 32752 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_356
timestamp 1644511149
transform 1 0 33856 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_373
timestamp 1644511149
transform 1 0 35420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_393
timestamp 1644511149
transform 1 0 37260 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1644511149
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_5
timestamp 1644511149
transform 1 0 1564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_16
timestamp 1644511149
transform 1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_38
timestamp 1644511149
transform 1 0 4600 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_46
timestamp 1644511149
transform 1 0 5336 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1644511149
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_90
timestamp 1644511149
transform 1 0 9384 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_102
timestamp 1644511149
transform 1 0 10488 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1644511149
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1644511149
transform 1 0 12972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_154
timestamp 1644511149
transform 1 0 15272 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1644511149
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_194
timestamp 1644511149
transform 1 0 18952 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_206
timestamp 1644511149
transform 1 0 20056 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1644511149
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_231
timestamp 1644511149
transform 1 0 22356 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_238
timestamp 1644511149
transform 1 0 23000 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_248
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_260
timestamp 1644511149
transform 1 0 25024 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_272
timestamp 1644511149
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_285
timestamp 1644511149
transform 1 0 27324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_297
timestamp 1644511149
transform 1 0 28428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_310
timestamp 1644511149
transform 1 0 29624 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_323
timestamp 1644511149
transform 1 0 30820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_330
timestamp 1644511149
transform 1 0 31464 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_377
timestamp 1644511149
transform 1 0 35788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1644511149
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_6
timestamp 1644511149
transform 1 0 1656 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_14
timestamp 1644511149
transform 1 0 2392 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1644511149
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_38
timestamp 1644511149
transform 1 0 4600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_42
timestamp 1644511149
transform 1 0 4968 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_64
timestamp 1644511149
transform 1 0 6992 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_74
timestamp 1644511149
transform 1 0 7912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_95
timestamp 1644511149
transform 1 0 9844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_102
timestamp 1644511149
transform 1 0 10488 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_114
timestamp 1644511149
transform 1 0 11592 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_120
timestamp 1644511149
transform 1 0 12144 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_127
timestamp 1644511149
transform 1 0 12788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_134
timestamp 1644511149
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1644511149
transform 1 0 14352 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_156
timestamp 1644511149
transform 1 0 15456 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1644511149
transform 1 0 16376 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_180
timestamp 1644511149
transform 1 0 17664 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1644511149
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_199
timestamp 1644511149
transform 1 0 19412 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_205
timestamp 1644511149
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1644511149
transform 1 0 21988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1644511149
transform 1 0 23092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_311
timestamp 1644511149
transform 1 0 29716 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_319
timestamp 1644511149
transform 1 0 30452 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_323
timestamp 1644511149
transform 1 0 30820 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_344
timestamp 1644511149
transform 1 0 32752 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_350
timestamp 1644511149
transform 1 0 33304 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1644511149
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_373
timestamp 1644511149
transform 1 0 35420 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_385
timestamp 1644511149
transform 1 0 36524 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_395
timestamp 1644511149
transform 1 0 37444 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1644511149
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_21
timestamp 1644511149
transform 1 0 3036 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_25
timestamp 1644511149
transform 1 0 3404 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_34
timestamp 1644511149
transform 1 0 4232 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_42
timestamp 1644511149
transform 1 0 4968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1644511149
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_63
timestamp 1644511149
transform 1 0 6900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_73
timestamp 1644511149
transform 1 0 7820 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_79
timestamp 1644511149
transform 1 0 8372 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1644511149
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_150
timestamp 1644511149
transform 1 0 14904 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1644511149
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_177
timestamp 1644511149
transform 1 0 17388 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_200
timestamp 1644511149
transform 1 0 19504 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_209
timestamp 1644511149
transform 1 0 20332 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_233
timestamp 1644511149
transform 1 0 22540 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1644511149
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_265
timestamp 1644511149
transform 1 0 25484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1644511149
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_302
timestamp 1644511149
transform 1 0 28888 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_308
timestamp 1644511149
transform 1 0 29440 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_318
timestamp 1644511149
transform 1 0 30360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_327
timestamp 1644511149
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_345
timestamp 1644511149
transform 1 0 32844 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_357
timestamp 1644511149
transform 1 0 33948 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_369
timestamp 1644511149
transform 1 0 35052 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_374
timestamp 1644511149
transform 1 0 35512 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_386
timestamp 1644511149
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_397
timestamp 1644511149
transform 1 0 37628 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_6
timestamp 1644511149
transform 1 0 1656 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_12
timestamp 1644511149
transform 1 0 2208 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1644511149
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_44
timestamp 1644511149
transform 1 0 5152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1644511149
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_58
timestamp 1644511149
transform 1 0 6440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1644511149
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_67
timestamp 1644511149
transform 1 0 7268 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1644511149
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_87
timestamp 1644511149
transform 1 0 9108 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1644511149
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_95
timestamp 1644511149
transform 1 0 9844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_107
timestamp 1644511149
transform 1 0 10948 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_115
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_131
timestamp 1644511149
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1644511149
transform 1 0 14352 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1644511149
transform 1 0 15456 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_168
timestamp 1644511149
transform 1 0 16560 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_176
timestamp 1644511149
transform 1 0 17296 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_182
timestamp 1644511149
transform 1 0 17848 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_186
timestamp 1644511149
transform 1 0 18216 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1644511149
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_214
timestamp 1644511149
transform 1 0 20792 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_222
timestamp 1644511149
transform 1 0 21528 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1644511149
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_240
timestamp 1644511149
transform 1 0 23184 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1644511149
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_259
timestamp 1644511149
transform 1 0 24932 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_267
timestamp 1644511149
transform 1 0 25668 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1644511149
transform 1 0 26036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_278
timestamp 1644511149
transform 1 0 26680 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_282
timestamp 1644511149
transform 1 0 27048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_311
timestamp 1644511149
transform 1 0 29716 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_319
timestamp 1644511149
transform 1 0 30452 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_338
timestamp 1644511149
transform 1 0 32200 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_349
timestamp 1644511149
transform 1 0 33212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_353
timestamp 1644511149
transform 1 0 33580 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1644511149
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_369
timestamp 1644511149
transform 1 0 35052 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_11
timestamp 1644511149
transform 1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_35
timestamp 1644511149
transform 1 0 4324 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_43
timestamp 1644511149
transform 1 0 5060 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1644511149
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_61
timestamp 1644511149
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_65
timestamp 1644511149
transform 1 0 7084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_71
timestamp 1644511149
transform 1 0 7636 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_119
timestamp 1644511149
transform 1 0 12052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1644511149
transform 1 0 12420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_130
timestamp 1644511149
transform 1 0 13064 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_148
timestamp 1644511149
transform 1 0 14720 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1644511149
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_184
timestamp 1644511149
transform 1 0 18032 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_187
timestamp 1644511149
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_195
timestamp 1644511149
transform 1 0 19044 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_201
timestamp 1644511149
transform 1 0 19596 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_206
timestamp 1644511149
transform 1 0 20056 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_228
timestamp 1644511149
transform 1 0 22080 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_235
timestamp 1644511149
transform 1 0 22724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_239
timestamp 1644511149
transform 1 0 23092 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_242
timestamp 1644511149
transform 1 0 23368 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_256
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_268
timestamp 1644511149
transform 1 0 25760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_342
timestamp 1644511149
transform 1 0 32568 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_348
timestamp 1644511149
transform 1 0 33120 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_360
timestamp 1644511149
transform 1 0 34224 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_368
timestamp 1644511149
transform 1 0 34960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_388
timestamp 1644511149
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_17
timestamp 1644511149
transform 1 0 2668 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1644511149
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_47
timestamp 1644511149
transform 1 0 5428 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_59
timestamp 1644511149
transform 1 0 6532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_71
timestamp 1644511149
transform 1 0 7636 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_117
timestamp 1644511149
transform 1 0 11868 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_120
timestamp 1644511149
transform 1 0 12144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_134
timestamp 1644511149
transform 1 0 13432 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_166
timestamp 1644511149
transform 1 0 16376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1644511149
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_231
timestamp 1644511149
transform 1 0 22356 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_238
timestamp 1644511149
transform 1 0 23000 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_259
timestamp 1644511149
transform 1 0 24932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_281
timestamp 1644511149
transform 1 0 26956 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_293
timestamp 1644511149
transform 1 0 28060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1644511149
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_387
timestamp 1644511149
transform 1 0 36708 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_400
timestamp 1644511149
transform 1 0 37904 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1644511149
transform 1 0 38456 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_6
timestamp 1644511149
transform 1 0 1656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_12
timestamp 1644511149
transform 1 0 2208 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_20
timestamp 1644511149
transform 1 0 2944 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_25
timestamp 1644511149
transform 1 0 3404 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_37
timestamp 1644511149
transform 1 0 4508 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_41
timestamp 1644511149
transform 1 0 4876 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1644511149
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_90
timestamp 1644511149
transform 1 0 9384 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1644511149
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1644511149
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_117
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_129
timestamp 1644511149
transform 1 0 12972 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1644511149
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_141
timestamp 1644511149
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_153
timestamp 1644511149
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1644511149
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_190
timestamp 1644511149
transform 1 0 18584 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_198
timestamp 1644511149
transform 1 0 19320 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_202
timestamp 1644511149
transform 1 0 19688 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1644511149
transform 1 0 20240 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_247
timestamp 1644511149
transform 1 0 23828 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1644511149
transform 1 0 24748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1644511149
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_39
timestamp 1644511149
transform 1 0 4692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_64
timestamp 1644511149
transform 1 0 6992 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_76
timestamp 1644511149
transform 1 0 8096 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_99
timestamp 1644511149
transform 1 0 10212 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_113
timestamp 1644511149
transform 1 0 11500 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_123
timestamp 1644511149
transform 1 0 12420 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_127
timestamp 1644511149
transform 1 0 12788 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 1644511149
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_161
timestamp 1644511149
transform 1 0 15916 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_166
timestamp 1644511149
transform 1 0 16376 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_174
timestamp 1644511149
transform 1 0 17112 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_186
timestamp 1644511149
transform 1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1644511149
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_201
timestamp 1644511149
transform 1 0 19596 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_205
timestamp 1644511149
transform 1 0 19964 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_217
timestamp 1644511149
transform 1 0 21068 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_229
timestamp 1644511149
transform 1 0 22172 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1644511149
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_259
timestamp 1644511149
transform 1 0 24932 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_266
timestamp 1644511149
transform 1 0 25576 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_272
timestamp 1644511149
transform 1 0 26128 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_280
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 1644511149
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_315
timestamp 1644511149
transform 1 0 30084 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_328
timestamp 1644511149
transform 1 0 31280 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_340
timestamp 1644511149
transform 1 0 32384 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_352
timestamp 1644511149
transform 1 0 33488 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_6
timestamp 1644511149
transform 1 0 1656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_12
timestamp 1644511149
transform 1 0 2208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_16
timestamp 1644511149
transform 1 0 2576 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_38
timestamp 1644511149
transform 1 0 4600 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_44
timestamp 1644511149
transform 1 0 5152 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1644511149
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_63
timestamp 1644511149
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_70
timestamp 1644511149
transform 1 0 7544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_77
timestamp 1644511149
transform 1 0 8188 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_83
timestamp 1644511149
transform 1 0 8740 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_86
timestamp 1644511149
transform 1 0 9016 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_100
timestamp 1644511149
transform 1 0 10304 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp 1644511149
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_134
timestamp 1644511149
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_142
timestamp 1644511149
transform 1 0 14168 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_148
timestamp 1644511149
transform 1 0 14720 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1644511149
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1644511149
transform 1 0 18032 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_196
timestamp 1644511149
transform 1 0 19136 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_263
timestamp 1644511149
transform 1 0 25300 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1644511149
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1644511149
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_339
timestamp 1644511149
transform 1 0 32292 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_351
timestamp 1644511149
transform 1 0 33396 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_363
timestamp 1644511149
transform 1 0 34500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_375
timestamp 1644511149
transform 1 0 35604 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_380
timestamp 1644511149
transform 1 0 36064 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_403
timestamp 1644511149
transform 1 0 38180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1644511149
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_37
timestamp 1644511149
transform 1 0 4508 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_45
timestamp 1644511149
transform 1 0 5244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_59
timestamp 1644511149
transform 1 0 6532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_67
timestamp 1644511149
transform 1 0 7268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_75
timestamp 1644511149
transform 1 0 8004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_87
timestamp 1644511149
transform 1 0 9108 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_94
timestamp 1644511149
transform 1 0 9752 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_105
timestamp 1644511149
transform 1 0 10764 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_130
timestamp 1644511149
transform 1 0 13064 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_149
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_171
timestamp 1644511149
transform 1 0 16836 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1644511149
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_188
timestamp 1644511149
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_203
timestamp 1644511149
transform 1 0 19780 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_228
timestamp 1644511149
transform 1 0 22080 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_234
timestamp 1644511149
transform 1 0 22632 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_269
timestamp 1644511149
transform 1 0 25852 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_291
timestamp 1644511149
transform 1 0 27876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_299
timestamp 1644511149
transform 1 0 28612 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_318
timestamp 1644511149
transform 1 0 30360 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_342
timestamp 1644511149
transform 1 0 32568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_348
timestamp 1644511149
transform 1 0 33120 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_354
timestamp 1644511149
transform 1 0 33672 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_374
timestamp 1644511149
transform 1 0 35512 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_397
timestamp 1644511149
transform 1 0 37628 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1644511149
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_5
timestamp 1644511149
transform 1 0 1564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_17
timestamp 1644511149
transform 1 0 2668 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_46
timestamp 1644511149
transform 1 0 5336 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1644511149
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_60
timestamp 1644511149
transform 1 0 6624 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_66
timestamp 1644511149
transform 1 0 7176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_72
timestamp 1644511149
transform 1 0 7728 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_84
timestamp 1644511149
transform 1 0 8832 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_92
timestamp 1644511149
transform 1 0 9568 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_116
timestamp 1644511149
transform 1 0 11776 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_123
timestamp 1644511149
transform 1 0 12420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_131
timestamp 1644511149
transform 1 0 13156 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_143
timestamp 1644511149
transform 1 0 14260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_154
timestamp 1644511149
transform 1 0 15272 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1644511149
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_172
timestamp 1644511149
transform 1 0 16928 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_186
timestamp 1644511149
transform 1 0 18216 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_196
timestamp 1644511149
transform 1 0 19136 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_203
timestamp 1644511149
transform 1 0 19780 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_211
timestamp 1644511149
transform 1 0 20516 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_215
timestamp 1644511149
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_229
timestamp 1644511149
transform 1 0 22172 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_232
timestamp 1644511149
transform 1 0 22448 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_242
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_254
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_260
timestamp 1644511149
transform 1 0 25024 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_272
timestamp 1644511149
transform 1 0 26128 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_289
timestamp 1644511149
transform 1 0 27692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_301
timestamp 1644511149
transform 1 0 28796 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_314
timestamp 1644511149
transform 1 0 29992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_327
timestamp 1644511149
transform 1 0 31188 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_345
timestamp 1644511149
transform 1 0 32844 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_348
timestamp 1644511149
transform 1 0 33120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_357
timestamp 1644511149
transform 1 0 33948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_363
timestamp 1644511149
transform 1 0 34500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_384
timestamp 1644511149
transform 1 0 36432 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_6
timestamp 1644511149
transform 1 0 1656 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_17
timestamp 1644511149
transform 1 0 2668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1644511149
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_37
timestamp 1644511149
transform 1 0 4508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_49
timestamp 1644511149
transform 1 0 5612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_57
timestamp 1644511149
transform 1 0 6348 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_62
timestamp 1644511149
transform 1 0 6808 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_74
timestamp 1644511149
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1644511149
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_107
timestamp 1644511149
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_114
timestamp 1644511149
transform 1 0 11592 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_122
timestamp 1644511149
transform 1 0 12328 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_127
timestamp 1644511149
transform 1 0 12788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1644511149
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1644511149
transform 1 0 14812 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_172
timestamp 1644511149
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_182
timestamp 1644511149
transform 1 0 17848 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_205
timestamp 1644511149
transform 1 0 19964 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_212
timestamp 1644511149
transform 1 0 20608 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_224
timestamp 1644511149
transform 1 0 21712 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_236
timestamp 1644511149
transform 1 0 22816 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1644511149
transform 1 0 23092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_261
timestamp 1644511149
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1644511149
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_316
timestamp 1644511149
transform 1 0 30176 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_320
timestamp 1644511149
transform 1 0 30544 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_326
timestamp 1644511149
transform 1 0 31096 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1644511149
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_383
timestamp 1644511149
transform 1 0 36340 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_395
timestamp 1644511149
transform 1 0 37444 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_41
timestamp 1644511149
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1644511149
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_65
timestamp 1644511149
transform 1 0 7084 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_70
timestamp 1644511149
transform 1 0 7544 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_82
timestamp 1644511149
transform 1 0 8648 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_94
timestamp 1644511149
transform 1 0 9752 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_106
timestamp 1644511149
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1644511149
transform 1 0 12420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1644511149
transform 1 0 13524 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_147
timestamp 1644511149
transform 1 0 14628 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_151
timestamp 1644511149
transform 1 0 14996 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_155
timestamp 1644511149
transform 1 0 15364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_175
timestamp 1644511149
transform 1 0 17204 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_185
timestamp 1644511149
transform 1 0 18124 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_196
timestamp 1644511149
transform 1 0 19136 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_210
timestamp 1644511149
transform 1 0 20424 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1644511149
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_235
timestamp 1644511149
transform 1 0 22724 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_245
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_251
timestamp 1644511149
transform 1 0 24196 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_265
timestamp 1644511149
transform 1 0 25484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_271
timestamp 1644511149
transform 1 0 26036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_284
timestamp 1644511149
transform 1 0 27232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_290
timestamp 1644511149
transform 1 0 27784 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_315
timestamp 1644511149
transform 1 0 30084 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_321
timestamp 1644511149
transform 1 0 30636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 1644511149
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_345
timestamp 1644511149
transform 1 0 32844 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_357
timestamp 1644511149
transform 1 0 33948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_364
timestamp 1644511149
transform 1 0 34592 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_370
timestamp 1644511149
transform 1 0 35144 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_382
timestamp 1644511149
transform 1 0 36248 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1644511149
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_6
timestamp 1644511149
transform 1 0 1656 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_12
timestamp 1644511149
transform 1 0 2208 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1644511149
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_36
timestamp 1644511149
transform 1 0 4416 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_43
timestamp 1644511149
transform 1 0 5060 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_50
timestamp 1644511149
transform 1 0 5704 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1644511149
transform 1 0 6256 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1644511149
transform 1 0 7360 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_80
timestamp 1644511149
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_144
timestamp 1644511149
transform 1 0 14352 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_152
timestamp 1644511149
transform 1 0 15088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_175
timestamp 1644511149
transform 1 0 17204 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_181
timestamp 1644511149
transform 1 0 17756 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_188
timestamp 1644511149
transform 1 0 18400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_200
timestamp 1644511149
transform 1 0 19504 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_206
timestamp 1644511149
transform 1 0 20056 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_217
timestamp 1644511149
transform 1 0 21068 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_231
timestamp 1644511149
transform 1 0 22356 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_238
timestamp 1644511149
transform 1 0 23000 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_244
timestamp 1644511149
transform 1 0 23552 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_256
timestamp 1644511149
transform 1 0 24656 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_262
timestamp 1644511149
transform 1 0 25208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_272
timestamp 1644511149
transform 1 0 26128 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1644511149
transform 1 0 26496 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_280
timestamp 1644511149
transform 1 0 26864 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_294
timestamp 1644511149
transform 1 0 28152 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1644511149
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_343
timestamp 1644511149
transform 1 0 32660 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_349
timestamp 1644511149
transform 1 0 33212 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_355
timestamp 1644511149
transform 1 0 33764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_37
timestamp 1644511149
transform 1 0 4508 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_41
timestamp 1644511149
transform 1 0 4876 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1644511149
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_59
timestamp 1644511149
transform 1 0 6532 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_71
timestamp 1644511149
transform 1 0 7636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_83
timestamp 1644511149
transform 1 0 8740 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_87
timestamp 1644511149
transform 1 0 9108 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_91
timestamp 1644511149
transform 1 0 9476 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_101
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1644511149
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_177
timestamp 1644511149
transform 1 0 17388 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_183
timestamp 1644511149
transform 1 0 17940 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_189
timestamp 1644511149
transform 1 0 18492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_201
timestamp 1644511149
transform 1 0 19596 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_219
timestamp 1644511149
transform 1 0 21252 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_231
timestamp 1644511149
transform 1 0 22356 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_259
timestamp 1644511149
transform 1 0 24932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_263
timestamp 1644511149
transform 1 0 25300 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_270
timestamp 1644511149
transform 1 0 25944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_287
timestamp 1644511149
transform 1 0 27508 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_316
timestamp 1644511149
transform 1 0 30176 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_324
timestamp 1644511149
transform 1 0 30912 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1644511149
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_343
timestamp 1644511149
transform 1 0 32660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_5
timestamp 1644511149
transform 1 0 1564 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_13
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_17
timestamp 1644511149
transform 1 0 2668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1644511149
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_36
timestamp 1644511149
transform 1 0 4416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_61
timestamp 1644511149
transform 1 0 6716 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_73
timestamp 1644511149
transform 1 0 7820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1644511149
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_106
timestamp 1644511149
transform 1 0 10856 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_116
timestamp 1644511149
transform 1 0 11776 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_128
timestamp 1644511149
transform 1 0 12880 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_200
timestamp 1644511149
transform 1 0 19504 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_212
timestamp 1644511149
transform 1 0 20608 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_220
timestamp 1644511149
transform 1 0 21344 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_228
timestamp 1644511149
transform 1 0 22080 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_236
timestamp 1644511149
transform 1 0 22816 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_257
timestamp 1644511149
transform 1 0 24748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_260
timestamp 1644511149
transform 1 0 25024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_270
timestamp 1644511149
transform 1 0 25944 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_280
timestamp 1644511149
transform 1 0 26864 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_288
timestamp 1644511149
transform 1 0 27600 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1644511149
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_314
timestamp 1644511149
transform 1 0 29992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_328
timestamp 1644511149
transform 1 0 31280 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_341
timestamp 1644511149
transform 1 0 32476 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_352
timestamp 1644511149
transform 1 0 33488 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_358
timestamp 1644511149
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_382
timestamp 1644511149
transform 1 0 36248 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_394
timestamp 1644511149
transform 1 0 37352 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1644511149
transform 1 0 38456 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_6
timestamp 1644511149
transform 1 0 1656 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_22
timestamp 1644511149
transform 1 0 3128 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_40
timestamp 1644511149
transform 1 0 4784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1644511149
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_60
timestamp 1644511149
transform 1 0 6624 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_72
timestamp 1644511149
transform 1 0 7728 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_84
timestamp 1644511149
transform 1 0 8832 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_91
timestamp 1644511149
transform 1 0 9476 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_101
timestamp 1644511149
transform 1 0 10396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1644511149
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_116
timestamp 1644511149
transform 1 0 11776 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_123
timestamp 1644511149
transform 1 0 12420 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_131
timestamp 1644511149
transform 1 0 13156 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_135
timestamp 1644511149
transform 1 0 13524 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_160
timestamp 1644511149
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_233
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_242
timestamp 1644511149
transform 1 0 23368 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_254
timestamp 1644511149
transform 1 0 24472 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_264
timestamp 1644511149
transform 1 0 25392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_270
timestamp 1644511149
transform 1 0 25944 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_291
timestamp 1644511149
transform 1 0 27876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_303
timestamp 1644511149
transform 1 0 28980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_327
timestamp 1644511149
transform 1 0 31188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_347
timestamp 1644511149
transform 1 0 33028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_353
timestamp 1644511149
transform 1 0 33580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_365
timestamp 1644511149
transform 1 0 34684 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_375
timestamp 1644511149
transform 1 0 35604 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1644511149
transform 1 0 36800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_399
timestamp 1644511149
transform 1 0 37812 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_40
timestamp 1644511149
transform 1 0 4784 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1644511149
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_108
timestamp 1644511149
transform 1 0 11040 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_145
timestamp 1644511149
transform 1 0 14444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_159
timestamp 1644511149
transform 1 0 15732 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_169
timestamp 1644511149
transform 1 0 16652 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_175
timestamp 1644511149
transform 1 0 17204 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_185
timestamp 1644511149
transform 1 0 18124 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_218
timestamp 1644511149
transform 1 0 21160 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_230
timestamp 1644511149
transform 1 0 22264 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_242
timestamp 1644511149
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1644511149
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_269
timestamp 1644511149
transform 1 0 25852 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_272
timestamp 1644511149
transform 1 0 26128 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_276
timestamp 1644511149
transform 1 0 26496 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_279
timestamp 1644511149
transform 1 0 26772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_287
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1644511149
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_330
timestamp 1644511149
transform 1 0 31464 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_343
timestamp 1644511149
transform 1 0 32660 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1644511149
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_380
timestamp 1644511149
transform 1 0 36064 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_393
timestamp 1644511149
transform 1 0 37260 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_403
timestamp 1644511149
transform 1 0 38180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_6
timestamp 1644511149
transform 1 0 1656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_12
timestamp 1644511149
transform 1 0 2208 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_24
timestamp 1644511149
transform 1 0 3312 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_36
timestamp 1644511149
transform 1 0 4416 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_40
timestamp 1644511149
transform 1 0 4784 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_47
timestamp 1644511149
transform 1 0 5428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_95
timestamp 1644511149
transform 1 0 9844 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1644511149
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_185
timestamp 1644511149
transform 1 0 18124 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_210
timestamp 1644511149
transform 1 0 20424 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1644511149
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_245
timestamp 1644511149
transform 1 0 23644 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_254
timestamp 1644511149
transform 1 0 24472 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_266
timestamp 1644511149
transform 1 0 25576 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1644511149
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_289
timestamp 1644511149
transform 1 0 27692 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_313
timestamp 1644511149
transform 1 0 29900 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_325
timestamp 1644511149
transform 1 0 31004 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_345
timestamp 1644511149
transform 1 0 32844 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_362
timestamp 1644511149
transform 1 0 34408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_368
timestamp 1644511149
transform 1 0 34960 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_376
timestamp 1644511149
transform 1 0 35696 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1644511149
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_401
timestamp 1644511149
transform 1 0 37996 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1644511149
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_35
timestamp 1644511149
transform 1 0 4324 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_47
timestamp 1644511149
transform 1 0 5428 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_59
timestamp 1644511149
transform 1 0 6532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_71
timestamp 1644511149
transform 1 0 7636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_96
timestamp 1644511149
transform 1 0 9936 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_103
timestamp 1644511149
transform 1 0 10580 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_110
timestamp 1644511149
transform 1 0 11224 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_122
timestamp 1644511149
transform 1 0 12328 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 1644511149
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_145
timestamp 1644511149
transform 1 0 14444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_167
timestamp 1644511149
transform 1 0 16468 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_181
timestamp 1644511149
transform 1 0 17756 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_185
timestamp 1644511149
transform 1 0 18124 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_201
timestamp 1644511149
transform 1 0 19596 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_206
timestamp 1644511149
transform 1 0 20056 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_220
timestamp 1644511149
transform 1 0 21344 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_232
timestamp 1644511149
transform 1 0 22448 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_244
timestamp 1644511149
transform 1 0 23552 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_274
timestamp 1644511149
transform 1 0 26312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_288
timestamp 1644511149
transform 1 0 27600 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_300
timestamp 1644511149
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_338
timestamp 1644511149
transform 1 0 32200 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_350
timestamp 1644511149
transform 1 0 33304 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_369
timestamp 1644511149
transform 1 0 35052 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_379
timestamp 1644511149
transform 1 0 35972 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_392
timestamp 1644511149
transform 1 0 37168 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_404
timestamp 1644511149
transform 1 0 38272 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_5
timestamp 1644511149
transform 1 0 1564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_17
timestamp 1644511149
transform 1 0 2668 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_46
timestamp 1644511149
transform 1 0 5336 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1644511149
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1644511149
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_135
timestamp 1644511149
transform 1 0 13524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_144
timestamp 1644511149
transform 1 0 14352 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_151
timestamp 1644511149
transform 1 0 14996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_172
timestamp 1644511149
transform 1 0 16928 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1644511149
transform 1 0 18032 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_196
timestamp 1644511149
transform 1 0 19136 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_209
timestamp 1644511149
transform 1 0 20332 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_215
timestamp 1644511149
transform 1 0 20884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_266
timestamp 1644511149
transform 1 0 25576 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_291
timestamp 1644511149
transform 1 0 27876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_303
timestamp 1644511149
transform 1 0 28980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_309
timestamp 1644511149
transform 1 0 29532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_319
timestamp 1644511149
transform 1 0 30452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_331
timestamp 1644511149
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_345
timestamp 1644511149
transform 1 0 32844 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_353
timestamp 1644511149
transform 1 0 33580 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_360
timestamp 1644511149
transform 1 0 34224 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_372
timestamp 1644511149
transform 1 0 35328 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1644511149
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_6
timestamp 1644511149
transform 1 0 1656 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_17
timestamp 1644511149
transform 1 0 2668 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_37
timestamp 1644511149
transform 1 0 4508 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_43
timestamp 1644511149
transform 1 0 5060 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_51
timestamp 1644511149
transform 1 0 5796 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_63
timestamp 1644511149
transform 1 0 6900 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_75
timestamp 1644511149
transform 1 0 8004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_106
timestamp 1644511149
transform 1 0 10856 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_118
timestamp 1644511149
transform 1 0 11960 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_122
timestamp 1644511149
transform 1 0 12328 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_151
timestamp 1644511149
transform 1 0 14996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_163
timestamp 1644511149
transform 1 0 16100 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_175
timestamp 1644511149
transform 1 0 17204 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_187
timestamp 1644511149
transform 1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_229
timestamp 1644511149
transform 1 0 22172 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_234
timestamp 1644511149
transform 1 0 22632 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1644511149
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_259
timestamp 1644511149
transform 1 0 24932 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_266
timestamp 1644511149
transform 1 0 25576 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_278
timestamp 1644511149
transform 1 0 26680 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_290
timestamp 1644511149
transform 1 0 27784 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1644511149
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_318
timestamp 1644511149
transform 1 0 30360 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_324
timestamp 1644511149
transform 1 0 30912 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_327
timestamp 1644511149
transform 1 0 31188 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_339
timestamp 1644511149
transform 1 0 32292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_351
timestamp 1644511149
transform 1 0 33396 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_356
timestamp 1644511149
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_22
timestamp 1644511149
transform 1 0 3128 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1644511149
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_77
timestamp 1644511149
transform 1 0 8188 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_83
timestamp 1644511149
transform 1 0 8740 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_87
timestamp 1644511149
transform 1 0 9108 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_91
timestamp 1644511149
transform 1 0 9476 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_103
timestamp 1644511149
transform 1 0 10580 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_116
timestamp 1644511149
transform 1 0 11776 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_141
timestamp 1644511149
transform 1 0 14076 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_155
timestamp 1644511149
transform 1 0 15364 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1644511149
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_177
timestamp 1644511149
transform 1 0 17388 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_183
timestamp 1644511149
transform 1 0 17940 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_188
timestamp 1644511149
transform 1 0 18400 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_202
timestamp 1644511149
transform 1 0 19688 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_209
timestamp 1644511149
transform 1 0 20332 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_215
timestamp 1644511149
transform 1 0 20884 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_239
timestamp 1644511149
transform 1 0 23092 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_246
timestamp 1644511149
transform 1 0 23736 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_253
timestamp 1644511149
transform 1 0 24380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_265
timestamp 1644511149
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1644511149
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_285
timestamp 1644511149
transform 1 0 27324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_307
timestamp 1644511149
transform 1 0 29348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_320
timestamp 1644511149
transform 1 0 30544 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_326
timestamp 1644511149
transform 1 0 31096 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1644511149
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_6
timestamp 1644511149
transform 1 0 1656 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_12
timestamp 1644511149
transform 1 0 2208 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1644511149
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_36
timestamp 1644511149
transform 1 0 4416 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_48
timestamp 1644511149
transform 1 0 5520 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_60
timestamp 1644511149
transform 1 0 6624 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_68
timestamp 1644511149
transform 1 0 7360 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_72
timestamp 1644511149
transform 1 0 7728 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_93
timestamp 1644511149
transform 1 0 9660 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_105
timestamp 1644511149
transform 1 0 10764 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_113
timestamp 1644511149
transform 1 0 11500 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_117
timestamp 1644511149
transform 1 0 11868 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_131
timestamp 1644511149
transform 1 0 13156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_143
timestamp 1644511149
transform 1 0 14260 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_151
timestamp 1644511149
transform 1 0 14996 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_154
timestamp 1644511149
transform 1 0 15272 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_168
timestamp 1644511149
transform 1 0 16560 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_174
timestamp 1644511149
transform 1 0 17112 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_185
timestamp 1644511149
transform 1 0 18124 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1644511149
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_214
timestamp 1644511149
transform 1 0 20792 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_226
timestamp 1644511149
transform 1 0 21896 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_236
timestamp 1644511149
transform 1 0 22816 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_243
timestamp 1644511149
transform 1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1644511149
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_313
timestamp 1644511149
transform 1 0 29900 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_319
timestamp 1644511149
transform 1 0 30452 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_324
timestamp 1644511149
transform 1 0 30912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_332
timestamp 1644511149
transform 1 0 31648 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_335
timestamp 1644511149
transform 1 0 31924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_341
timestamp 1644511149
transform 1 0 32476 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_353
timestamp 1644511149
transform 1 0 33580 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_361
timestamp 1644511149
transform 1 0 34316 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_370
timestamp 1644511149
transform 1 0 35144 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_378
timestamp 1644511149
transform 1 0 35880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_390
timestamp 1644511149
transform 1 0 36984 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1644511149
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_36
timestamp 1644511149
transform 1 0 4416 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_46
timestamp 1644511149
transform 1 0 5336 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1644511149
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_90
timestamp 1644511149
transform 1 0 9384 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_102
timestamp 1644511149
transform 1 0 10488 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1644511149
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_117
timestamp 1644511149
transform 1 0 11868 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_124
timestamp 1644511149
transform 1 0 12512 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_130
timestamp 1644511149
transform 1 0 13064 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_135
timestamp 1644511149
transform 1 0 13524 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_143
timestamp 1644511149
transform 1 0 14260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_151
timestamp 1644511149
transform 1 0 14996 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_163
timestamp 1644511149
transform 1 0 16100 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_177
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_188
timestamp 1644511149
transform 1 0 18400 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_198
timestamp 1644511149
transform 1 0 19320 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_204
timestamp 1644511149
transform 1 0 19872 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_213
timestamp 1644511149
transform 1 0 20700 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1644511149
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_230
timestamp 1644511149
transform 1 0 22264 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_255
timestamp 1644511149
transform 1 0 24564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_267
timestamp 1644511149
transform 1 0 25668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_297
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_300
timestamp 1644511149
transform 1 0 28704 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_311
timestamp 1644511149
transform 1 0 29716 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_315
timestamp 1644511149
transform 1 0 30084 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_326
timestamp 1644511149
transform 1 0 31096 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_342
timestamp 1644511149
transform 1 0 32568 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_354
timestamp 1644511149
transform 1 0 33672 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_366
timestamp 1644511149
transform 1 0 34776 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_370
timestamp 1644511149
transform 1 0 35144 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1644511149
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_399
timestamp 1644511149
transform 1 0 37812 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1644511149
transform 1 0 38180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_5
timestamp 1644511149
transform 1 0 1564 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_17
timestamp 1644511149
transform 1 0 2668 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1644511149
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_50
timestamp 1644511149
transform 1 0 5704 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_62
timestamp 1644511149
transform 1 0 6808 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_66
timestamp 1644511149
transform 1 0 7176 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_70
timestamp 1644511149
transform 1 0 7544 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1644511149
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_91
timestamp 1644511149
transform 1 0 9476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_101
timestamp 1644511149
transform 1 0 10396 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_130
timestamp 1644511149
transform 1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1644511149
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_149
timestamp 1644511149
transform 1 0 14812 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_156
timestamp 1644511149
transform 1 0 15456 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_170
timestamp 1644511149
transform 1 0 16744 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_184
timestamp 1644511149
transform 1 0 18032 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1644511149
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_203
timestamp 1644511149
transform 1 0 19780 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_211
timestamp 1644511149
transform 1 0 20516 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_218
timestamp 1644511149
transform 1 0 21160 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_228
timestamp 1644511149
transform 1 0 22080 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_234
timestamp 1644511149
transform 1 0 22632 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_238
timestamp 1644511149
transform 1 0 23000 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_259
timestamp 1644511149
transform 1 0 24932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_293
timestamp 1644511149
transform 1 0 28060 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_318
timestamp 1644511149
transform 1 0 30360 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_331
timestamp 1644511149
transform 1 0 31556 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_342
timestamp 1644511149
transform 1 0 32568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_346
timestamp 1644511149
transform 1 0 32936 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_356
timestamp 1644511149
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_376
timestamp 1644511149
transform 1 0 35696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_388
timestamp 1644511149
transform 1 0 36800 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_400
timestamp 1644511149
transform 1 0 37904 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1644511149
transform 1 0 38456 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_6
timestamp 1644511149
transform 1 0 1656 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_14
timestamp 1644511149
transform 1 0 2392 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_24
timestamp 1644511149
transform 1 0 3312 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_31
timestamp 1644511149
transform 1 0 3956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_38
timestamp 1644511149
transform 1 0 4600 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1644511149
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_63
timestamp 1644511149
transform 1 0 6900 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_88
timestamp 1644511149
transform 1 0 9200 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_100
timestamp 1644511149
transform 1 0 10304 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1644511149
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_123
timestamp 1644511149
transform 1 0 12420 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_148
timestamp 1644511149
transform 1 0 14720 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_160
timestamp 1644511149
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_177
timestamp 1644511149
transform 1 0 17388 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_183
timestamp 1644511149
transform 1 0 17940 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_231
timestamp 1644511149
transform 1 0 22356 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_239
timestamp 1644511149
transform 1 0 23092 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_262
timestamp 1644511149
transform 1 0 25208 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_272
timestamp 1644511149
transform 1 0 26128 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_314
timestamp 1644511149
transform 1 0 29992 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_318
timestamp 1644511149
transform 1 0 30360 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_321
timestamp 1644511149
transform 1 0 30636 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_350
timestamp 1644511149
transform 1 0 33304 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_358
timestamp 1644511149
transform 1 0 34040 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_364
timestamp 1644511149
transform 1 0 34592 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_370
timestamp 1644511149
transform 1 0 35144 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1644511149
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_22
timestamp 1644511149
transform 1 0 3128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_52
timestamp 1644511149
transform 1 0 5888 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_56
timestamp 1644511149
transform 1 0 6256 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_67
timestamp 1644511149
transform 1 0 7268 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_79
timestamp 1644511149
transform 1 0 8372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_123
timestamp 1644511149
transform 1 0 12420 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_130
timestamp 1644511149
transform 1 0 13064 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1644511149
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_144
timestamp 1644511149
transform 1 0 14352 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_159
timestamp 1644511149
transform 1 0 15732 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_184
timestamp 1644511149
transform 1 0 18032 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_200
timestamp 1644511149
transform 1 0 19504 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_212
timestamp 1644511149
transform 1 0 20608 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_224
timestamp 1644511149
transform 1 0 21712 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_236
timestamp 1644511149
transform 1 0 22816 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_244
timestamp 1644511149
transform 1 0 23552 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1644511149
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_259
timestamp 1644511149
transform 1 0 24932 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_263
timestamp 1644511149
transform 1 0 25300 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_266
timestamp 1644511149
transform 1 0 25576 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_278
timestamp 1644511149
transform 1 0 26680 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_290
timestamp 1644511149
transform 1 0 27784 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_302
timestamp 1644511149
transform 1 0 28888 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_318
timestamp 1644511149
transform 1 0 30360 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_324
timestamp 1644511149
transform 1 0 30912 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_332
timestamp 1644511149
transform 1 0 31648 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_342
timestamp 1644511149
transform 1 0 32568 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_355
timestamp 1644511149
transform 1 0 33764 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_381
timestamp 1644511149
transform 1 0 36156 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_398
timestamp 1644511149
transform 1 0 37720 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1644511149
transform 1 0 38456 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_6
timestamp 1644511149
transform 1 0 1656 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_12
timestamp 1644511149
transform 1 0 2208 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_18
timestamp 1644511149
transform 1 0 2760 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_40
timestamp 1644511149
transform 1 0 4784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_47
timestamp 1644511149
transform 1 0 5428 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_65
timestamp 1644511149
transform 1 0 7084 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_87
timestamp 1644511149
transform 1 0 9108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_99
timestamp 1644511149
transform 1 0 10212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_121
timestamp 1644511149
transform 1 0 12236 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_144
timestamp 1644511149
transform 1 0 14352 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_156
timestamp 1644511149
transform 1 0 15456 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_187
timestamp 1644511149
transform 1 0 18308 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_194
timestamp 1644511149
transform 1 0 18952 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_200
timestamp 1644511149
transform 1 0 19504 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_212
timestamp 1644511149
transform 1 0 20608 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_241
timestamp 1644511149
transform 1 0 23276 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_252
timestamp 1644511149
transform 1 0 24288 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_267
timestamp 1644511149
transform 1 0 25668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_39
timestamp 1644511149
transform 1 0 4692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_51
timestamp 1644511149
transform 1 0 5796 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_63
timestamp 1644511149
transform 1 0 6900 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_69
timestamp 1644511149
transform 1 0 7452 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_73
timestamp 1644511149
transform 1 0 7820 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_81
timestamp 1644511149
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_118
timestamp 1644511149
transform 1 0 11960 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_122
timestamp 1644511149
transform 1 0 12328 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_126
timestamp 1644511149
transform 1 0 12696 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1644511149
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_151
timestamp 1644511149
transform 1 0 14996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_157
timestamp 1644511149
transform 1 0 15548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_169
timestamp 1644511149
transform 1 0 16652 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_176
timestamp 1644511149
transform 1 0 17296 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_184
timestamp 1644511149
transform 1 0 18032 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_188
timestamp 1644511149
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_199
timestamp 1644511149
transform 1 0 19412 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_205
timestamp 1644511149
transform 1 0 19964 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_217
timestamp 1644511149
transform 1 0 21068 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_229
timestamp 1644511149
transform 1 0 22172 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_243
timestamp 1644511149
transform 1 0 23460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_258
timestamp 1644511149
transform 1 0 24840 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_287
timestamp 1644511149
transform 1 0 27508 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_299
timestamp 1644511149
transform 1 0 28612 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_66
timestamp 1644511149
transform 1 0 7176 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_76
timestamp 1644511149
transform 1 0 8096 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_88
timestamp 1644511149
transform 1 0 9200 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_96
timestamp 1644511149
transform 1 0 9936 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_102
timestamp 1644511149
transform 1 0 10488 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1644511149
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_116
timestamp 1644511149
transform 1 0 11776 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_130
timestamp 1644511149
transform 1 0 13064 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_142
timestamp 1644511149
transform 1 0 14168 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_154
timestamp 1644511149
transform 1 0 15272 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_179
timestamp 1644511149
transform 1 0 17572 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_187
timestamp 1644511149
transform 1 0 18308 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_194
timestamp 1644511149
transform 1 0 18952 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_204
timestamp 1644511149
transform 1 0 19872 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_210
timestamp 1644511149
transform 1 0 20424 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1644511149
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_253
timestamp 1644511149
transform 1 0 24380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1644511149
transform 1 0 26404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_284
timestamp 1644511149
transform 1 0 27232 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_296
timestamp 1644511149
transform 1 0 28336 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_308
timestamp 1644511149
transform 1 0 29440 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_320
timestamp 1644511149
transform 1 0 30544 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1644511149
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_342
timestamp 1644511149
transform 1 0 32568 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_354
timestamp 1644511149
transform 1 0 33672 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_366
timestamp 1644511149
transform 1 0 34776 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_378
timestamp 1644511149
transform 1 0 35880 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1644511149
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_12
timestamp 1644511149
transform 1 0 2208 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1644511149
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_35
timestamp 1644511149
transform 1 0 4324 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_57
timestamp 1644511149
transform 1 0 6348 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_73
timestamp 1644511149
transform 1 0 7820 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_81
timestamp 1644511149
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_112
timestamp 1644511149
transform 1 0 11408 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_126
timestamp 1644511149
transform 1 0 12696 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_159
timestamp 1644511149
transform 1 0 15732 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_166
timestamp 1644511149
transform 1 0 16376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_172
timestamp 1644511149
transform 1 0 16928 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_182
timestamp 1644511149
transform 1 0 17848 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1644511149
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_203
timestamp 1644511149
transform 1 0 19780 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_211
timestamp 1644511149
transform 1 0 20516 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_216
timestamp 1644511149
transform 1 0 20976 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_224
timestamp 1644511149
transform 1 0 21712 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_228
timestamp 1644511149
transform 1 0 22080 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_243
timestamp 1644511149
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_281
timestamp 1644511149
transform 1 0 26956 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_295
timestamp 1644511149
transform 1 0 28244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_316
timestamp 1644511149
transform 1 0 30176 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_325
timestamp 1644511149
transform 1 0 31004 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_329
timestamp 1644511149
transform 1 0 31372 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_335
timestamp 1644511149
transform 1 0 31924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_346
timestamp 1644511149
transform 1 0 32936 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_358
timestamp 1644511149
transform 1 0 34040 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_393
timestamp 1644511149
transform 1 0 37260 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_396
timestamp 1644511149
transform 1 0 37536 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_403
timestamp 1644511149
transform 1 0 38180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_18
timestamp 1644511149
transform 1 0 2760 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_43
timestamp 1644511149
transform 1 0 5060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1644511149
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_67
timestamp 1644511149
transform 1 0 7268 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_77
timestamp 1644511149
transform 1 0 8188 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_89
timestamp 1644511149
transform 1 0 9292 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_101
timestamp 1644511149
transform 1 0 10396 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_109
timestamp 1644511149
transform 1 0 11132 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_119
timestamp 1644511149
transform 1 0 12052 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_129
timestamp 1644511149
transform 1 0 12972 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_136
timestamp 1644511149
transform 1 0 13616 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_148
timestamp 1644511149
transform 1 0 14720 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_160
timestamp 1644511149
transform 1 0 15824 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_175
timestamp 1644511149
transform 1 0 17204 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_185
timestamp 1644511149
transform 1 0 18124 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_195
timestamp 1644511149
transform 1 0 19044 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_201
timestamp 1644511149
transform 1 0 19596 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_213
timestamp 1644511149
transform 1 0 20700 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_219
timestamp 1644511149
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_246
timestamp 1644511149
transform 1 0 23736 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_309
timestamp 1644511149
transform 1 0 29532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_313
timestamp 1644511149
transform 1 0 29900 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_320
timestamp 1644511149
transform 1 0 30544 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1644511149
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_345
timestamp 1644511149
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_362
timestamp 1644511149
transform 1 0 34408 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_374
timestamp 1644511149
transform 1 0 35512 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_386
timestamp 1644511149
transform 1 0 36616 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_24
timestamp 1644511149
transform 1 0 3312 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_32
timestamp 1644511149
transform 1 0 4048 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_57
timestamp 1644511149
transform 1 0 6348 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_71
timestamp 1644511149
transform 1 0 7636 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_78
timestamp 1644511149
transform 1 0 8280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_108
timestamp 1644511149
transform 1 0 11040 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_122
timestamp 1644511149
transform 1 0 12328 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_132
timestamp 1644511149
transform 1 0 13248 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_162
timestamp 1644511149
transform 1 0 16008 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_172
timestamp 1644511149
transform 1 0 16928 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_180
timestamp 1644511149
transform 1 0 17664 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_187
timestamp 1644511149
transform 1 0 18308 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_225
timestamp 1644511149
transform 1 0 21804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_247
timestamp 1644511149
transform 1 0 23828 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_263
timestamp 1644511149
transform 1 0 25300 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_272
timestamp 1644511149
transform 1 0 26128 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_299
timestamp 1644511149
transform 1 0 28612 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_325
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_338
timestamp 1644511149
transform 1 0 32200 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_350
timestamp 1644511149
transform 1 0 33304 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1644511149
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_21
timestamp 1644511149
transform 1 0 3036 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_46
timestamp 1644511149
transform 1 0 5336 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_91
timestamp 1644511149
transform 1 0 9476 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_100
timestamp 1644511149
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_119
timestamp 1644511149
transform 1 0 12052 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_144
timestamp 1644511149
transform 1 0 14352 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_156
timestamp 1644511149
transform 1 0 15456 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_160
timestamp 1644511149
transform 1 0 15824 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1644511149
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_190
timestamp 1644511149
transform 1 0 18584 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_198
timestamp 1644511149
transform 1 0 19320 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_203
timestamp 1644511149
transform 1 0 19780 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_211
timestamp 1644511149
transform 1 0 20516 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_215
timestamp 1644511149
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_228
timestamp 1644511149
transform 1 0 22080 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_235
timestamp 1644511149
transform 1 0 22724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_260
timestamp 1644511149
transform 1 0 25024 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_272
timestamp 1644511149
transform 1 0 26128 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_302
timestamp 1644511149
transform 1 0 28888 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_330
timestamp 1644511149
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_353
timestamp 1644511149
transform 1 0 33580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_365
timestamp 1644511149
transform 1 0 34684 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_377
timestamp 1644511149
transform 1 0 35788 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_389
timestamp 1644511149
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_50
timestamp 1644511149
transform 1 0 5704 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_62
timestamp 1644511149
transform 1 0 6808 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_70
timestamp 1644511149
transform 1 0 7544 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_74
timestamp 1644511149
transform 1 0 7912 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1644511149
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_106
timestamp 1644511149
transform 1 0 10856 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_114
timestamp 1644511149
transform 1 0 11592 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_119
timestamp 1644511149
transform 1 0 12052 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_129
timestamp 1644511149
transform 1 0 12972 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1644511149
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_144
timestamp 1644511149
transform 1 0 14352 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_156
timestamp 1644511149
transform 1 0 15456 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_163
timestamp 1644511149
transform 1 0 16100 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_175
timestamp 1644511149
transform 1 0 17204 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_179
timestamp 1644511149
transform 1 0 17572 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_186
timestamp 1644511149
transform 1 0 18216 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1644511149
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_220
timestamp 1644511149
transform 1 0 21344 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_256
timestamp 1644511149
transform 1 0 24656 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_262
timestamp 1644511149
transform 1 0 25208 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_266
timestamp 1644511149
transform 1 0 25576 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_273
timestamp 1644511149
transform 1 0 26220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_298
timestamp 1644511149
transform 1 0 28520 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1644511149
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_21
timestamp 1644511149
transform 1 0 3036 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_25
timestamp 1644511149
transform 1 0 3404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_29
timestamp 1644511149
transform 1 0 3772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_33
timestamp 1644511149
transform 1 0 4140 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1644511149
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_77
timestamp 1644511149
transform 1 0 8188 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_83
timestamp 1644511149
transform 1 0 8740 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_90
timestamp 1644511149
transform 1 0 9384 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_102
timestamp 1644511149
transform 1 0 10488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1644511149
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_121
timestamp 1644511149
transform 1 0 12236 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_177
timestamp 1644511149
transform 1 0 17388 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_199
timestamp 1644511149
transform 1 0 19412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1644511149
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1644511149
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_284
timestamp 1644511149
transform 1 0 27232 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_296
timestamp 1644511149
transform 1 0 28336 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_308
timestamp 1644511149
transform 1 0 29440 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_314
timestamp 1644511149
transform 1 0 29992 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_326
timestamp 1644511149
transform 1 0 31096 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1644511149
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1644511149
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1644511149
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1644511149
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_181
timestamp 1644511149
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1644511149
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_237
timestamp 1644511149
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1644511149
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_293
timestamp 1644511149
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1644511149
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_313
timestamp 1644511149
transform 1 0 29900 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_318
timestamp 1644511149
transform 1 0 30360 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_330
timestamp 1644511149
transform 1 0 31464 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1644511149
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1644511149
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_393
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0726_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0727_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0728_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0729_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0730_
timestamp 1644511149
transform -1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0731_
timestamp 1644511149
transform 1 0 20148 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0732_
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1644511149
transform 1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0734_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0735_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0736_
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _0737_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2852 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0738_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18032 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0739_
timestamp 1644511149
transform 1 0 19688 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0740_
timestamp 1644511149
transform 1 0 22172 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1644511149
transform 1 0 3128 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0742_
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_2  _0743_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3128 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0744_
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0745_
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0746_
timestamp 1644511149
transform 1 0 16928 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0747_
timestamp 1644511149
transform -1 0 17296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0748_
timestamp 1644511149
transform -1 0 17204 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0749_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0750_
timestamp 1644511149
transform 1 0 17664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0751_
timestamp 1644511149
transform 1 0 18032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0752_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3404 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0753_
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0754_
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0755_
timestamp 1644511149
transform 1 0 2576 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0756_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4048 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0757_
timestamp 1644511149
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0758_
timestamp 1644511149
transform 1 0 19412 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0759_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0760_
timestamp 1644511149
transform -1 0 18124 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0761_
timestamp 1644511149
transform -1 0 17388 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0762_
timestamp 1644511149
transform -1 0 17204 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0763_
timestamp 1644511149
transform -1 0 16284 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0764_
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0765_
timestamp 1644511149
transform -1 0 20424 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0766_
timestamp 1644511149
transform -1 0 18216 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0767_
timestamp 1644511149
transform 1 0 17112 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0768_
timestamp 1644511149
transform -1 0 19136 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0769_
timestamp 1644511149
transform -1 0 18216 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0770_
timestamp 1644511149
transform 1 0 17204 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0771_
timestamp 1644511149
transform 1 0 18216 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0772_
timestamp 1644511149
transform -1 0 19780 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0773_
timestamp 1644511149
transform 1 0 17848 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0774_
timestamp 1644511149
transform -1 0 19504 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0775_
timestamp 1644511149
transform -1 0 17848 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0776_
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0777_
timestamp 1644511149
transform -1 0 13524 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0778_
timestamp 1644511149
transform -1 0 16008 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0779_
timestamp 1644511149
transform -1 0 14260 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0780_
timestamp 1644511149
transform 1 0 15640 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0781_
timestamp 1644511149
transform -1 0 16652 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0782_
timestamp 1644511149
transform 1 0 14720 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0783_
timestamp 1644511149
transform 1 0 18308 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0784_
timestamp 1644511149
transform -1 0 17388 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0785_
timestamp 1644511149
transform -1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0786_
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0787_
timestamp 1644511149
transform 1 0 16836 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0788_
timestamp 1644511149
transform -1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0789_
timestamp 1644511149
transform 1 0 15548 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0790_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0791_
timestamp 1644511149
transform -1 0 16376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0792_
timestamp 1644511149
transform 1 0 14444 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0793_
timestamp 1644511149
transform -1 0 15364 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0794_
timestamp 1644511149
transform -1 0 14996 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0795_
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0796_
timestamp 1644511149
transform -1 0 12696 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0797_
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0798_
timestamp 1644511149
transform -1 0 11960 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0799_
timestamp 1644511149
transform 1 0 11500 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0800_
timestamp 1644511149
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0801_
timestamp 1644511149
transform -1 0 10488 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0802_
timestamp 1644511149
transform 1 0 7636 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0803_
timestamp 1644511149
transform 1 0 8004 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0804_
timestamp 1644511149
transform -1 0 7820 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0805_
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0806_
timestamp 1644511149
transform -1 0 8096 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0807_
timestamp 1644511149
transform 1 0 7544 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0808_
timestamp 1644511149
transform -1 0 7268 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0809_
timestamp 1644511149
transform 1 0 6716 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0810_
timestamp 1644511149
transform 1 0 13340 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0811_
timestamp 1644511149
transform 1 0 13064 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0812_
timestamp 1644511149
transform -1 0 14996 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0813_
timestamp 1644511149
transform -1 0 12052 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0814_
timestamp 1644511149
transform 1 0 10028 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0815_
timestamp 1644511149
transform 1 0 12144 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0816_
timestamp 1644511149
transform -1 0 13248 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0817_
timestamp 1644511149
transform -1 0 12604 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0818_
timestamp 1644511149
transform -1 0 12972 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0819_
timestamp 1644511149
transform -1 0 12328 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0820_
timestamp 1644511149
transform 1 0 12420 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0821_
timestamp 1644511149
transform -1 0 13616 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0822_
timestamp 1644511149
transform -1 0 18308 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0823_
timestamp 1644511149
transform -1 0 12052 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0824_
timestamp 1644511149
transform -1 0 3312 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0825_
timestamp 1644511149
transform -1 0 16192 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0826_
timestamp 1644511149
transform -1 0 16376 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0827_
timestamp 1644511149
transform 1 0 17756 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0828_
timestamp 1644511149
transform -1 0 20884 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0829_
timestamp 1644511149
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0830_
timestamp 1644511149
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1644511149
transform 1 0 3128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0832_
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0833_
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0834_
timestamp 1644511149
transform 1 0 20424 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0835_
timestamp 1644511149
transform 1 0 22448 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0836_
timestamp 1644511149
transform 1 0 22816 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0837_
timestamp 1644511149
transform -1 0 25024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0838_
timestamp 1644511149
transform -1 0 16928 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0839_
timestamp 1644511149
transform 1 0 3864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0840_
timestamp 1644511149
transform -1 0 17204 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0841_
timestamp 1644511149
transform -1 0 16192 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0842_
timestamp 1644511149
transform -1 0 18400 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0843_
timestamp 1644511149
transform 1 0 17572 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0844_
timestamp 1644511149
transform 1 0 17940 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0845_
timestamp 1644511149
transform 1 0 18492 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0846_
timestamp 1644511149
transform -1 0 19780 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0847_
timestamp 1644511149
transform 1 0 23092 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0848_
timestamp 1644511149
transform 1 0 24564 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 1644511149
transform -1 0 17296 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0850_
timestamp 1644511149
transform -1 0 15732 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0851_
timestamp 1644511149
transform 1 0 18400 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0852_
timestamp 1644511149
transform -1 0 18952 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0853_
timestamp 1644511149
transform -1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0854_
timestamp 1644511149
transform 1 0 18216 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0855_
timestamp 1644511149
transform -1 0 26128 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0856_
timestamp 1644511149
transform 1 0 15088 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0857_
timestamp 1644511149
transform 1 0 17296 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0858_
timestamp 1644511149
transform -1 0 20976 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0859_
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0860_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0861_
timestamp 1644511149
transform 1 0 19320 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0862_
timestamp 1644511149
transform -1 0 21252 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0863_
timestamp 1644511149
transform 1 0 13524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0864_
timestamp 1644511149
transform -1 0 18584 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0865_
timestamp 1644511149
transform 1 0 12880 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0866_
timestamp 1644511149
transform -1 0 18584 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0867_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0868_
timestamp 1644511149
transform 1 0 19228 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0869_
timestamp 1644511149
transform 1 0 19872 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0870_
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0871_
timestamp 1644511149
transform 1 0 16744 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1644511149
transform -1 0 16928 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0873_
timestamp 1644511149
transform 1 0 19320 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0874_
timestamp 1644511149
transform -1 0 20608 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0875_
timestamp 1644511149
transform 1 0 15824 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0876_
timestamp 1644511149
transform 1 0 17296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0877_
timestamp 1644511149
transform -1 0 19596 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0878_
timestamp 1644511149
transform 1 0 19688 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0879_
timestamp 1644511149
transform -1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0880_
timestamp 1644511149
transform -1 0 19780 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1644511149
transform -1 0 20424 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0882_
timestamp 1644511149
transform 1 0 20516 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0883_
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0884_
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0885_
timestamp 1644511149
transform 1 0 23736 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0886_
timestamp 1644511149
transform -1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0887_
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0888_
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0889_
timestamp 1644511149
transform 1 0 21252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0890_
timestamp 1644511149
transform 1 0 22632 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0891_
timestamp 1644511149
transform -1 0 19688 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0892_
timestamp 1644511149
transform 1 0 19412 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 1644511149
transform 1 0 19688 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0894_
timestamp 1644511149
transform -1 0 19504 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1644511149
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0896_
timestamp 1644511149
transform 1 0 21252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0897_
timestamp 1644511149
transform -1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0898_
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0899_
timestamp 1644511149
transform -1 0 23276 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0900_
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1644511149
transform 1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0902_
timestamp 1644511149
transform -1 0 20424 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0903_
timestamp 1644511149
transform -1 0 14996 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0904_
timestamp 1644511149
transform 1 0 22172 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0905_
timestamp 1644511149
transform 1 0 23920 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0906_
timestamp 1644511149
transform -1 0 14444 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0907_
timestamp 1644511149
transform -1 0 14260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0908_
timestamp 1644511149
transform 1 0 14904 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0909_
timestamp 1644511149
transform 1 0 15272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0910_
timestamp 1644511149
transform -1 0 15916 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0912_
timestamp 1644511149
transform 1 0 14996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0913_
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0914_
timestamp 1644511149
transform -1 0 12604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0915_
timestamp 1644511149
transform -1 0 13524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0916_
timestamp 1644511149
transform 1 0 12696 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0917_
timestamp 1644511149
transform -1 0 11684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0918_
timestamp 1644511149
transform -1 0 12604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0919_
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0920_
timestamp 1644511149
transform 1 0 12420 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0921_
timestamp 1644511149
transform -1 0 13156 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0922_
timestamp 1644511149
transform -1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0923_
timestamp 1644511149
transform -1 0 9660 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0924_
timestamp 1644511149
transform -1 0 11316 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0925_
timestamp 1644511149
transform 1 0 10672 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0926_
timestamp 1644511149
transform -1 0 12236 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0927_
timestamp 1644511149
transform -1 0 12144 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0928_
timestamp 1644511149
transform -1 0 12420 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0929_
timestamp 1644511149
transform 1 0 10488 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0930_
timestamp 1644511149
transform -1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0932_
timestamp 1644511149
transform -1 0 11040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0933_
timestamp 1644511149
transform -1 0 10120 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0934_
timestamp 1644511149
transform 1 0 6900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0935_
timestamp 1644511149
transform 1 0 9384 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0936_
timestamp 1644511149
transform 1 0 7636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0937_
timestamp 1644511149
transform 1 0 9292 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0938_
timestamp 1644511149
transform -1 0 9752 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1644511149
transform 1 0 9016 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0940_
timestamp 1644511149
transform -1 0 10672 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0941_
timestamp 1644511149
transform -1 0 7360 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0942_
timestamp 1644511149
transform -1 0 10212 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1644511149
transform 1 0 9384 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0944_
timestamp 1644511149
transform 1 0 4600 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0945_
timestamp 1644511149
transform 1 0 8188 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0946_
timestamp 1644511149
transform 1 0 9292 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 1644511149
transform 1 0 10212 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0948_
timestamp 1644511149
transform 1 0 10120 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0949_
timestamp 1644511149
transform 1 0 27232 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0950_
timestamp 1644511149
transform -1 0 24656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 1644511149
transform -1 0 23920 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0952_
timestamp 1644511149
transform 1 0 25392 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0953_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0954_
timestamp 1644511149
transform 1 0 25392 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0955_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0956_
timestamp 1644511149
transform 1 0 5428 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0957_
timestamp 1644511149
transform 1 0 7544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0958_
timestamp 1644511149
transform 1 0 26312 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0959_
timestamp 1644511149
transform 1 0 26680 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0960_
timestamp 1644511149
transform 1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0961_
timestamp 1644511149
transform 1 0 25576 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0962_
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0963_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0964_
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0965_
timestamp 1644511149
transform -1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0966_
timestamp 1644511149
transform -1 0 7636 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _0967_
timestamp 1644511149
transform 1 0 7636 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0968_
timestamp 1644511149
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0969_
timestamp 1644511149
transform 1 0 7268 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0970_
timestamp 1644511149
transform 1 0 7544 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0971_
timestamp 1644511149
transform -1 0 5244 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0972_
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0973_
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0974_
timestamp 1644511149
transform 1 0 5336 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0975_
timestamp 1644511149
transform -1 0 5888 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0976_
timestamp 1644511149
transform -1 0 5428 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0977_
timestamp 1644511149
transform -1 0 6072 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0978_
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0979_
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0980_
timestamp 1644511149
transform 1 0 5612 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0981_
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0982_
timestamp 1644511149
transform -1 0 7544 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0983_
timestamp 1644511149
transform -1 0 4692 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 1644511149
transform 1 0 3128 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0985_
timestamp 1644511149
transform 1 0 4968 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1644511149
transform 1 0 5244 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0987_
timestamp 1644511149
transform 1 0 4784 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1644511149
transform 1 0 4600 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0989_
timestamp 1644511149
transform 1 0 3956 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1644511149
transform 1 0 5060 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0991_
timestamp 1644511149
transform -1 0 4508 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1644511149
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1644511149
transform 1 0 5428 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0994_
timestamp 1644511149
transform -1 0 5888 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0995_
timestamp 1644511149
transform -1 0 4416 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1644511149
transform 1 0 3036 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0997_
timestamp 1644511149
transform 1 0 3864 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1644511149
transform -1 0 5428 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0999_
timestamp 1644511149
transform 1 0 4232 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1644511149
transform 1 0 4508 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1644511149
transform 1 0 5060 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1003_
timestamp 1644511149
transform -1 0 4324 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1644511149
transform 1 0 3036 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1005_
timestamp 1644511149
transform -1 0 4508 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1644511149
transform -1 0 3312 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1007_
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1008_
timestamp 1644511149
transform -1 0 13340 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1009_
timestamp 1644511149
transform 1 0 13800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1010_
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1644511149
transform -1 0 4416 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1644511149
transform 1 0 3680 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1013_
timestamp 1644511149
transform -1 0 5336 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1644511149
transform 1 0 4324 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1015_
timestamp 1644511149
transform -1 0 4416 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1016_
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1017_
timestamp 1644511149
transform -1 0 18400 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1018_
timestamp 1644511149
transform 1 0 9292 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1019_
timestamp 1644511149
transform 1 0 11960 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1644511149
transform -1 0 13064 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1021_
timestamp 1644511149
transform 1 0 11868 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1644511149
transform -1 0 23736 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1024_
timestamp 1644511149
transform 1 0 23000 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1025_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1644511149
transform -1 0 25668 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1027_
timestamp 1644511149
transform -1 0 24932 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1028_
timestamp 1644511149
transform 1 0 24564 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1029_
timestamp 1644511149
transform 1 0 25576 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1030_
timestamp 1644511149
transform 1 0 26036 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1031_
timestamp 1644511149
transform -1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1032_
timestamp 1644511149
transform 1 0 22632 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1033_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1644511149
transform -1 0 23920 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1035_
timestamp 1644511149
transform 1 0 23920 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1644511149
transform -1 0 24380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1644511149
transform -1 0 23644 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1644511149
transform -1 0 23000 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1039_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1644511149
transform 1 0 25300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1041_
timestamp 1644511149
transform 1 0 24196 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1644511149
transform -1 0 26128 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1043_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1044_
timestamp 1644511149
transform 1 0 26036 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1644511149
transform -1 0 22080 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1046_
timestamp 1644511149
transform -1 0 22724 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1047_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1048_
timestamp 1644511149
transform -1 0 26036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1049_
timestamp 1644511149
transform 1 0 24104 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1050_
timestamp 1644511149
transform -1 0 26680 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1051_
timestamp 1644511149
transform -1 0 23184 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1052_
timestamp 1644511149
transform -1 0 22540 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1053_
timestamp 1644511149
transform 1 0 23368 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1054_
timestamp 1644511149
transform 1 0 25116 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1055_
timestamp 1644511149
transform 1 0 23092 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1056_
timestamp 1644511149
transform -1 0 25116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1057_
timestamp 1644511149
transform 1 0 22448 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1058_
timestamp 1644511149
transform 1 0 23184 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1059_
timestamp 1644511149
transform -1 0 12236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1060_
timestamp 1644511149
transform -1 0 12420 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1061_
timestamp 1644511149
transform 1 0 12420 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1062_
timestamp 1644511149
transform 1 0 12696 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1063_
timestamp 1644511149
transform 1 0 12604 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1064_
timestamp 1644511149
transform -1 0 5796 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1065_
timestamp 1644511149
transform 1 0 12696 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1066_
timestamp 1644511149
transform 1 0 12512 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1067_
timestamp 1644511149
transform 1 0 12052 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1644511149
transform -1 0 13432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1069_
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1070_
timestamp 1644511149
transform -1 0 13064 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1071_
timestamp 1644511149
transform 1 0 12604 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1644511149
transform -1 0 14352 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1073_
timestamp 1644511149
transform 1 0 10672 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1644511149
transform -1 0 9752 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1075_
timestamp 1644511149
transform 1 0 10948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1644511149
transform 1 0 11592 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1077_
timestamp 1644511149
transform 1 0 11868 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 1644511149
transform -1 0 11776 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1079_
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1080_
timestamp 1644511149
transform 1 0 12144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1081_
timestamp 1644511149
transform -1 0 10396 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1644511149
transform 1 0 9200 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1083_
timestamp 1644511149
transform 1 0 9844 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1084_
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1085_
timestamp 1644511149
transform -1 0 11776 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1644511149
transform -1 0 10672 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1087_
timestamp 1644511149
transform -1 0 10948 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1088_
timestamp 1644511149
transform 1 0 9844 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1089_
timestamp 1644511149
transform 1 0 9292 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1644511149
transform 1 0 10304 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1091_
timestamp 1644511149
transform -1 0 9476 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1092_
timestamp 1644511149
transform 1 0 9016 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1093_
timestamp 1644511149
transform -1 0 18400 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1644511149
transform -1 0 18124 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1095_
timestamp 1644511149
transform -1 0 9476 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1096_
timestamp 1644511149
transform -1 0 5888 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1097_
timestamp 1644511149
transform -1 0 8464 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1098_
timestamp 1644511149
transform -1 0 7544 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1099_
timestamp 1644511149
transform -1 0 10396 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1100_
timestamp 1644511149
transform -1 0 7268 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1101_
timestamp 1644511149
transform 1 0 18768 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1644511149
transform -1 0 20332 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1103_
timestamp 1644511149
transform -1 0 19780 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1104_
timestamp 1644511149
transform -1 0 18032 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1105_
timestamp 1644511149
transform -1 0 19320 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1644511149
transform -1 0 18952 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1107_
timestamp 1644511149
transform -1 0 20792 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1108_
timestamp 1644511149
transform -1 0 20700 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1109_
timestamp 1644511149
transform 1 0 21528 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1110_
timestamp 1644511149
transform 1 0 23368 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1111_
timestamp 1644511149
transform 1 0 20608 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1112_
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1113_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1114_
timestamp 1644511149
transform 1 0 27324 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1115_
timestamp 1644511149
transform 1 0 21344 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1116_
timestamp 1644511149
transform -1 0 22264 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1117_
timestamp 1644511149
transform 1 0 22264 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1118_
timestamp 1644511149
transform -1 0 23000 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1119_
timestamp 1644511149
transform 1 0 21528 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1120_
timestamp 1644511149
transform -1 0 23000 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1121_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1122_
timestamp 1644511149
transform -1 0 26864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1123_
timestamp 1644511149
transform 1 0 20056 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1124_
timestamp 1644511149
transform 1 0 20608 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1125_
timestamp 1644511149
transform -1 0 36616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1126_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34592 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1127_
timestamp 1644511149
transform -1 0 35052 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1128_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31832 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1129_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29808 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1130_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31280 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _1131_
timestamp 1644511149
transform 1 0 30452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1132_
timestamp 1644511149
transform -1 0 31740 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1644511149
transform -1 0 30912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1134_
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1135_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32752 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1136_
timestamp 1644511149
transform -1 0 32660 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1137_
timestamp 1644511149
transform -1 0 37996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1138_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36156 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1139_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35880 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1140_
timestamp 1644511149
transform 1 0 35144 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1141_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1142_
timestamp 1644511149
transform 1 0 17112 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_4  _1143_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20792 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _1144_
timestamp 1644511149
transform 1 0 31188 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1145_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25852 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1146_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32384 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1147_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33488 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1148_
timestamp 1644511149
transform -1 0 34224 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1149_
timestamp 1644511149
transform 1 0 30360 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1150_
timestamp 1644511149
transform -1 0 31096 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1151_
timestamp 1644511149
transform 1 0 30544 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1152_
timestamp 1644511149
transform 1 0 29624 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1153_
timestamp 1644511149
transform -1 0 33856 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1154_
timestamp 1644511149
transform -1 0 30360 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1155_
timestamp 1644511149
transform -1 0 32844 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1156_
timestamp 1644511149
transform 1 0 29900 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1157_
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1158_
timestamp 1644511149
transform -1 0 34592 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1159_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1160_
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1161_
timestamp 1644511149
transform 1 0 28428 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1162_
timestamp 1644511149
transform -1 0 30176 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1163_
timestamp 1644511149
transform -1 0 29900 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1164_
timestamp 1644511149
transform 1 0 30728 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1165_
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1166_
timestamp 1644511149
transform 1 0 29072 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1167_
timestamp 1644511149
transform -1 0 31004 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1168_
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1169_
timestamp 1644511149
transform 1 0 32476 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1170_
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1171_
timestamp 1644511149
transform 1 0 31004 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1172_
timestamp 1644511149
transform 1 0 31464 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1173_
timestamp 1644511149
transform -1 0 32200 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1174_
timestamp 1644511149
transform 1 0 33028 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1175_
timestamp 1644511149
transform 1 0 32936 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1176_
timestamp 1644511149
transform -1 0 32568 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1177_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1178_
timestamp 1644511149
transform -1 0 32936 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1179_
timestamp 1644511149
transform 1 0 30360 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1180_
timestamp 1644511149
transform 1 0 33580 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1181_
timestamp 1644511149
transform 1 0 33028 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1182_
timestamp 1644511149
transform 1 0 32200 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1183_
timestamp 1644511149
transform 1 0 33488 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1184_
timestamp 1644511149
transform -1 0 35144 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1185_
timestamp 1644511149
transform 1 0 23092 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1186_
timestamp 1644511149
transform 1 0 37352 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1187_
timestamp 1644511149
transform 1 0 35236 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1188_
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1189_
timestamp 1644511149
transform 1 0 33304 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1190_
timestamp 1644511149
transform -1 0 34592 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1191_
timestamp 1644511149
transform 1 0 36432 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1192_
timestamp 1644511149
transform 1 0 35972 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1193_
timestamp 1644511149
transform -1 0 36800 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1194_
timestamp 1644511149
transform 1 0 37076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1195_
timestamp 1644511149
transform 1 0 36340 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1196_
timestamp 1644511149
transform -1 0 32476 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1197_
timestamp 1644511149
transform 1 0 32016 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1198_
timestamp 1644511149
transform 1 0 33764 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1199_
timestamp 1644511149
transform -1 0 35696 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1200_
timestamp 1644511149
transform 1 0 2576 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1201_
timestamp 1644511149
transform 1 0 2944 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _1202_
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1203_
timestamp 1644511149
transform 1 0 29900 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1204_
timestamp 1644511149
transform 1 0 30452 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1205_
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1206_
timestamp 1644511149
transform 1 0 31464 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1207_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1208_
timestamp 1644511149
transform 1 0 29532 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1644511149
transform -1 0 30176 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1210_
timestamp 1644511149
transform 1 0 30912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1211_
timestamp 1644511149
transform -1 0 30360 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1212_
timestamp 1644511149
transform 1 0 30728 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1213_
timestamp 1644511149
transform -1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1214_
timestamp 1644511149
transform -1 0 30084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1215_
timestamp 1644511149
transform 1 0 27968 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1216_
timestamp 1644511149
transform -1 0 27600 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1217_
timestamp 1644511149
transform 1 0 27048 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1218_
timestamp 1644511149
transform 1 0 29992 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1219_
timestamp 1644511149
transform 1 0 30084 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1220_
timestamp 1644511149
transform -1 0 31464 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1221_
timestamp 1644511149
transform -1 0 31188 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 1644511149
transform 1 0 33764 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1644511149
transform -1 0 35512 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1224_
timestamp 1644511149
transform 1 0 30176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1225_
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1226_
timestamp 1644511149
transform -1 0 26128 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1227_
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1228_
timestamp 1644511149
transform 1 0 29716 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1229_
timestamp 1644511149
transform 1 0 28980 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1230_
timestamp 1644511149
transform 1 0 29808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1231_
timestamp 1644511149
transform 1 0 32660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1232_
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1233_
timestamp 1644511149
transform 1 0 32384 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1234_
timestamp 1644511149
transform 1 0 32292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1235_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 33212 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1236_
timestamp 1644511149
transform 1 0 35696 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1237_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35880 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1238_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35052 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1239_
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1240_
timestamp 1644511149
transform 1 0 37260 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 1644511149
transform -1 0 35512 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1242_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1243_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34868 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1244_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1245_
timestamp 1644511149
transform -1 0 35052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1246_
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1247_
timestamp 1644511149
transform 1 0 33764 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1248_
timestamp 1644511149
transform -1 0 34776 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _1249_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35512 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1250_
timestamp 1644511149
transform -1 0 33396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1251_
timestamp 1644511149
transform -1 0 33488 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1252_
timestamp 1644511149
transform -1 0 32476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1253_
timestamp 1644511149
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1254_
timestamp 1644511149
transform -1 0 17388 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1255_
timestamp 1644511149
transform 1 0 14904 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1256_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24104 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1257_
timestamp 1644511149
transform 1 0 14168 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _1258_
timestamp 1644511149
transform -1 0 18676 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _1259_
timestamp 1644511149
transform -1 0 17388 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1260_
timestamp 1644511149
transform -1 0 14720 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1261_
timestamp 1644511149
transform -1 0 14536 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1644511149
transform 1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1263_
timestamp 1644511149
transform 1 0 20424 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1264_
timestamp 1644511149
transform 1 0 11868 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1265_
timestamp 1644511149
transform 1 0 10120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1266_
timestamp 1644511149
transform -1 0 11040 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1267_
timestamp 1644511149
transform -1 0 20332 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1268_
timestamp 1644511149
transform 1 0 10488 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1269_
timestamp 1644511149
transform -1 0 11960 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1270_
timestamp 1644511149
transform -1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1271_
timestamp 1644511149
transform -1 0 26220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1272_
timestamp 1644511149
transform 1 0 8372 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1273_
timestamp 1644511149
transform 1 0 6440 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1274_
timestamp 1644511149
transform -1 0 5612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1275_
timestamp 1644511149
transform 1 0 4048 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1276_
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1277_
timestamp 1644511149
transform 1 0 6808 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1278_
timestamp 1644511149
transform 1 0 5336 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1279_
timestamp 1644511149
transform -1 0 4968 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1280_
timestamp 1644511149
transform -1 0 4232 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1281_
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1282_
timestamp 1644511149
transform 1 0 6164 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1283_
timestamp 1644511149
transform 1 0 4968 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1284_
timestamp 1644511149
transform -1 0 5060 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1285_
timestamp 1644511149
transform -1 0 4048 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1286_
timestamp 1644511149
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1287_
timestamp 1644511149
transform 1 0 6900 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1288_
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1289_
timestamp 1644511149
transform -1 0 5888 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1290_
timestamp 1644511149
transform 1 0 5152 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1291_
timestamp 1644511149
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1292_
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1293_
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1294_
timestamp 1644511149
transform -1 0 8372 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1295_
timestamp 1644511149
transform -1 0 8188 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1296_
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1297_
timestamp 1644511149
transform 1 0 26680 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1298_
timestamp 1644511149
transform -1 0 16284 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1299_
timestamp 1644511149
transform -1 0 17480 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1300_
timestamp 1644511149
transform -1 0 18492 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1644511149
transform -1 0 18308 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1644511149
transform -1 0 17572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1303_
timestamp 1644511149
transform -1 0 15916 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1304_
timestamp 1644511149
transform -1 0 15916 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1305_
timestamp 1644511149
transform -1 0 16008 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1306_
timestamp 1644511149
transform 1 0 22908 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1307_
timestamp 1644511149
transform 1 0 19688 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1308_
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1309_
timestamp 1644511149
transform 1 0 18216 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1310_
timestamp 1644511149
transform 1 0 18952 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1311_
timestamp 1644511149
transform -1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1312_
timestamp 1644511149
transform 1 0 3956 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _1313_
timestamp 1644511149
transform 1 0 15916 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1314_
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1315_
timestamp 1644511149
transform 1 0 27232 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1316_
timestamp 1644511149
transform 1 0 26772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1317_
timestamp 1644511149
transform -1 0 29072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1318_
timestamp 1644511149
transform 1 0 27600 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1319_
timestamp 1644511149
transform 1 0 27140 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1320_
timestamp 1644511149
transform -1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1321_
timestamp 1644511149
transform 1 0 25576 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1322_
timestamp 1644511149
transform 1 0 25852 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 1644511149
transform -1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1324_
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1325_
timestamp 1644511149
transform -1 0 24932 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1327_
timestamp 1644511149
transform -1 0 30820 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1328_
timestamp 1644511149
transform -1 0 31648 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1329_
timestamp 1644511149
transform -1 0 31280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1330_
timestamp 1644511149
transform -1 0 21344 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1331_
timestamp 1644511149
transform 1 0 21804 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1332_
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1333_
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1644511149
transform 1 0 25668 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1335_
timestamp 1644511149
transform -1 0 27232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1336_
timestamp 1644511149
transform -1 0 30452 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1337_
timestamp 1644511149
transform -1 0 30268 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1338_
timestamp 1644511149
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1339_
timestamp 1644511149
transform -1 0 36156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1340_
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1341_
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1342_
timestamp 1644511149
transform -1 0 30728 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1343_
timestamp 1644511149
transform 1 0 35144 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1344_
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1345_
timestamp 1644511149
transform -1 0 34132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1346_
timestamp 1644511149
transform -1 0 37260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1347_
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1348_
timestamp 1644511149
transform -1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1349_
timestamp 1644511149
transform -1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1350_
timestamp 1644511149
transform 1 0 35604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1351_
timestamp 1644511149
transform -1 0 36524 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1352_
timestamp 1644511149
transform 1 0 34960 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1353_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1354_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33304 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1355_
timestamp 1644511149
transform -1 0 35052 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1356_
timestamp 1644511149
transform 1 0 34040 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1357_
timestamp 1644511149
transform -1 0 33580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1358_
timestamp 1644511149
transform 1 0 33672 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1359_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34776 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1360_
timestamp 1644511149
transform 1 0 35236 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1361_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1644511149
transform 1 0 29992 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1364_
timestamp 1644511149
transform 1 0 32936 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1365_
timestamp 1644511149
transform 1 0 35236 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1366_
timestamp 1644511149
transform 1 0 34868 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1367_
timestamp 1644511149
transform 1 0 36248 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1368_
timestamp 1644511149
transform 1 0 31096 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1369_
timestamp 1644511149
transform 1 0 29716 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1370_
timestamp 1644511149
transform 1 0 30728 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1371_
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1372_
timestamp 1644511149
transform 1 0 31188 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1373_
timestamp 1644511149
transform 1 0 36064 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1644511149
transform 1 0 26496 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1375_
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1644511149
transform 1 0 35328 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1644511149
transform 1 0 35420 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1644511149
transform 1 0 35052 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1644511149
transform 1 0 35972 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1644511149
transform -1 0 33672 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1644511149
transform 1 0 13156 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1644511149
transform -1 0 11224 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1644511149
transform 1 0 2208 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1644511149
transform 1 0 2852 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1644511149
transform 1 0 5244 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1388_
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1644511149
transform -1 0 17848 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1390_
timestamp 1644511149
transform 1 0 19596 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1644511149
transform -1 0 29440 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1644511149
transform 1 0 27600 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1644511149
transform 1 0 23368 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1395_
timestamp 1644511149
transform 1 0 31096 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1396_
timestamp 1644511149
transform -1 0 22264 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1644511149
transform 1 0 27232 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1644511149
transform 1 0 29992 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1644511149
transform 1 0 33304 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1644511149
transform 1 0 34868 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1644511149
transform 1 0 36340 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1644511149
transform 1 0 34960 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1644511149
transform 1 0 34960 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1644511149
transform -1 0 33304 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1405__37 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1406__38
timestamp 1644511149
transform -1 0 6440 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1407__39
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1408__40
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1409__41
timestamp 1644511149
transform -1 0 2668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1410__42
timestamp 1644511149
transform -1 0 5428 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1411__43
timestamp 1644511149
transform -1 0 2944 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1412__44
timestamp 1644511149
transform 1 0 2392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1413__45
timestamp 1644511149
transform 1 0 2392 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1414__46
timestamp 1644511149
transform -1 0 5428 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1415__47
timestamp 1644511149
transform 1 0 4508 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1416__48
timestamp 1644511149
transform 1 0 2392 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1417__49
timestamp 1644511149
transform 1 0 2852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1418__50
timestamp 1644511149
transform -1 0 3128 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1419__51
timestamp 1644511149
transform 1 0 3036 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1420__52
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1421__53
timestamp 1644511149
transform -1 0 14352 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1422__54
timestamp 1644511149
transform -1 0 12696 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1423__55
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1424__56
timestamp 1644511149
transform -1 0 24656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1425__57
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1426__58
timestamp 1644511149
transform 1 0 25300 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1427__59
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1428__60
timestamp 1644511149
transform 1 0 23368 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1429__61
timestamp 1644511149
transform -1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1430__62
timestamp 1644511149
transform -1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1431__63
timestamp 1644511149
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1432__64
timestamp 1644511149
transform -1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1433__65
timestamp 1644511149
transform -1 0 13708 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1434__66
timestamp 1644511149
transform -1 0 14720 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1435__67
timestamp 1644511149
transform -1 0 11592 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1436__68
timestamp 1644511149
transform -1 0 12420 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1437__69
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1438__70
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1439__71
timestamp 1644511149
transform 1 0 10948 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1440__72
timestamp 1644511149
transform -1 0 9476 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1441__73
timestamp 1644511149
transform 1 0 8464 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1442__74
timestamp 1644511149
transform 1 0 5152 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1443__75
timestamp 1644511149
transform 1 0 6624 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1444__76
timestamp 1644511149
transform 1 0 5428 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1445__77
timestamp 1644511149
transform 1 0 15456 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1446__78
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1447__79
timestamp 1644511149
transform -1 0 24840 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1448__80
timestamp 1644511149
transform -1 0 23460 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1449__81
timestamp 1644511149
transform 1 0 25944 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1450__82
timestamp 1644511149
transform -1 0 23460 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1451__83
timestamp 1644511149
transform -1 0 23644 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1452__84
timestamp 1644511149
transform -1 0 23368 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1453__85
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1454__86
timestamp 1644511149
transform -1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1455__87
timestamp 1644511149
transform 1 0 5244 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1456__88
timestamp 1644511149
transform -1 0 9384 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1457__89
timestamp 1644511149
transform -1 0 9844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1458__90
timestamp 1644511149
transform -1 0 8188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1459__91
timestamp 1644511149
transform 1 0 19504 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1460__92
timestamp 1644511149
transform -1 0 15272 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1461__93
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1462__94
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1463__95
timestamp 1644511149
transform 1 0 14168 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1464__96
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1465__97
timestamp 1644511149
transform -1 0 7912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1466__98
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1467__99
timestamp 1644511149
transform 1 0 6900 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1468__100
timestamp 1644511149
transform 1 0 4508 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1469__101
timestamp 1644511149
transform -1 0 9384 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1470__102
timestamp 1644511149
transform 1 0 11776 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1471__103
timestamp 1644511149
transform -1 0 14352 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1472__104
timestamp 1644511149
transform -1 0 22080 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1473__105
timestamp 1644511149
transform -1 0 27232 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1474__106
timestamp 1644511149
transform -1 0 22080 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1475__107
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1476__108
timestamp 1644511149
transform 1 0 15548 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1477__109
timestamp 1644511149
transform -1 0 22632 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1478__110
timestamp 1644511149
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1479__111
timestamp 1644511149
transform 1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1480__112
timestamp 1644511149
transform -1 0 17848 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1481__113
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1482__114
timestamp 1644511149
transform 1 0 16100 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1483__115
timestamp 1644511149
transform -1 0 19964 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1484__116
timestamp 1644511149
transform 1 0 15088 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1485__117
timestamp 1644511149
transform 1 0 13248 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1486__118
timestamp 1644511149
transform -1 0 18768 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1487__119
timestamp 1644511149
transform 1 0 14076 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1488__120
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1489__121
timestamp 1644511149
transform 1 0 8464 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1490__122
timestamp 1644511149
transform 1 0 3036 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1491__123
timestamp 1644511149
transform 1 0 7452 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1492__124
timestamp 1644511149
transform -1 0 3404 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1493__125
timestamp 1644511149
transform 1 0 15824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1494__126
timestamp 1644511149
transform 1 0 17296 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1495__127
timestamp 1644511149
transform -1 0 20792 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1496__128
timestamp 1644511149
transform -1 0 22724 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1497__129
timestamp 1644511149
transform -1 0 25576 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1498__130
timestamp 1644511149
transform -1 0 20332 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1499__131
timestamp 1644511149
transform -1 0 21068 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1500__132
timestamp 1644511149
transform 1 0 20976 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1501__133
timestamp 1644511149
transform 1 0 37904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1502__134
timestamp 1644511149
transform 1 0 37904 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1503_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27692 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1504_
timestamp 1644511149
transform -1 0 30176 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1505_
timestamp 1644511149
transform -1 0 29900 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1506_
timestamp 1644511149
transform -1 0 29072 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1507_
timestamp 1644511149
transform -1 0 29348 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1508_
timestamp 1644511149
transform -1 0 31464 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1509_
timestamp 1644511149
transform -1 0 31188 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1510_
timestamp 1644511149
transform -1 0 24932 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1511_
timestamp 1644511149
transform 1 0 7360 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1512_
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1513_
timestamp 1644511149
transform -1 0 5428 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1514_
timestamp 1644511149
transform 1 0 5060 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1515_
timestamp 1644511149
transform 1 0 2392 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1516_
timestamp 1644511149
transform 1 0 5060 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1517_
timestamp 1644511149
transform 1 0 2668 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1518_
timestamp 1644511149
transform 1 0 2760 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1519_
timestamp 1644511149
transform 1 0 2576 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1520_
timestamp 1644511149
transform 1 0 5152 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1521_
timestamp 1644511149
transform 1 0 4784 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1522_
timestamp 1644511149
transform 1 0 2760 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1523_
timestamp 1644511149
transform 1 0 3496 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1524_
timestamp 1644511149
transform 1 0 2852 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1525_
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1526_
timestamp 1644511149
transform 1 0 2760 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1527_
timestamp 1644511149
transform 1 0 12788 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1528_
timestamp 1644511149
transform 1 0 12420 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1529_
timestamp 1644511149
transform -1 0 27508 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1530_
timestamp 1644511149
transform 1 0 24288 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1531_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1532_
timestamp 1644511149
transform -1 0 25576 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1533_
timestamp 1644511149
transform -1 0 26312 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1534_
timestamp 1644511149
transform -1 0 25300 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1535_
timestamp 1644511149
transform -1 0 27876 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1536_
timestamp 1644511149
transform -1 0 28980 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1537_
timestamp 1644511149
transform -1 0 29164 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1538_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1539_
timestamp 1644511149
transform -1 0 29072 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1540_
timestamp 1644511149
transform -1 0 30084 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1541_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1542_
timestamp 1644511149
transform -1 0 26312 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1543_
timestamp 1644511149
transform 1 0 22540 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1544_
timestamp 1644511149
transform 1 0 12512 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1545_
timestamp 1644511149
transform 1 0 3956 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1546_
timestamp 1644511149
transform 1 0 13340 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1547_
timestamp 1644511149
transform 1 0 12972 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1548_
timestamp 1644511149
transform 1 0 14444 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1549_
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1550_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1551_
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1552_
timestamp 1644511149
transform 1 0 9108 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1553_
timestamp 1644511149
transform 1 0 11408 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1554_
timestamp 1644511149
transform 1 0 9108 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1555_
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1556_
timestamp 1644511149
transform -1 0 5888 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1557_
timestamp 1644511149
transform 1 0 7268 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1558_
timestamp 1644511149
transform -1 0 6348 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1559_
timestamp 1644511149
transform 1 0 16100 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1560_
timestamp 1644511149
transform -1 0 19964 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1561_
timestamp 1644511149
transform 1 0 24472 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1562_
timestamp 1644511149
transform 1 0 23092 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1563_
timestamp 1644511149
transform 1 0 26680 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1564_
timestamp 1644511149
transform 1 0 22632 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1565_
timestamp 1644511149
transform 1 0 23276 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1566_
timestamp 1644511149
transform 1 0 23000 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1567_
timestamp 1644511149
transform 1 0 15088 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1568_
timestamp 1644511149
transform 1 0 15364 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1569_
timestamp 1644511149
transform 1 0 12420 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1570_
timestamp 1644511149
transform 1 0 9108 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1571_
timestamp 1644511149
transform 1 0 7636 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1572_
timestamp 1644511149
transform 1 0 10120 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1573_
timestamp 1644511149
transform 1 0 11960 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1574_
timestamp 1644511149
transform 1 0 10948 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1575_
timestamp 1644511149
transform 1 0 8372 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1576_
timestamp 1644511149
transform 1 0 8648 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1577_
timestamp 1644511149
transform -1 0 7084 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1578_
timestamp 1644511149
transform 1 0 9108 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1579_
timestamp 1644511149
transform 1 0 9108 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1580_
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1581_
timestamp 1644511149
transform 1 0 20148 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1582_
timestamp 1644511149
transform 1 0 14904 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1583_
timestamp 1644511149
transform -1 0 15916 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1584_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1585_
timestamp 1644511149
transform 1 0 14260 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1586_
timestamp 1644511149
transform -1 0 14076 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1587_
timestamp 1644511149
transform 1 0 7544 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1588_
timestamp 1644511149
transform 1 0 3404 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1589_
timestamp 1644511149
transform 1 0 7176 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1590_
timestamp 1644511149
transform -1 0 6348 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1591_
timestamp 1644511149
transform 1 0 9108 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1592_
timestamp 1644511149
transform 1 0 12420 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1593_
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1594_
timestamp 1644511149
transform 1 0 21712 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1595_
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1596_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1597_
timestamp 1644511149
transform 1 0 16744 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1598_
timestamp 1644511149
transform 1 0 16192 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1599_
timestamp 1644511149
transform -1 0 27232 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1600_
timestamp 1644511149
transform 1 0 27784 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1601_
timestamp 1644511149
transform 1 0 25208 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1602_
timestamp 1644511149
transform 1 0 21988 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1603_
timestamp 1644511149
transform -1 0 25852 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1604_
timestamp 1644511149
transform 1 0 19320 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1605_
timestamp 1644511149
transform 1 0 24932 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1606_
timestamp 1644511149
transform -1 0 26312 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1607_
timestamp 1644511149
transform 1 0 22264 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1608_
timestamp 1644511149
transform -1 0 14904 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1609_
timestamp 1644511149
transform 1 0 5244 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1610_
timestamp 1644511149
transform 1 0 17572 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1611_
timestamp 1644511149
transform 1 0 16744 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1612_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1613_
timestamp 1644511149
transform 1 0 19412 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1614_
timestamp 1644511149
transform -1 0 16928 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1615_
timestamp 1644511149
transform 1 0 13892 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1616_
timestamp 1644511149
transform 1 0 18492 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1617_
timestamp 1644511149
transform 1 0 14536 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1618_
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1619_
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1620_
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1621_
timestamp 1644511149
transform -1 0 9384 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1622_
timestamp 1644511149
transform 1 0 3128 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1623_
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1624_
timestamp 1644511149
transform 1 0 17480 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1625_
timestamp 1644511149
transform 1 0 19412 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1626_
timestamp 1644511149
transform 1 0 21896 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1627_
timestamp 1644511149
transform 1 0 24564 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1628_
timestamp 1644511149
transform 1 0 20056 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1629_
timestamp 1644511149
transform 1 0 20792 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1630_
timestamp 1644511149
transform 1 0 21620 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk
timestamp 1644511149
transform -1 0 22448 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 1644511149
transform 1 0 27324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_clk
timestamp 1644511149
transform -1 0 17020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_clk
timestamp 1644511149
transform 1 0 29256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_clk
timestamp 1644511149
transform 1 0 33672 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_clk
timestamp 1644511149
transform -1 0 30912 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform -1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform -1 0 1656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform -1 0 1656 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform -1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform -1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform -1 0 1656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform -1 0 1656 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform -1 0 1656 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform -1 0 1656 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform -1 0 1656 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform -1 0 1656 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1644511149
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1644511149
transform -1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 37904 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1644511149
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1644511149
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1644511149
transform 1 0 37812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1644511149
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1644511149
transform 1 0 37812 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1644511149
transform 1 0 37812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1644511149
transform 1 0 37812 0 1 36992
box -38 -48 406 592
<< labels >>
rlabel metal2 s 9954 39200 10010 40000 6 clk
port 0 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 peripheralBus_address[0]
port 1 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 peripheralBus_address[10]
port 2 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 peripheralBus_address[11]
port 3 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 peripheralBus_address[12]
port 4 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 peripheralBus_address[13]
port 5 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 peripheralBus_address[14]
port 6 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 peripheralBus_address[15]
port 7 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 peripheralBus_address[16]
port 8 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 peripheralBus_address[17]
port 9 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 peripheralBus_address[18]
port 10 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 peripheralBus_address[19]
port 11 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 peripheralBus_address[1]
port 12 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 peripheralBus_address[20]
port 13 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 peripheralBus_address[21]
port 14 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 peripheralBus_address[22]
port 15 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 peripheralBus_address[23]
port 16 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 peripheralBus_address[2]
port 17 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 peripheralBus_address[3]
port 18 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 peripheralBus_address[4]
port 19 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 peripheralBus_address[5]
port 20 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 peripheralBus_address[6]
port 21 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 peripheralBus_address[7]
port 22 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 peripheralBus_address[8]
port 23 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 peripheralBus_address[9]
port 24 nsew signal input
rlabel metal3 s 0 280 800 400 6 peripheralBus_busy
port 25 nsew signal tristate
rlabel metal3 s 0 2864 800 2984 6 peripheralBus_data[0]
port 26 nsew signal bidirectional
rlabel metal3 s 0 16464 800 16584 6 peripheralBus_data[10]
port 27 nsew signal bidirectional
rlabel metal3 s 0 17824 800 17944 6 peripheralBus_data[11]
port 28 nsew signal bidirectional
rlabel metal3 s 0 19184 800 19304 6 peripheralBus_data[12]
port 29 nsew signal bidirectional
rlabel metal3 s 0 20544 800 20664 6 peripheralBus_data[13]
port 30 nsew signal bidirectional
rlabel metal3 s 0 21904 800 22024 6 peripheralBus_data[14]
port 31 nsew signal bidirectional
rlabel metal3 s 0 23264 800 23384 6 peripheralBus_data[15]
port 32 nsew signal bidirectional
rlabel metal3 s 0 24624 800 24744 6 peripheralBus_data[16]
port 33 nsew signal bidirectional
rlabel metal3 s 0 25984 800 26104 6 peripheralBus_data[17]
port 34 nsew signal bidirectional
rlabel metal3 s 0 27344 800 27464 6 peripheralBus_data[18]
port 35 nsew signal bidirectional
rlabel metal3 s 0 28704 800 28824 6 peripheralBus_data[19]
port 36 nsew signal bidirectional
rlabel metal3 s 0 4224 800 4344 6 peripheralBus_data[1]
port 37 nsew signal bidirectional
rlabel metal3 s 0 30064 800 30184 6 peripheralBus_data[20]
port 38 nsew signal bidirectional
rlabel metal3 s 0 31424 800 31544 6 peripheralBus_data[21]
port 39 nsew signal bidirectional
rlabel metal3 s 0 32784 800 32904 6 peripheralBus_data[22]
port 40 nsew signal bidirectional
rlabel metal3 s 0 34144 800 34264 6 peripheralBus_data[23]
port 41 nsew signal bidirectional
rlabel metal3 s 0 34824 800 34944 6 peripheralBus_data[24]
port 42 nsew signal bidirectional
rlabel metal3 s 0 35504 800 35624 6 peripheralBus_data[25]
port 43 nsew signal bidirectional
rlabel metal3 s 0 36184 800 36304 6 peripheralBus_data[26]
port 44 nsew signal bidirectional
rlabel metal3 s 0 36864 800 36984 6 peripheralBus_data[27]
port 45 nsew signal bidirectional
rlabel metal3 s 0 37544 800 37664 6 peripheralBus_data[28]
port 46 nsew signal bidirectional
rlabel metal3 s 0 38224 800 38344 6 peripheralBus_data[29]
port 47 nsew signal bidirectional
rlabel metal3 s 0 5584 800 5704 6 peripheralBus_data[2]
port 48 nsew signal bidirectional
rlabel metal3 s 0 38904 800 39024 6 peripheralBus_data[30]
port 49 nsew signal bidirectional
rlabel metal3 s 0 39584 800 39704 6 peripheralBus_data[31]
port 50 nsew signal bidirectional
rlabel metal3 s 0 6944 800 7064 6 peripheralBus_data[3]
port 51 nsew signal bidirectional
rlabel metal3 s 0 8304 800 8424 6 peripheralBus_data[4]
port 52 nsew signal bidirectional
rlabel metal3 s 0 9664 800 9784 6 peripheralBus_data[5]
port 53 nsew signal bidirectional
rlabel metal3 s 0 11024 800 11144 6 peripheralBus_data[6]
port 54 nsew signal bidirectional
rlabel metal3 s 0 12384 800 12504 6 peripheralBus_data[7]
port 55 nsew signal bidirectional
rlabel metal3 s 0 13744 800 13864 6 peripheralBus_data[8]
port 56 nsew signal bidirectional
rlabel metal3 s 0 15104 800 15224 6 peripheralBus_data[9]
port 57 nsew signal bidirectional
rlabel metal3 s 0 824 800 944 6 peripheralBus_oe
port 58 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 peripheralBus_we
port 59 nsew signal input
rlabel metal2 s 29918 39200 29974 40000 6 rst
port 60 nsew signal input
rlabel metal3 s 39200 1912 40000 2032 6 spi_clk[0]
port 61 nsew signal tristate
rlabel metal3 s 39200 21904 40000 22024 6 spi_clk[1]
port 62 nsew signal tristate
rlabel metal3 s 39200 5856 40000 5976 6 spi_cs[0]
port 63 nsew signal tristate
rlabel metal3 s 39200 25848 40000 25968 6 spi_cs[1]
port 64 nsew signal tristate
rlabel metal3 s 39200 9800 40000 9920 6 spi_en[0]
port 65 nsew signal tristate
rlabel metal3 s 39200 29792 40000 29912 6 spi_en[1]
port 66 nsew signal tristate
rlabel metal3 s 39200 13880 40000 14000 6 spi_miso[0]
port 67 nsew signal input
rlabel metal3 s 39200 33872 40000 33992 6 spi_miso[1]
port 68 nsew signal input
rlabel metal3 s 39200 17824 40000 17944 6 spi_mosi[0]
port 69 nsew signal tristate
rlabel metal3 s 39200 37816 40000 37936 6 spi_mosi[1]
port 70 nsew signal tristate
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 71 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 71 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 72 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
