magic
tech sky130A
magscale 1 2
timestamp 1650726245
<< viali >>
rect 5273 11305 5307 11339
rect 5457 11305 5491 11339
rect 7389 11305 7423 11339
rect 3985 11237 4019 11271
rect 4629 11237 4663 11271
rect 7573 11237 7607 11271
rect 3065 11101 3099 11135
rect 3249 11101 3283 11135
rect 3801 11101 3835 11135
rect 4445 11101 4479 11135
rect 4629 11101 4663 11135
rect 6561 11101 6595 11135
rect 6745 11101 6779 11135
rect 8033 11101 8067 11135
rect 8217 11101 8251 11135
rect 3157 11033 3191 11067
rect 5089 11033 5123 11067
rect 7205 11033 7239 11067
rect 7421 11033 7455 11067
rect 8125 11033 8159 11067
rect 1409 10965 1443 10999
rect 5289 10965 5323 10999
rect 6377 10965 6411 10999
rect 6653 10761 6687 10795
rect 7757 10761 7791 10795
rect 5089 10693 5123 10727
rect 6745 10693 6779 10727
rect 2697 10625 2731 10659
rect 3341 10625 3375 10659
rect 4261 10625 4295 10659
rect 4709 10625 4743 10659
rect 4813 10625 4847 10659
rect 4951 10625 4985 10659
rect 5197 10625 5231 10659
rect 6561 10625 6595 10659
rect 7389 10625 7423 10659
rect 7573 10625 7607 10659
rect 8217 10625 8251 10659
rect 8401 10625 8435 10659
rect 8493 10625 8527 10659
rect 9137 10625 9171 10659
rect 1409 10557 1443 10591
rect 1685 10557 1719 10591
rect 3985 10557 4019 10591
rect 3525 10489 3559 10523
rect 6929 10489 6963 10523
rect 2881 10421 2915 10455
rect 4077 10421 4111 10455
rect 4169 10421 4203 10455
rect 4721 10421 4755 10455
rect 6377 10421 6411 10455
rect 8217 10421 8251 10455
rect 8953 10421 8987 10455
rect 7665 10217 7699 10251
rect 8309 10217 8343 10251
rect 4261 10149 4295 10183
rect 6653 10149 6687 10183
rect 4445 10081 4479 10115
rect 4538 10081 4572 10115
rect 4629 10081 4663 10115
rect 7297 10081 7331 10115
rect 7389 10081 7423 10115
rect 8125 10081 8159 10115
rect 1777 10013 1811 10047
rect 1961 10013 1995 10047
rect 2421 10013 2455 10047
rect 3065 10013 3099 10047
rect 4721 10013 4755 10047
rect 5273 10013 5307 10047
rect 7205 10013 7239 10047
rect 7481 10013 7515 10047
rect 8401 10013 8435 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 9597 10013 9631 10047
rect 1869 9945 1903 9979
rect 5540 9945 5574 9979
rect 8125 9945 8159 9979
rect 2605 9877 2639 9911
rect 3157 9877 3191 9911
rect 9045 9877 9079 9911
rect 9689 9877 9723 9911
rect 6377 9673 6411 9707
rect 3893 9605 3927 9639
rect 7512 9605 7546 9639
rect 9229 9605 9263 9639
rect 1501 9537 1535 9571
rect 2145 9537 2179 9571
rect 2329 9537 2363 9571
rect 3065 9537 3099 9571
rect 3709 9537 3743 9571
rect 3985 9537 4019 9571
rect 4445 9537 4479 9571
rect 4701 9537 4735 9571
rect 8401 9537 8435 9571
rect 8585 9537 8619 9571
rect 9413 9537 9447 9571
rect 2789 9469 2823 9503
rect 3525 9469 3559 9503
rect 7757 9469 7791 9503
rect 8493 9469 8527 9503
rect 8677 9469 8711 9503
rect 2881 9401 2915 9435
rect 9597 9401 9631 9435
rect 1685 9333 1719 9367
rect 2329 9333 2363 9367
rect 2973 9333 3007 9367
rect 5825 9333 5859 9367
rect 8217 9333 8251 9367
rect 2237 9129 2271 9163
rect 3026 9129 3060 9163
rect 3249 9129 3283 9163
rect 3985 9129 4019 9163
rect 9965 9129 9999 9163
rect 6837 9061 6871 9095
rect 4997 8993 5031 9027
rect 8953 8993 8987 9027
rect 1961 8925 1995 8959
rect 2053 8925 2087 8959
rect 2697 8925 2731 8959
rect 4261 8925 4295 8959
rect 8217 8925 8251 8959
rect 9045 8925 9079 8959
rect 9137 8925 9171 8959
rect 9413 8925 9447 8959
rect 9505 8925 9539 8959
rect 10149 8925 10183 8959
rect 2237 8857 2271 8891
rect 4353 8857 4387 8891
rect 4537 8857 4571 8891
rect 5264 8857 5298 8891
rect 7972 8857 8006 8891
rect 9229 8857 9263 8891
rect 3065 8789 3099 8823
rect 4169 8789 4203 8823
rect 6377 8789 6411 8823
rect 5273 8585 5307 8619
rect 6377 8585 6411 8619
rect 1777 8517 1811 8551
rect 1961 8517 1995 8551
rect 7512 8517 7546 8551
rect 2145 8449 2179 8483
rect 2881 8449 2915 8483
rect 3893 8449 3927 8483
rect 4149 8449 4183 8483
rect 7757 8449 7791 8483
rect 9341 8449 9375 8483
rect 2605 8381 2639 8415
rect 9597 8381 9631 8415
rect 5733 8313 5767 8347
rect 8217 8313 8251 8347
rect 1961 8041 1995 8075
rect 4077 8041 4111 8075
rect 1593 7905 1627 7939
rect 1777 7905 1811 7939
rect 3249 7905 3283 7939
rect 7297 7905 7331 7939
rect 8953 7905 8987 7939
rect 9229 7905 9263 7939
rect 1501 7837 1535 7871
rect 1685 7837 1719 7871
rect 2973 7837 3007 7871
rect 5457 7837 5491 7871
rect 7030 7837 7064 7871
rect 7941 7837 7975 7871
rect 5190 7769 5224 7803
rect 8309 7769 8343 7803
rect 5917 7701 5951 7735
rect 7757 7701 7791 7735
rect 8033 7701 8067 7735
rect 8125 7701 8159 7735
rect 1501 7497 1535 7531
rect 5365 7497 5399 7531
rect 8217 7497 8251 7531
rect 1685 7429 1719 7463
rect 3258 7429 3292 7463
rect 9330 7429 9364 7463
rect 1409 7361 1443 7395
rect 3525 7361 3559 7395
rect 3985 7361 4019 7395
rect 4241 7361 4275 7395
rect 6644 7361 6678 7395
rect 9597 7361 9631 7395
rect 6377 7293 6411 7327
rect 1685 7225 1719 7259
rect 2145 7157 2179 7191
rect 7757 7157 7791 7191
rect 4721 6953 4755 6987
rect 3801 6885 3835 6919
rect 8401 6885 8435 6919
rect 1869 6749 1903 6783
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 8953 6749 8987 6783
rect 9965 6749 9999 6783
rect 10149 6749 10183 6783
rect 2136 6681 2170 6715
rect 4813 6681 4847 6715
rect 5825 6681 5859 6715
rect 8219 6681 8253 6715
rect 9229 6681 9263 6715
rect 3249 6613 3283 6647
rect 7113 6613 7147 6647
rect 9137 6613 9171 6647
rect 9321 6613 9355 6647
rect 9505 6613 9539 6647
rect 10057 6613 10091 6647
rect 1961 6341 1995 6375
rect 8576 6341 8610 6375
rect 3718 6273 3752 6307
rect 3985 6273 4019 6307
rect 5569 6273 5603 6307
rect 5825 6273 5859 6307
rect 6469 6273 6503 6307
rect 6725 6273 6759 6307
rect 8309 6273 8343 6307
rect 1593 6137 1627 6171
rect 1961 6069 1995 6103
rect 2145 6069 2179 6103
rect 2605 6069 2639 6103
rect 4445 6069 4479 6103
rect 7849 6069 7883 6103
rect 9689 6069 9723 6103
rect 3065 5865 3099 5899
rect 8953 5865 8987 5899
rect 10057 5865 10091 5899
rect 5825 5729 5859 5763
rect 7757 5729 7791 5763
rect 9229 5729 9263 5763
rect 9413 5729 9447 5763
rect 2053 5661 2087 5695
rect 2145 5661 2179 5695
rect 2697 5661 2731 5695
rect 5558 5661 5592 5695
rect 9137 5661 9171 5695
rect 9321 5661 9355 5695
rect 9965 5661 9999 5695
rect 10149 5661 10183 5695
rect 7512 5593 7546 5627
rect 1869 5525 1903 5559
rect 3065 5525 3099 5559
rect 3249 5525 3283 5559
rect 4445 5525 4479 5559
rect 6377 5525 6411 5559
rect 2529 5321 2563 5355
rect 2697 5321 2731 5355
rect 5549 5321 5583 5355
rect 8493 5321 8527 5355
rect 8769 5321 8803 5355
rect 2329 5253 2363 5287
rect 1593 5185 1627 5219
rect 3248 5185 3282 5219
rect 3433 5185 3467 5219
rect 4169 5185 4203 5219
rect 4436 5185 4470 5219
rect 6377 5185 6411 5219
rect 6644 5185 6678 5219
rect 8217 5185 8251 5219
rect 8401 5185 8435 5219
rect 8585 5185 8619 5219
rect 9413 5185 9447 5219
rect 9597 5185 9631 5219
rect 1869 5117 1903 5151
rect 3341 5117 3375 5151
rect 3525 5117 3559 5151
rect 1777 5049 1811 5083
rect 9229 5049 9263 5083
rect 1685 4981 1719 5015
rect 2513 4981 2547 5015
rect 3709 4981 3743 5015
rect 7757 4981 7791 5015
rect 3157 4777 3191 4811
rect 5641 4777 5675 4811
rect 8217 4777 8251 4811
rect 9229 4777 9263 4811
rect 1777 4709 1811 4743
rect 2329 4709 2363 4743
rect 9781 4709 9815 4743
rect 2513 4641 2547 4675
rect 2973 4641 3007 4675
rect 4261 4641 4295 4675
rect 6377 4641 6411 4675
rect 9045 4641 9079 4675
rect 1593 4573 1627 4607
rect 2237 4573 2271 4607
rect 3249 4573 3283 4607
rect 8401 4573 8435 4607
rect 9321 4573 9355 4607
rect 10057 4573 10091 4607
rect 4528 4505 4562 4539
rect 6644 4505 6678 4539
rect 9781 4505 9815 4539
rect 2513 4437 2547 4471
rect 2973 4437 3007 4471
rect 7757 4437 7791 4471
rect 9045 4437 9079 4471
rect 9965 4437 9999 4471
rect 2815 4233 2849 4267
rect 3985 4233 4019 4267
rect 8953 4233 8987 4267
rect 2605 4165 2639 4199
rect 3801 4165 3835 4199
rect 1961 4097 1995 4131
rect 2145 4097 2179 4131
rect 4445 4097 4479 4131
rect 4712 4097 4746 4131
rect 8125 4097 8159 4131
rect 8769 4097 8803 4131
rect 9045 4097 9079 4131
rect 9873 4097 9907 4131
rect 2053 4029 2087 4063
rect 7205 4029 7239 4063
rect 7481 4029 7515 4063
rect 7941 4029 7975 4063
rect 8309 4029 8343 4063
rect 3433 3961 3467 3995
rect 5825 3961 5859 3995
rect 10057 3961 10091 3995
rect 2789 3893 2823 3927
rect 2973 3893 3007 3927
rect 3801 3893 3835 3927
rect 8769 3893 8803 3927
rect 2145 3689 2179 3723
rect 2881 3689 2915 3723
rect 6469 3689 6503 3723
rect 7113 3689 7147 3723
rect 7297 3689 7331 3723
rect 9137 3689 9171 3723
rect 5641 3621 5675 3655
rect 8309 3621 8343 3655
rect 4261 3553 4295 3587
rect 6101 3553 6135 3587
rect 2145 3485 2179 3519
rect 2329 3485 2363 3519
rect 2973 3485 3007 3519
rect 4445 3485 4479 3519
rect 5365 3485 5399 3519
rect 5457 3485 5491 3519
rect 7205 3485 7239 3519
rect 7481 3485 7515 3519
rect 8033 3485 8067 3519
rect 8309 3485 8343 3519
rect 8953 3485 8987 3519
rect 9137 3485 9171 3519
rect 4629 3417 4663 3451
rect 5273 3417 5307 3451
rect 7573 3417 7607 3451
rect 5089 3349 5123 3383
rect 6469 3349 6503 3383
rect 6653 3349 6687 3383
rect 8125 3349 8159 3383
rect 3249 3145 3283 3179
rect 4737 3145 4771 3179
rect 7665 3145 7699 3179
rect 8585 3145 8619 3179
rect 4537 3077 4571 3111
rect 3065 3009 3099 3043
rect 3801 3009 3835 3043
rect 3985 3009 4019 3043
rect 4077 3009 4111 3043
rect 5365 3009 5399 3043
rect 5549 3009 5583 3043
rect 5641 3009 5675 3043
rect 7205 3009 7239 3043
rect 7941 3009 7975 3043
rect 8401 3009 8435 3043
rect 6929 2941 6963 2975
rect 7665 2941 7699 2975
rect 3801 2873 3835 2907
rect 4905 2873 4939 2907
rect 7113 2873 7147 2907
rect 7849 2873 7883 2907
rect 4721 2805 4755 2839
rect 7021 2805 7055 2839
rect 4261 2601 4295 2635
rect 4353 2601 4387 2635
rect 5089 2601 5123 2635
rect 5181 2601 5215 2635
rect 6561 2601 6595 2635
rect 7113 2601 7147 2635
rect 7941 2601 7975 2635
rect 6469 2533 6503 2567
rect 4169 2465 4203 2499
rect 4997 2465 5031 2499
rect 6377 2465 6411 2499
rect 2421 2397 2455 2431
rect 2605 2397 2639 2431
rect 3065 2397 3099 2431
rect 3249 2397 3283 2431
rect 4445 2397 4479 2431
rect 5273 2397 5307 2431
rect 6653 2397 6687 2431
rect 7297 2397 7331 2431
rect 7757 2397 7791 2431
rect 3157 2329 3191 2363
rect 2513 2261 2547 2295
<< metal1 >>
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 10134 11540 10140 11552
rect 5500 11512 10140 11540
rect 5500 11500 5506 11512
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 1104 11450 10856 11472
rect 1104 11398 2582 11450
rect 2634 11398 2646 11450
rect 2698 11398 2710 11450
rect 2762 11398 2774 11450
rect 2826 11398 2838 11450
rect 2890 11398 5846 11450
rect 5898 11398 5910 11450
rect 5962 11398 5974 11450
rect 6026 11398 6038 11450
rect 6090 11398 6102 11450
rect 6154 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 9238 11450
rect 9290 11398 9302 11450
rect 9354 11398 9366 11450
rect 9418 11398 10856 11450
rect 1104 11376 10856 11398
rect 4798 11296 4804 11348
rect 4856 11336 4862 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 4856 11308 5273 11336
rect 4856 11296 4862 11308
rect 5261 11305 5273 11308
rect 5307 11305 5319 11339
rect 5442 11336 5448 11348
rect 5403 11308 5448 11336
rect 5261 11299 5319 11305
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 7377 11339 7435 11345
rect 7377 11305 7389 11339
rect 7423 11336 7435 11339
rect 8110 11336 8116 11348
rect 7423 11308 8116 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 3970 11268 3976 11280
rect 3931 11240 3976 11268
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 4617 11271 4675 11277
rect 4617 11237 4629 11271
rect 4663 11268 4675 11271
rect 5166 11268 5172 11280
rect 4663 11240 5172 11268
rect 4663 11237 4675 11240
rect 4617 11231 4675 11237
rect 5166 11228 5172 11240
rect 5224 11228 5230 11280
rect 7561 11271 7619 11277
rect 7561 11237 7573 11271
rect 7607 11268 7619 11271
rect 9122 11268 9128 11280
rect 7607 11240 9128 11268
rect 7607 11237 7619 11240
rect 7561 11231 7619 11237
rect 9122 11228 9128 11240
rect 9180 11228 9186 11280
rect 4522 11200 4528 11212
rect 3068 11172 4528 11200
rect 3068 11141 3096 11172
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 6822 11200 6828 11212
rect 6564 11172 6828 11200
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 3234 11132 3240 11144
rect 3195 11104 3240 11132
rect 3053 11095 3111 11101
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 3786 11132 3792 11144
rect 3747 11104 3792 11132
rect 3786 11092 3792 11104
rect 3844 11092 3850 11144
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 4212 11104 4445 11132
rect 4212 11092 4218 11104
rect 4433 11101 4445 11104
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 4982 11132 4988 11144
rect 4663 11104 4988 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5350 11092 5356 11144
rect 5408 11092 5414 11144
rect 6564 11141 6592 11172
rect 6822 11160 6828 11172
rect 6880 11200 6886 11212
rect 8754 11200 8760 11212
rect 6880 11172 8760 11200
rect 6880 11160 6886 11172
rect 6549 11135 6607 11141
rect 6549 11101 6561 11135
rect 6595 11101 6607 11135
rect 6730 11132 6736 11144
rect 6691 11104 6736 11132
rect 6549 11095 6607 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 8036 11141 8064 11172
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8202 11132 8208 11144
rect 8163 11104 8208 11132
rect 8021 11095 8079 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 3142 11064 3148 11076
rect 3103 11036 3148 11064
rect 3142 11024 3148 11036
rect 3200 11024 3206 11076
rect 5077 11067 5135 11073
rect 5077 11033 5089 11067
rect 5123 11064 5135 11067
rect 5368 11064 5396 11092
rect 7193 11067 7251 11073
rect 7193 11064 7205 11067
rect 5123 11036 7205 11064
rect 5123 11033 5135 11036
rect 5077 11027 5135 11033
rect 7193 11033 7205 11036
rect 7239 11033 7251 11067
rect 7193 11027 7251 11033
rect 7409 11067 7467 11073
rect 7409 11033 7421 11067
rect 7455 11064 7467 11067
rect 8113 11067 8171 11073
rect 8113 11064 8125 11067
rect 7455 11036 8125 11064
rect 7455 11033 7467 11036
rect 7409 11027 7467 11033
rect 8113 11033 8125 11036
rect 8159 11064 8171 11067
rect 8478 11064 8484 11076
rect 8159 11036 8484 11064
rect 8159 11033 8171 11036
rect 8113 11027 8171 11033
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 1394 10996 1400 11008
rect 1355 10968 1400 10996
rect 1394 10956 1400 10968
rect 1452 10956 1458 11008
rect 4890 10956 4896 11008
rect 4948 10996 4954 11008
rect 5258 10996 5264 11008
rect 5316 11005 5322 11008
rect 5316 10999 5335 11005
rect 4948 10968 5264 10996
rect 4948 10956 4954 10968
rect 5258 10956 5264 10968
rect 5323 10965 5335 10999
rect 5316 10959 5335 10965
rect 6365 10999 6423 11005
rect 6365 10965 6377 10999
rect 6411 10996 6423 10999
rect 6546 10996 6552 11008
rect 6411 10968 6552 10996
rect 6411 10965 6423 10968
rect 6365 10959 6423 10965
rect 5316 10956 5322 10959
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 1104 10906 10856 10928
rect 1104 10854 4214 10906
rect 4266 10854 4278 10906
rect 4330 10854 4342 10906
rect 4394 10854 4406 10906
rect 4458 10854 4470 10906
rect 4522 10854 7478 10906
rect 7530 10854 7542 10906
rect 7594 10854 7606 10906
rect 7658 10854 7670 10906
rect 7722 10854 7734 10906
rect 7786 10854 10856 10906
rect 1104 10832 10856 10854
rect 6641 10795 6699 10801
rect 6641 10792 6653 10795
rect 2746 10764 6653 10792
rect 1762 10684 1768 10736
rect 1820 10724 1826 10736
rect 2746 10724 2774 10764
rect 6641 10761 6653 10764
rect 6687 10792 6699 10795
rect 7745 10795 7803 10801
rect 6687 10764 7696 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 1820 10696 2774 10724
rect 1820 10684 1826 10696
rect 5074 10684 5080 10736
rect 5132 10724 5138 10736
rect 5132 10696 5177 10724
rect 5132 10684 5138 10696
rect 6362 10684 6368 10736
rect 6420 10724 6426 10736
rect 6733 10727 6791 10733
rect 6733 10724 6745 10727
rect 6420 10696 6745 10724
rect 6420 10684 6426 10696
rect 6733 10693 6745 10696
rect 6779 10724 6791 10727
rect 7668 10724 7696 10764
rect 7745 10761 7757 10795
rect 7791 10792 7803 10795
rect 8202 10792 8208 10804
rect 7791 10764 8208 10792
rect 7791 10761 7803 10764
rect 7745 10755 7803 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8662 10724 8668 10736
rect 6779 10696 7420 10724
rect 6779 10693 6791 10696
rect 6733 10687 6791 10693
rect 2498 10656 2504 10668
rect 1688 10628 2504 10656
rect 1688 10600 1716 10628
rect 2498 10616 2504 10628
rect 2556 10656 2562 10668
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2556 10628 2697 10656
rect 2556 10616 2562 10628
rect 2685 10625 2697 10628
rect 2731 10656 2743 10659
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 2731 10628 3341 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 4430 10656 4436 10668
rect 4295 10628 4436 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 4697 10659 4755 10665
rect 4580 10654 4660 10656
rect 4697 10654 4709 10659
rect 4580 10628 4709 10654
rect 4580 10616 4586 10628
rect 4632 10626 4709 10628
rect 4697 10625 4709 10626
rect 4743 10625 4755 10659
rect 4697 10619 4755 10625
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 1670 10588 1676 10600
rect 1631 10560 1676 10588
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 3970 10588 3976 10600
rect 3528 10560 3976 10588
rect 3326 10480 3332 10532
rect 3384 10520 3390 10532
rect 3528 10529 3556 10560
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 4816 10588 4844 10619
rect 4890 10616 4896 10668
rect 4948 10665 4954 10668
rect 4948 10659 4997 10665
rect 4948 10625 4951 10659
rect 4985 10625 4997 10659
rect 4948 10619 4997 10625
rect 5185 10659 5243 10665
rect 5185 10625 5197 10659
rect 5231 10656 5243 10659
rect 6546 10656 6552 10668
rect 5231 10628 5304 10656
rect 6507 10628 6552 10656
rect 5231 10625 5243 10628
rect 5185 10619 5243 10625
rect 4948 10616 4954 10619
rect 4816 10560 4936 10588
rect 4908 10532 4936 10560
rect 5276 10532 5304 10628
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 7392 10665 7420 10696
rect 7668 10696 8668 10724
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7668 10656 7696 10696
rect 8662 10684 8668 10696
rect 8720 10684 8726 10736
rect 7607 10628 7696 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 8018 10616 8024 10668
rect 8076 10656 8082 10668
rect 8205 10659 8263 10665
rect 8205 10656 8217 10659
rect 8076 10628 8217 10656
rect 8076 10616 8082 10628
rect 8205 10625 8217 10628
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 9122 10656 9128 10668
rect 9083 10628 9128 10656
rect 8481 10619 8539 10625
rect 7098 10548 7104 10600
rect 7156 10588 7162 10600
rect 8404 10588 8432 10619
rect 7156 10560 8432 10588
rect 7156 10548 7162 10560
rect 3513 10523 3571 10529
rect 3513 10520 3525 10523
rect 3384 10492 3525 10520
rect 3384 10480 3390 10492
rect 3513 10489 3525 10492
rect 3559 10489 3571 10523
rect 3513 10483 3571 10489
rect 4890 10480 4896 10532
rect 4948 10480 4954 10532
rect 5258 10480 5264 10532
rect 5316 10480 5322 10532
rect 6914 10520 6920 10532
rect 6875 10492 6920 10520
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 8496 10520 8524 10619
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 7484 10492 8524 10520
rect 7484 10464 7512 10492
rect 2869 10455 2927 10461
rect 2869 10421 2881 10455
rect 2915 10452 2927 10455
rect 3050 10452 3056 10464
rect 2915 10424 3056 10452
rect 2915 10421 2927 10424
rect 2869 10415 2927 10421
rect 3050 10412 3056 10424
rect 3108 10412 3114 10464
rect 4062 10452 4068 10464
rect 4023 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 4614 10452 4620 10464
rect 4203 10424 4620 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 4709 10455 4767 10461
rect 4709 10421 4721 10455
rect 4755 10452 4767 10455
rect 5534 10452 5540 10464
rect 4755 10424 5540 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 6328 10424 6377 10452
rect 6328 10412 6334 10424
rect 6365 10421 6377 10424
rect 6411 10452 6423 10455
rect 7466 10452 7472 10464
rect 6411 10424 7472 10452
rect 6411 10421 6423 10424
rect 6365 10415 6423 10421
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 8205 10455 8263 10461
rect 8205 10421 8217 10455
rect 8251 10452 8263 10455
rect 8294 10452 8300 10464
rect 8251 10424 8300 10452
rect 8251 10421 8263 10424
rect 8205 10415 8263 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8938 10452 8944 10464
rect 8899 10424 8944 10452
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 1104 10362 10856 10384
rect 1104 10310 2582 10362
rect 2634 10310 2646 10362
rect 2698 10310 2710 10362
rect 2762 10310 2774 10362
rect 2826 10310 2838 10362
rect 2890 10310 5846 10362
rect 5898 10310 5910 10362
rect 5962 10310 5974 10362
rect 6026 10310 6038 10362
rect 6090 10310 6102 10362
rect 6154 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 9238 10362
rect 9290 10310 9302 10362
rect 9354 10310 9366 10362
rect 9418 10310 10856 10362
rect 1104 10288 10856 10310
rect 3510 10208 3516 10260
rect 3568 10248 3574 10260
rect 5442 10248 5448 10260
rect 3568 10220 5448 10248
rect 3568 10208 3574 10220
rect 2314 10140 2320 10192
rect 2372 10180 2378 10192
rect 4249 10183 4307 10189
rect 4249 10180 4261 10183
rect 2372 10152 4261 10180
rect 2372 10140 2378 10152
rect 4249 10149 4261 10152
rect 4295 10149 4307 10183
rect 4249 10143 4307 10149
rect 4062 10112 4068 10124
rect 1964 10084 4068 10112
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 1964 10053 1992 10084
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 4540 10121 4568 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 7653 10251 7711 10257
rect 7653 10217 7665 10251
rect 7699 10248 7711 10251
rect 7926 10248 7932 10260
rect 7699 10220 7932 10248
rect 7699 10217 7711 10220
rect 7653 10211 7711 10217
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8297 10251 8355 10257
rect 8297 10217 8309 10251
rect 8343 10248 8355 10251
rect 8662 10248 8668 10260
rect 8343 10220 8668 10248
rect 8343 10217 8355 10220
rect 8297 10211 8355 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 6641 10183 6699 10189
rect 6641 10149 6653 10183
rect 6687 10180 6699 10183
rect 6730 10180 6736 10192
rect 6687 10152 6736 10180
rect 6687 10149 6699 10152
rect 6641 10143 6699 10149
rect 6730 10140 6736 10152
rect 6788 10180 6794 10192
rect 6788 10152 9628 10180
rect 6788 10140 6794 10152
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 4212 10084 4445 10112
rect 4212 10072 4218 10084
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 4526 10115 4584 10121
rect 4526 10081 4538 10115
rect 4572 10081 4584 10115
rect 4526 10075 4584 10081
rect 4617 10115 4675 10121
rect 4617 10081 4629 10115
rect 4663 10112 4675 10115
rect 4890 10112 4896 10124
rect 4663 10084 4896 10112
rect 4663 10081 4675 10084
rect 4617 10075 4675 10081
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 7285 10115 7343 10121
rect 7285 10112 7297 10115
rect 7156 10084 7297 10112
rect 7156 10072 7162 10084
rect 7285 10081 7297 10084
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 7834 10112 7840 10124
rect 7423 10084 7840 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 8113 10115 8171 10121
rect 8113 10081 8125 10115
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10013 2007 10047
rect 2406 10044 2412 10056
rect 2367 10016 2412 10044
rect 1949 10007 2007 10013
rect 2406 10004 2412 10016
rect 2464 10004 2470 10056
rect 2498 10004 2504 10056
rect 2556 10044 2562 10056
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 2556 10016 3065 10044
rect 2556 10004 2562 10016
rect 3053 10013 3065 10016
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 3418 10004 3424 10056
rect 3476 10044 3482 10056
rect 4172 10044 4200 10072
rect 4709 10047 4767 10053
rect 4709 10044 4721 10047
rect 3476 10016 4200 10044
rect 4264 10016 4721 10044
rect 3476 10004 3482 10016
rect 1857 9979 1915 9985
rect 1857 9945 1869 9979
rect 1903 9976 1915 9979
rect 3602 9976 3608 9988
rect 1903 9948 3608 9976
rect 1903 9945 1915 9948
rect 1857 9939 1915 9945
rect 3602 9936 3608 9948
rect 3660 9936 3666 9988
rect 2590 9908 2596 9920
rect 2551 9880 2596 9908
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 3145 9911 3203 9917
rect 3145 9877 3157 9911
rect 3191 9908 3203 9911
rect 3234 9908 3240 9920
rect 3191 9880 3240 9908
rect 3191 9877 3203 9880
rect 3145 9871 3203 9877
rect 3234 9868 3240 9880
rect 3292 9908 3298 9920
rect 4264 9908 4292 10016
rect 4709 10013 4721 10016
rect 4755 10013 4767 10047
rect 5258 10044 5264 10056
rect 5219 10016 5264 10044
rect 4709 10007 4767 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 7064 10016 7205 10044
rect 7064 10004 7070 10016
rect 7193 10013 7205 10016
rect 7239 10013 7251 10047
rect 7466 10044 7472 10056
rect 7427 10016 7472 10044
rect 7193 10007 7251 10013
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 7558 10004 7564 10056
rect 7616 10044 7622 10056
rect 8128 10044 8156 10075
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 8260 10084 9168 10112
rect 8260 10072 8266 10084
rect 7616 10016 8156 10044
rect 8389 10047 8447 10053
rect 7616 10004 7622 10016
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 8570 10044 8576 10056
rect 8435 10016 8576 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 9140 10053 9168 10084
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9214 10044 9220 10056
rect 9171 10016 9220 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 4430 9936 4436 9988
rect 4488 9936 4494 9988
rect 5528 9979 5586 9985
rect 5528 9945 5540 9979
rect 5574 9976 5586 9979
rect 8113 9979 8171 9985
rect 5574 9948 7696 9976
rect 5574 9945 5586 9948
rect 5528 9939 5586 9945
rect 3292 9880 4292 9908
rect 4448 9908 4476 9936
rect 6178 9908 6184 9920
rect 4448 9880 6184 9908
rect 3292 9868 3298 9880
rect 6178 9868 6184 9880
rect 6236 9868 6242 9920
rect 7668 9908 7696 9948
rect 8113 9945 8125 9979
rect 8159 9976 8171 9979
rect 8956 9976 8984 10007
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9600 10053 9628 10152
rect 9585 10047 9643 10053
rect 9585 10013 9597 10047
rect 9631 10013 9643 10047
rect 9585 10007 9643 10013
rect 8159 9948 8984 9976
rect 8159 9945 8171 9948
rect 8113 9939 8171 9945
rect 8386 9908 8392 9920
rect 7668 9880 8392 9908
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 9030 9908 9036 9920
rect 8991 9880 9036 9908
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9582 9868 9588 9920
rect 9640 9908 9646 9920
rect 9677 9911 9735 9917
rect 9677 9908 9689 9911
rect 9640 9880 9689 9908
rect 9640 9868 9646 9880
rect 9677 9877 9689 9880
rect 9723 9877 9735 9911
rect 9677 9871 9735 9877
rect 1104 9818 10856 9840
rect 1104 9766 4214 9818
rect 4266 9766 4278 9818
rect 4330 9766 4342 9818
rect 4394 9766 4406 9818
rect 4458 9766 4470 9818
rect 4522 9766 7478 9818
rect 7530 9766 7542 9818
rect 7594 9766 7606 9818
rect 7658 9766 7670 9818
rect 7722 9766 7734 9818
rect 7786 9766 10856 9818
rect 1104 9744 10856 9766
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 5074 9704 5080 9716
rect 2648 9676 5080 9704
rect 2648 9664 2654 9676
rect 3326 9636 3332 9648
rect 2792 9608 3332 9636
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9568 1547 9571
rect 1670 9568 1676 9580
rect 1535 9540 1676 9568
rect 1535 9537 1547 9540
rect 1489 9531 1547 9537
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2314 9568 2320 9580
rect 2275 9540 2320 9568
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 2792 9509 2820 9608
rect 3326 9596 3332 9608
rect 3384 9596 3390 9648
rect 3510 9636 3516 9648
rect 3436 9608 3516 9636
rect 2958 9528 2964 9580
rect 3016 9568 3022 9580
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 3016 9540 3065 9568
rect 3016 9528 3022 9540
rect 3053 9537 3065 9540
rect 3099 9568 3111 9571
rect 3436 9568 3464 9608
rect 3510 9596 3516 9608
rect 3568 9596 3574 9648
rect 3896 9645 3924 9676
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 6365 9707 6423 9713
rect 6365 9673 6377 9707
rect 6411 9673 6423 9707
rect 6365 9667 6423 9673
rect 3881 9639 3939 9645
rect 3881 9605 3893 9639
rect 3927 9636 3939 9639
rect 4982 9636 4988 9648
rect 3927 9608 3961 9636
rect 4448 9608 4988 9636
rect 3927 9605 3939 9608
rect 3881 9599 3939 9605
rect 3694 9568 3700 9580
rect 3099 9540 3464 9568
rect 3655 9540 3700 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 3970 9568 3976 9580
rect 3883 9540 3976 9568
rect 3970 9528 3976 9540
rect 4028 9568 4034 9580
rect 4154 9568 4160 9580
rect 4028 9540 4160 9568
rect 4028 9528 4034 9540
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4448 9577 4476 9608
rect 4982 9596 4988 9608
rect 5040 9636 5046 9648
rect 5258 9636 5264 9648
rect 5040 9608 5264 9636
rect 5040 9596 5046 9608
rect 5258 9596 5264 9608
rect 5316 9596 5322 9648
rect 6380 9636 6408 9667
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 8570 9704 8576 9716
rect 6512 9676 8576 9704
rect 6512 9664 6518 9676
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 8662 9664 8668 9716
rect 8720 9664 8726 9716
rect 7098 9636 7104 9648
rect 6380 9608 7104 9636
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 7500 9639 7558 9645
rect 7500 9605 7512 9639
rect 7546 9636 7558 9639
rect 8294 9636 8300 9648
rect 7546 9608 8300 9636
rect 7546 9605 7558 9608
rect 7500 9599 7558 9605
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 8680 9636 8708 9664
rect 8496 9608 8708 9636
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4522 9528 4528 9580
rect 4580 9568 4586 9580
rect 4689 9571 4747 9577
rect 4689 9568 4701 9571
rect 4580 9540 4701 9568
rect 4580 9528 4586 9540
rect 4689 9537 4701 9540
rect 4735 9537 4747 9571
rect 4689 9531 4747 9537
rect 6546 9528 6552 9580
rect 6604 9568 6610 9580
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 6604 9540 8401 9568
rect 6604 9528 6610 9540
rect 8312 9512 8340 9540
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9469 2835 9503
rect 3418 9492 3424 9512
rect 2777 9463 2835 9469
rect 3344 9464 3424 9492
rect 1946 9392 1952 9444
rect 2004 9432 2010 9444
rect 2869 9435 2927 9441
rect 2869 9432 2881 9435
rect 2004 9404 2881 9432
rect 2004 9392 2010 9404
rect 2869 9401 2881 9404
rect 2915 9401 2927 9435
rect 2869 9395 2927 9401
rect 1670 9364 1676 9376
rect 1631 9336 1676 9364
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 2314 9364 2320 9376
rect 2275 9336 2320 9364
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 2961 9367 3019 9373
rect 2961 9333 2973 9367
rect 3007 9364 3019 9367
rect 3344 9364 3372 9464
rect 3418 9460 3424 9464
rect 3476 9460 3482 9512
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9500 3571 9503
rect 7742 9500 7748 9512
rect 3559 9472 3648 9500
rect 7703 9472 7748 9500
rect 3559 9469 3571 9472
rect 3513 9463 3571 9469
rect 3620 9376 3648 9472
rect 7742 9460 7748 9472
rect 7800 9460 7806 9512
rect 8294 9460 8300 9512
rect 8352 9460 8358 9512
rect 8496 9509 8524 9608
rect 8846 9596 8852 9648
rect 8904 9636 8910 9648
rect 9214 9636 9220 9648
rect 8904 9608 9220 9636
rect 8904 9596 8910 9608
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 8570 9528 8576 9580
rect 8628 9568 8634 9580
rect 8628 9540 8673 9568
rect 8628 9528 8634 9540
rect 8754 9528 8760 9580
rect 8812 9568 8818 9580
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 8812 9540 9413 9568
rect 8812 9528 8818 9540
rect 9401 9537 9413 9540
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 8481 9503 8539 9509
rect 8481 9469 8493 9503
rect 8527 9469 8539 9503
rect 8481 9463 8539 9469
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 9122 9500 9128 9512
rect 8711 9472 9128 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 9585 9435 9643 9441
rect 9585 9432 9597 9435
rect 9548 9404 9597 9432
rect 9548 9392 9554 9404
rect 9585 9401 9597 9404
rect 9631 9401 9643 9435
rect 9585 9395 9643 9401
rect 3418 9364 3424 9376
rect 3007 9336 3424 9364
rect 3007 9333 3019 9336
rect 2961 9327 3019 9333
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3602 9324 3608 9376
rect 3660 9324 3666 9376
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9364 5871 9367
rect 6178 9364 6184 9376
rect 5859 9336 6184 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6454 9324 6460 9376
rect 6512 9364 6518 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 6512 9336 8217 9364
rect 6512 9324 6518 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8205 9327 8263 9333
rect 1104 9274 10856 9296
rect 1104 9222 2582 9274
rect 2634 9222 2646 9274
rect 2698 9222 2710 9274
rect 2762 9222 2774 9274
rect 2826 9222 2838 9274
rect 2890 9222 5846 9274
rect 5898 9222 5910 9274
rect 5962 9222 5974 9274
rect 6026 9222 6038 9274
rect 6090 9222 6102 9274
rect 6154 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 9238 9274
rect 9290 9222 9302 9274
rect 9354 9222 9366 9274
rect 9418 9222 10856 9274
rect 1104 9200 10856 9222
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 2225 9163 2283 9169
rect 2225 9160 2237 9163
rect 2188 9132 2237 9160
rect 2188 9120 2194 9132
rect 2225 9129 2237 9132
rect 2271 9129 2283 9163
rect 3014 9163 3072 9169
rect 3014 9160 3026 9163
rect 2225 9123 2283 9129
rect 2884 9132 3026 9160
rect 2774 9024 2780 9036
rect 2056 8996 2780 9024
rect 2056 8968 2084 8996
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 1394 8916 1400 8968
rect 1452 8956 1458 8968
rect 1949 8959 2007 8965
rect 1949 8956 1961 8959
rect 1452 8928 1961 8956
rect 1452 8916 1458 8928
rect 1949 8925 1961 8928
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2038 8916 2044 8968
rect 2096 8956 2102 8968
rect 2096 8928 2189 8956
rect 2096 8916 2102 8928
rect 2498 8916 2504 8968
rect 2556 8956 2562 8968
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2556 8928 2697 8956
rect 2556 8916 2562 8928
rect 2685 8925 2697 8928
rect 2731 8925 2743 8959
rect 2884 8956 2912 9132
rect 3014 9129 3026 9132
rect 3060 9129 3072 9163
rect 3014 9123 3072 9129
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3786 9160 3792 9172
rect 3283 9132 3792 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 4246 9160 4252 9172
rect 4019 9132 4252 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 4246 9120 4252 9132
rect 4304 9160 4310 9172
rect 5626 9160 5632 9172
rect 4304 9132 5632 9160
rect 4304 9120 4310 9132
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 8662 9120 8668 9172
rect 8720 9160 8726 9172
rect 9953 9163 10011 9169
rect 9953 9160 9965 9163
rect 8720 9132 9965 9160
rect 8720 9120 8726 9132
rect 9953 9129 9965 9132
rect 9999 9129 10011 9163
rect 9953 9123 10011 9129
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 4614 9092 4620 9104
rect 3384 9064 4620 9092
rect 3384 9052 3390 9064
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 6822 9092 6828 9104
rect 6783 9064 6828 9092
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 8846 9052 8852 9104
rect 8904 9092 8910 9104
rect 8904 9064 9168 9092
rect 8904 9052 8910 9064
rect 4982 9024 4988 9036
rect 4943 8996 4988 9024
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 8941 9027 8999 9033
rect 8941 9024 8953 9027
rect 8444 8996 8953 9024
rect 8444 8984 8450 8996
rect 8941 8993 8953 8996
rect 8987 8993 8999 9027
rect 8941 8987 8999 8993
rect 2958 8956 2964 8968
rect 2884 8928 2964 8956
rect 2685 8919 2743 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 5074 8956 5080 8968
rect 4295 8928 5080 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 8110 8956 8116 8968
rect 7852 8928 8116 8956
rect 1578 8848 1584 8900
rect 1636 8888 1642 8900
rect 2225 8891 2283 8897
rect 2225 8888 2237 8891
rect 1636 8860 2237 8888
rect 1636 8848 1642 8860
rect 2225 8857 2237 8860
rect 2271 8888 2283 8891
rect 4341 8891 4399 8897
rect 4341 8888 4353 8891
rect 2271 8860 4353 8888
rect 2271 8857 2283 8860
rect 2225 8851 2283 8857
rect 4341 8857 4353 8860
rect 4387 8857 4399 8891
rect 4341 8851 4399 8857
rect 4525 8891 4583 8897
rect 4525 8857 4537 8891
rect 4571 8888 4583 8891
rect 4614 8888 4620 8900
rect 4571 8860 4620 8888
rect 4571 8857 4583 8860
rect 4525 8851 4583 8857
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 3053 8823 3111 8829
rect 3053 8820 3065 8823
rect 1728 8792 3065 8820
rect 1728 8780 1734 8792
rect 3053 8789 3065 8792
rect 3099 8820 3111 8823
rect 3510 8820 3516 8832
rect 3099 8792 3516 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 4157 8823 4215 8829
rect 4157 8820 4169 8823
rect 4120 8792 4169 8820
rect 4120 8780 4126 8792
rect 4157 8789 4169 8792
rect 4203 8789 4215 8823
rect 4356 8820 4384 8851
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 5252 8891 5310 8897
rect 5252 8857 5264 8891
rect 5298 8888 5310 8891
rect 5350 8888 5356 8900
rect 5298 8860 5356 8888
rect 5298 8857 5310 8860
rect 5252 8851 5310 8857
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 7742 8848 7748 8900
rect 7800 8888 7806 8900
rect 7852 8888 7880 8928
rect 8110 8916 8116 8928
rect 8168 8956 8174 8968
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 8168 8928 8217 8956
rect 8168 8916 8174 8928
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 9140 8965 9168 9064
rect 9582 9024 9588 9036
rect 9416 8996 9588 9024
rect 9416 8965 9444 8996
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 8352 8928 9045 8956
rect 8352 8916 8358 8928
rect 9033 8925 9045 8928
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 10134 8956 10140 8968
rect 9548 8928 9593 8956
rect 10095 8928 10140 8956
rect 9548 8916 9554 8928
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 7800 8860 7880 8888
rect 7960 8891 8018 8897
rect 7800 8848 7806 8860
rect 7960 8857 7972 8891
rect 8006 8888 8018 8891
rect 8938 8888 8944 8900
rect 8006 8860 8944 8888
rect 8006 8857 8018 8860
rect 7960 8851 8018 8857
rect 8938 8848 8944 8860
rect 8996 8848 9002 8900
rect 9217 8891 9275 8897
rect 9217 8857 9229 8891
rect 9263 8857 9275 8891
rect 9217 8851 9275 8857
rect 4890 8820 4896 8832
rect 4356 8792 4896 8820
rect 4157 8783 4215 8789
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 6365 8823 6423 8829
rect 6365 8789 6377 8823
rect 6411 8820 6423 8823
rect 7282 8820 7288 8832
rect 6411 8792 7288 8820
rect 6411 8789 6423 8792
rect 6365 8783 6423 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 9232 8820 9260 8851
rect 8536 8792 9260 8820
rect 8536 8780 8542 8792
rect 1104 8730 10856 8752
rect 1104 8678 4214 8730
rect 4266 8678 4278 8730
rect 4330 8678 4342 8730
rect 4394 8678 4406 8730
rect 4458 8678 4470 8730
rect 4522 8678 7478 8730
rect 7530 8678 7542 8730
rect 7594 8678 7606 8730
rect 7658 8678 7670 8730
rect 7722 8678 7734 8730
rect 7786 8678 10856 8730
rect 1104 8656 10856 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 3418 8616 3424 8628
rect 1452 8588 3424 8616
rect 1452 8576 1458 8588
rect 1762 8548 1768 8560
rect 1723 8520 1768 8548
rect 1762 8508 1768 8520
rect 1820 8508 1826 8560
rect 1949 8551 2007 8557
rect 1949 8517 1961 8551
rect 1995 8548 2007 8551
rect 1995 8520 2820 8548
rect 1995 8517 2007 8520
rect 1949 8511 2007 8517
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 2314 8440 2320 8492
rect 2372 8480 2378 8492
rect 2372 8452 2728 8480
rect 2372 8440 2378 8452
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8381 2651 8415
rect 2593 8375 2651 8381
rect 1854 8236 1860 8288
rect 1912 8276 1918 8288
rect 2608 8276 2636 8375
rect 2700 8344 2728 8452
rect 2792 8412 2820 8520
rect 2884 8489 2912 8588
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 3510 8576 3516 8628
rect 3568 8616 3574 8628
rect 4706 8616 4712 8628
rect 3568 8588 4712 8616
rect 3568 8576 3574 8588
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 4948 8588 5273 8616
rect 4948 8576 4954 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 6362 8616 6368 8628
rect 6323 8588 6368 8616
rect 5261 8579 5319 8585
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 9030 8616 9036 8628
rect 7668 8588 9036 8616
rect 4982 8548 4988 8560
rect 3896 8520 4988 8548
rect 3896 8489 3924 8520
rect 4982 8508 4988 8520
rect 5040 8508 5046 8560
rect 7500 8551 7558 8557
rect 7500 8517 7512 8551
rect 7546 8548 7558 8551
rect 7668 8548 7696 8588
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 8110 8548 8116 8560
rect 7546 8520 7696 8548
rect 7760 8520 8116 8548
rect 7546 8517 7558 8520
rect 7500 8511 7558 8517
rect 7760 8492 7788 8520
rect 8110 8508 8116 8520
rect 8168 8548 8174 8560
rect 8168 8520 9628 8548
rect 8168 8508 8174 8520
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 4137 8483 4195 8489
rect 4137 8480 4149 8483
rect 3881 8443 3939 8449
rect 3988 8452 4149 8480
rect 3786 8412 3792 8424
rect 2792 8384 3792 8412
rect 3786 8372 3792 8384
rect 3844 8372 3850 8424
rect 3988 8412 4016 8452
rect 4137 8449 4149 8452
rect 4183 8449 4195 8483
rect 4137 8443 4195 8449
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 4890 8480 4896 8492
rect 4764 8452 4896 8480
rect 4764 8440 4770 8452
rect 4890 8440 4896 8452
rect 4948 8480 4954 8492
rect 5258 8480 5264 8492
rect 4948 8452 5264 8480
rect 4948 8440 4954 8452
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 7742 8480 7748 8492
rect 7655 8452 7748 8480
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 9329 8483 9387 8489
rect 9329 8449 9341 8483
rect 9375 8480 9387 8483
rect 9490 8480 9496 8492
rect 9375 8452 9496 8480
rect 9375 8449 9387 8452
rect 9329 8443 9387 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9600 8424 9628 8520
rect 9582 8412 9588 8424
rect 3896 8384 4016 8412
rect 9543 8384 9588 8412
rect 3896 8344 3924 8384
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 5718 8344 5724 8356
rect 2700 8316 3924 8344
rect 5679 8316 5724 8344
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 7834 8304 7840 8356
rect 7892 8344 7898 8356
rect 8205 8347 8263 8353
rect 8205 8344 8217 8347
rect 7892 8316 8217 8344
rect 7892 8304 7898 8316
rect 8205 8313 8217 8316
rect 8251 8344 8263 8347
rect 8386 8344 8392 8356
rect 8251 8316 8392 8344
rect 8251 8313 8263 8316
rect 8205 8307 8263 8313
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 4154 8276 4160 8288
rect 1912 8248 4160 8276
rect 1912 8236 1918 8248
rect 4154 8236 4160 8248
rect 4212 8236 4218 8288
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 8478 8276 8484 8288
rect 5500 8248 8484 8276
rect 5500 8236 5506 8248
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 1104 8186 10856 8208
rect 1104 8134 2582 8186
rect 2634 8134 2646 8186
rect 2698 8134 2710 8186
rect 2762 8134 2774 8186
rect 2826 8134 2838 8186
rect 2890 8134 5846 8186
rect 5898 8134 5910 8186
rect 5962 8134 5974 8186
rect 6026 8134 6038 8186
rect 6090 8134 6102 8186
rect 6154 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 9238 8186
rect 9290 8134 9302 8186
rect 9354 8134 9366 8186
rect 9418 8134 10856 8186
rect 1104 8112 10856 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2958 8072 2964 8084
rect 1995 8044 2964 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8072 4123 8075
rect 4154 8072 4160 8084
rect 4111 8044 4160 8072
rect 4111 8041 4123 8044
rect 4065 8035 4123 8041
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 5132 8044 8432 8072
rect 5132 8032 5138 8044
rect 1578 7936 1584 7948
rect 1539 7908 1584 7936
rect 1578 7896 1584 7908
rect 1636 7896 1642 7948
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7936 1823 7939
rect 1854 7936 1860 7948
rect 1811 7908 1860 7936
rect 1811 7905 1823 7908
rect 1765 7899 1823 7905
rect 1854 7896 1860 7908
rect 1912 7896 1918 7948
rect 3234 7936 3240 7948
rect 3195 7908 3240 7936
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 7742 7936 7748 7948
rect 7331 7908 7748 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 8404 7936 8432 8044
rect 8478 7964 8484 8016
rect 8536 8004 8542 8016
rect 8536 7976 9260 8004
rect 8536 7964 8542 7976
rect 9232 7945 9260 7976
rect 8941 7939 8999 7945
rect 8941 7936 8953 7939
rect 8404 7908 8953 7936
rect 8941 7905 8953 7908
rect 8987 7905 8999 7939
rect 8941 7899 8999 7905
rect 9217 7939 9275 7945
rect 9217 7905 9229 7939
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7837 1547 7871
rect 1489 7831 1547 7837
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 2038 7868 2044 7880
rect 1719 7840 2044 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 1504 7800 1532 7831
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3326 7868 3332 7880
rect 3007 7840 3332 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 5445 7871 5503 7877
rect 5445 7868 5457 7871
rect 5000 7840 5457 7868
rect 5000 7812 5028 7840
rect 5445 7837 5457 7840
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 7006 7828 7012 7880
rect 7064 7877 7070 7880
rect 7064 7868 7076 7877
rect 7929 7871 7987 7877
rect 7064 7840 7109 7868
rect 7064 7831 7076 7840
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 9030 7868 9036 7880
rect 7975 7840 9036 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 7064 7828 7070 7831
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 4614 7800 4620 7812
rect 1504 7772 4620 7800
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 4982 7760 4988 7812
rect 5040 7760 5046 7812
rect 5166 7760 5172 7812
rect 5224 7809 5230 7812
rect 5224 7800 5236 7809
rect 8297 7803 8355 7809
rect 5224 7772 5269 7800
rect 5224 7763 5236 7772
rect 8297 7769 8309 7803
rect 8343 7800 8355 7803
rect 8846 7800 8852 7812
rect 8343 7772 8852 7800
rect 8343 7769 8355 7772
rect 8297 7763 8355 7769
rect 5224 7760 5230 7763
rect 8846 7760 8852 7772
rect 8904 7760 8910 7812
rect 4632 7732 4660 7760
rect 5905 7735 5963 7741
rect 5905 7732 5917 7735
rect 4632 7704 5917 7732
rect 5905 7701 5917 7704
rect 5951 7701 5963 7735
rect 5905 7695 5963 7701
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 7745 7735 7803 7741
rect 7745 7732 7757 7735
rect 7248 7704 7757 7732
rect 7248 7692 7254 7704
rect 7745 7701 7757 7704
rect 7791 7701 7803 7735
rect 7745 7695 7803 7701
rect 7834 7692 7840 7744
rect 7892 7732 7898 7744
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 7892 7704 8033 7732
rect 7892 7692 7898 7704
rect 8021 7701 8033 7704
rect 8067 7701 8079 7735
rect 8021 7695 8079 7701
rect 8113 7735 8171 7741
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 8478 7732 8484 7744
rect 8159 7704 8484 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 1104 7642 10856 7664
rect 1104 7590 4214 7642
rect 4266 7590 4278 7642
rect 4330 7590 4342 7642
rect 4394 7590 4406 7642
rect 4458 7590 4470 7642
rect 4522 7590 7478 7642
rect 7530 7590 7542 7642
rect 7594 7590 7606 7642
rect 7658 7590 7670 7642
rect 7722 7590 7734 7642
rect 7786 7590 10856 7642
rect 1104 7568 10856 7590
rect 1489 7531 1547 7537
rect 1489 7497 1501 7531
rect 1535 7528 1547 7531
rect 2038 7528 2044 7540
rect 1535 7500 2044 7528
rect 1535 7497 1547 7500
rect 1489 7491 1547 7497
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 5074 7488 5080 7540
rect 5132 7528 5138 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 5132 7500 5365 7528
rect 5132 7488 5138 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 8202 7528 8208 7540
rect 8163 7500 8208 7528
rect 5353 7491 5411 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7460 1731 7463
rect 1946 7460 1952 7472
rect 1719 7432 1952 7460
rect 1719 7429 1731 7432
rect 1673 7423 1731 7429
rect 1946 7420 1952 7432
rect 2004 7420 2010 7472
rect 3142 7420 3148 7472
rect 3200 7460 3206 7472
rect 3246 7463 3304 7469
rect 3246 7460 3258 7463
rect 3200 7432 3258 7460
rect 3200 7420 3206 7432
rect 3246 7429 3258 7432
rect 3292 7429 3304 7463
rect 4982 7460 4988 7472
rect 3246 7423 3304 7429
rect 3988 7432 4988 7460
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 3988 7401 4016 7432
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 7834 7420 7840 7472
rect 7892 7460 7898 7472
rect 8294 7460 8300 7472
rect 7892 7432 8300 7460
rect 7892 7420 7898 7432
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 8662 7420 8668 7472
rect 8720 7460 8726 7472
rect 9318 7463 9376 7469
rect 9318 7460 9330 7463
rect 8720 7432 9330 7460
rect 8720 7420 8726 7432
rect 9318 7429 9330 7432
rect 9364 7429 9376 7463
rect 9318 7423 9376 7429
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7392 3571 7395
rect 3973 7395 4031 7401
rect 3973 7392 3985 7395
rect 3559 7364 3985 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 3973 7361 3985 7364
rect 4019 7361 4031 7395
rect 4229 7395 4287 7401
rect 4229 7392 4241 7395
rect 3973 7355 4031 7361
rect 4080 7364 4241 7392
rect 4080 7324 4108 7364
rect 4229 7361 4241 7364
rect 4275 7361 4287 7395
rect 4229 7355 4287 7361
rect 6632 7395 6690 7401
rect 6632 7361 6644 7395
rect 6678 7392 6690 7395
rect 7374 7392 7380 7404
rect 6678 7364 7380 7392
rect 6678 7361 6690 7364
rect 6632 7355 6690 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 9582 7392 9588 7404
rect 9543 7364 9588 7392
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 6362 7324 6368 7336
rect 3528 7296 4108 7324
rect 6323 7296 6368 7324
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 1719 7228 2636 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 1762 7148 1768 7200
rect 1820 7188 1826 7200
rect 2133 7191 2191 7197
rect 2133 7188 2145 7191
rect 1820 7160 2145 7188
rect 1820 7148 1826 7160
rect 2133 7157 2145 7160
rect 2179 7157 2191 7191
rect 2608 7188 2636 7228
rect 3528 7188 3556 7296
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 2608 7160 3556 7188
rect 7745 7191 7803 7197
rect 2133 7151 2191 7157
rect 7745 7157 7757 7191
rect 7791 7188 7803 7191
rect 8938 7188 8944 7200
rect 7791 7160 8944 7188
rect 7791 7157 7803 7160
rect 7745 7151 7803 7157
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 1104 7098 10856 7120
rect 1104 7046 2582 7098
rect 2634 7046 2646 7098
rect 2698 7046 2710 7098
rect 2762 7046 2774 7098
rect 2826 7046 2838 7098
rect 2890 7046 5846 7098
rect 5898 7046 5910 7098
rect 5962 7046 5974 7098
rect 6026 7046 6038 7098
rect 6090 7046 6102 7098
rect 6154 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 9238 7098
rect 9290 7046 9302 7098
rect 9354 7046 9366 7098
rect 9418 7046 10856 7098
rect 1104 7024 10856 7046
rect 1854 6944 1860 6996
rect 1912 6984 1918 6996
rect 4062 6984 4068 6996
rect 1912 6956 4068 6984
rect 1912 6944 1918 6956
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 4709 6987 4767 6993
rect 4709 6953 4721 6987
rect 4755 6984 4767 6987
rect 4982 6984 4988 6996
rect 4755 6956 4988 6984
rect 4755 6953 4767 6956
rect 4709 6947 4767 6953
rect 3789 6919 3847 6925
rect 3789 6885 3801 6919
rect 3835 6916 3847 6919
rect 4154 6916 4160 6928
rect 3835 6888 4160 6916
rect 3835 6885 3847 6888
rect 3789 6879 3847 6885
rect 4154 6876 4160 6888
rect 4212 6876 4218 6928
rect 4724 6848 4752 6947
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 8389 6919 8447 6925
rect 8389 6916 8401 6919
rect 8352 6888 8401 6916
rect 8352 6876 8358 6888
rect 8389 6885 8401 6888
rect 8435 6916 8447 6919
rect 9582 6916 9588 6928
rect 8435 6888 9588 6916
rect 8435 6885 8447 6888
rect 8389 6879 8447 6885
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 3896 6820 4752 6848
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 3896 6780 3924 6820
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 5684 6820 9076 6848
rect 5684 6808 5690 6820
rect 1903 6752 3924 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4157 6783 4215 6789
rect 4028 6752 4073 6780
rect 4028 6740 4034 6752
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 2124 6715 2182 6721
rect 2124 6681 2136 6715
rect 2170 6712 2182 6715
rect 2222 6712 2228 6724
rect 2170 6684 2228 6712
rect 2170 6681 2182 6684
rect 2124 6675 2182 6681
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 3878 6672 3884 6724
rect 3936 6712 3942 6724
rect 4172 6712 4200 6743
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 7892 6752 8953 6780
rect 7892 6740 7898 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 3936 6684 4200 6712
rect 4801 6715 4859 6721
rect 3936 6672 3942 6684
rect 4801 6681 4813 6715
rect 4847 6681 4859 6715
rect 4801 6675 4859 6681
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 3200 6616 3249 6644
rect 3200 6604 3206 6616
rect 3237 6613 3249 6616
rect 3283 6613 3295 6647
rect 3237 6607 3295 6613
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 3694 6644 3700 6656
rect 3384 6616 3700 6644
rect 3384 6604 3390 6616
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 4816 6644 4844 6675
rect 5718 6672 5724 6724
rect 5776 6712 5782 6724
rect 5813 6715 5871 6721
rect 5813 6712 5825 6715
rect 5776 6684 5825 6712
rect 5776 6672 5782 6684
rect 5813 6681 5825 6684
rect 5859 6681 5871 6715
rect 5813 6675 5871 6681
rect 8207 6715 8265 6721
rect 8207 6681 8219 6715
rect 8253 6681 8265 6715
rect 9048 6712 9076 6820
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 9364 6820 10180 6848
rect 9364 6808 9370 6820
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 10152 6789 10180 6820
rect 9953 6783 10011 6789
rect 9953 6780 9965 6783
rect 9456 6752 9965 6780
rect 9456 6740 9462 6752
rect 9953 6749 9965 6752
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 9217 6715 9275 6721
rect 9217 6712 9229 6715
rect 9048 6684 9229 6712
rect 8207 6675 8265 6681
rect 9217 6681 9229 6684
rect 9263 6681 9275 6715
rect 9217 6675 9275 6681
rect 7101 6647 7159 6653
rect 7101 6644 7113 6647
rect 4816 6616 7113 6644
rect 7101 6613 7113 6616
rect 7147 6644 7159 6647
rect 8220 6644 8248 6675
rect 9122 6644 9128 6656
rect 7147 6616 8248 6644
rect 9083 6616 9128 6644
rect 7147 6613 7159 6616
rect 7101 6607 7159 6613
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9306 6644 9312 6656
rect 9267 6616 9312 6644
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 9490 6644 9496 6656
rect 9451 6616 9496 6644
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 9582 6604 9588 6656
rect 9640 6644 9646 6656
rect 10045 6647 10103 6653
rect 10045 6644 10057 6647
rect 9640 6616 10057 6644
rect 9640 6604 9646 6616
rect 10045 6613 10057 6616
rect 10091 6613 10103 6647
rect 10045 6607 10103 6613
rect 1104 6554 10856 6576
rect 1104 6502 4214 6554
rect 4266 6502 4278 6554
rect 4330 6502 4342 6554
rect 4394 6502 4406 6554
rect 4458 6502 4470 6554
rect 4522 6502 7478 6554
rect 7530 6502 7542 6554
rect 7594 6502 7606 6554
rect 7658 6502 7670 6554
rect 7722 6502 7734 6554
rect 7786 6502 10856 6554
rect 1104 6480 10856 6502
rect 2314 6400 2320 6452
rect 2372 6440 2378 6452
rect 10134 6440 10140 6452
rect 2372 6412 10140 6440
rect 2372 6400 2378 6412
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 1949 6375 2007 6381
rect 1949 6341 1961 6375
rect 1995 6372 2007 6375
rect 2958 6372 2964 6384
rect 1995 6344 2964 6372
rect 1995 6341 2007 6344
rect 1949 6335 2007 6341
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 6362 6332 6368 6384
rect 6420 6372 6426 6384
rect 8564 6375 8622 6381
rect 6420 6344 8340 6372
rect 6420 6332 6426 6344
rect 3694 6304 3700 6316
rect 3752 6313 3758 6316
rect 3664 6276 3700 6304
rect 3694 6264 3700 6276
rect 3752 6267 3764 6313
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6304 4031 6307
rect 4982 6304 4988 6316
rect 4019 6276 4988 6304
rect 4019 6273 4031 6276
rect 3973 6267 4031 6273
rect 3752 6264 3758 6267
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 6472 6313 6500 6344
rect 8312 6316 8340 6344
rect 8564 6341 8576 6375
rect 8610 6372 8622 6375
rect 9582 6372 9588 6384
rect 8610 6344 9588 6372
rect 8610 6341 8622 6344
rect 8564 6335 8622 6341
rect 9582 6332 9588 6344
rect 9640 6332 9646 6384
rect 5557 6307 5615 6313
rect 5557 6273 5569 6307
rect 5603 6304 5615 6307
rect 5813 6307 5871 6313
rect 5603 6276 5764 6304
rect 5603 6273 5615 6276
rect 5557 6267 5615 6273
rect 5736 6236 5764 6276
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 6457 6307 6515 6313
rect 6457 6304 6469 6307
rect 5859 6276 6469 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6457 6273 6469 6276
rect 6503 6273 6515 6307
rect 6457 6267 6515 6273
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 6713 6307 6771 6313
rect 6713 6304 6725 6307
rect 6604 6276 6725 6304
rect 6604 6264 6610 6276
rect 6713 6273 6725 6276
rect 6759 6273 6771 6307
rect 8294 6304 8300 6316
rect 8255 6276 8300 6304
rect 6713 6267 6771 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 5736 6208 5856 6236
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 1670 6168 1676 6180
rect 1627 6140 1676 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 1670 6128 1676 6140
rect 1728 6128 1734 6180
rect 1946 6100 1952 6112
rect 1907 6072 1952 6100
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2130 6100 2136 6112
rect 2091 6072 2136 6100
rect 2130 6060 2136 6072
rect 2188 6060 2194 6112
rect 2406 6060 2412 6112
rect 2464 6100 2470 6112
rect 2593 6103 2651 6109
rect 2593 6100 2605 6103
rect 2464 6072 2605 6100
rect 2464 6060 2470 6072
rect 2593 6069 2605 6072
rect 2639 6069 2651 6103
rect 2593 6063 2651 6069
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4433 6103 4491 6109
rect 4433 6100 4445 6103
rect 4028 6072 4445 6100
rect 4028 6060 4034 6072
rect 4433 6069 4445 6072
rect 4479 6100 4491 6103
rect 4706 6100 4712 6112
rect 4479 6072 4712 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 5828 6100 5856 6208
rect 7392 6140 7972 6168
rect 7392 6100 7420 6140
rect 7834 6100 7840 6112
rect 5828 6072 7420 6100
rect 7795 6072 7840 6100
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 7944 6100 7972 6140
rect 8570 6100 8576 6112
rect 7944 6072 8576 6100
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 9858 6100 9864 6112
rect 9723 6072 9864 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 1104 6010 10856 6032
rect 1104 5958 2582 6010
rect 2634 5958 2646 6010
rect 2698 5958 2710 6010
rect 2762 5958 2774 6010
rect 2826 5958 2838 6010
rect 2890 5958 5846 6010
rect 5898 5958 5910 6010
rect 5962 5958 5974 6010
rect 6026 5958 6038 6010
rect 6090 5958 6102 6010
rect 6154 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 9238 6010
rect 9290 5958 9302 6010
rect 9354 5958 9366 6010
rect 9418 5958 10856 6010
rect 1104 5936 10856 5958
rect 3053 5899 3111 5905
rect 3053 5865 3065 5899
rect 3099 5896 3111 5899
rect 3602 5896 3608 5908
rect 3099 5868 3608 5896
rect 3099 5865 3111 5868
rect 3053 5859 3111 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 4908 5868 8953 5896
rect 1946 5788 1952 5840
rect 2004 5828 2010 5840
rect 4908 5828 4936 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 9674 5856 9680 5908
rect 9732 5896 9738 5908
rect 10045 5899 10103 5905
rect 10045 5896 10057 5899
rect 9732 5868 10057 5896
rect 9732 5856 9738 5868
rect 10045 5865 10057 5868
rect 10091 5865 10103 5899
rect 10045 5859 10103 5865
rect 2004 5800 4936 5828
rect 2004 5788 2010 5800
rect 8202 5788 8208 5840
rect 8260 5828 8266 5840
rect 8570 5828 8576 5840
rect 8260 5800 8576 5828
rect 8260 5788 8266 5800
rect 8570 5788 8576 5800
rect 8628 5828 8634 5840
rect 8628 5800 9260 5828
rect 8628 5788 8634 5800
rect 3418 5760 3424 5772
rect 2148 5732 3424 5760
rect 2038 5692 2044 5704
rect 1999 5664 2044 5692
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2148 5701 2176 5732
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5760 5871 5763
rect 6362 5760 6368 5772
rect 5859 5732 6368 5760
rect 5859 5729 5871 5732
rect 5813 5723 5871 5729
rect 6362 5720 6368 5732
rect 6420 5720 6426 5772
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 8294 5760 8300 5772
rect 7791 5732 8300 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 9232 5769 9260 5800
rect 9217 5763 9275 5769
rect 9217 5729 9229 5763
rect 9263 5729 9275 5763
rect 9398 5760 9404 5772
rect 9359 5732 9404 5760
rect 9217 5723 9275 5729
rect 9398 5720 9404 5732
rect 9456 5720 9462 5772
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2682 5692 2688 5704
rect 2643 5664 2688 5692
rect 2133 5655 2191 5661
rect 2148 5568 2176 5655
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 5258 5692 5264 5704
rect 3344 5664 5264 5692
rect 3344 5636 3372 5664
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5534 5652 5540 5704
rect 5592 5701 5598 5704
rect 5592 5692 5604 5701
rect 7834 5692 7840 5704
rect 5592 5664 5637 5692
rect 5828 5664 7840 5692
rect 5592 5655 5604 5664
rect 5592 5652 5598 5655
rect 2774 5584 2780 5636
rect 2832 5624 2838 5636
rect 3326 5624 3332 5636
rect 2832 5596 3332 5624
rect 2832 5584 2838 5596
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 5828 5624 5856 5664
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 9122 5692 9128 5704
rect 9083 5664 9128 5692
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5692 9367 5695
rect 9490 5692 9496 5704
rect 9355 5664 9496 5692
rect 9355 5661 9367 5664
rect 9309 5655 9367 5661
rect 4120 5596 5856 5624
rect 7500 5627 7558 5633
rect 4120 5584 4126 5596
rect 7500 5593 7512 5627
rect 7546 5624 7558 5627
rect 8202 5624 8208 5636
rect 7546 5596 8208 5624
rect 7546 5593 7558 5596
rect 7500 5587 7558 5593
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 8478 5584 8484 5636
rect 8536 5624 8542 5636
rect 9324 5624 9352 5655
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 9953 5655 10011 5661
rect 8536 5596 9352 5624
rect 8536 5584 8542 5596
rect 1857 5559 1915 5565
rect 1857 5525 1869 5559
rect 1903 5556 1915 5559
rect 1946 5556 1952 5568
rect 1903 5528 1952 5556
rect 1903 5525 1915 5528
rect 1857 5519 1915 5525
rect 1946 5516 1952 5528
rect 2004 5516 2010 5568
rect 2130 5516 2136 5568
rect 2188 5516 2194 5568
rect 2958 5516 2964 5568
rect 3016 5556 3022 5568
rect 3053 5559 3111 5565
rect 3053 5556 3065 5559
rect 3016 5528 3065 5556
rect 3016 5516 3022 5528
rect 3053 5525 3065 5528
rect 3099 5525 3111 5559
rect 3234 5556 3240 5568
rect 3195 5528 3240 5556
rect 3053 5519 3111 5525
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 4433 5559 4491 5565
rect 4433 5556 4445 5559
rect 3936 5528 4445 5556
rect 3936 5516 3942 5528
rect 4433 5525 4445 5528
rect 4479 5525 4491 5559
rect 4433 5519 4491 5525
rect 5350 5516 5356 5568
rect 5408 5556 5414 5568
rect 6365 5559 6423 5565
rect 6365 5556 6377 5559
rect 5408 5528 6377 5556
rect 5408 5516 5414 5528
rect 6365 5525 6377 5528
rect 6411 5525 6423 5559
rect 6365 5519 6423 5525
rect 6638 5516 6644 5568
rect 6696 5556 6702 5568
rect 9968 5556 9996 5655
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 6696 5528 9996 5556
rect 6696 5516 6702 5528
rect 1104 5466 10856 5488
rect 1104 5414 4214 5466
rect 4266 5414 4278 5466
rect 4330 5414 4342 5466
rect 4394 5414 4406 5466
rect 4458 5414 4470 5466
rect 4522 5414 7478 5466
rect 7530 5414 7542 5466
rect 7594 5414 7606 5466
rect 7658 5414 7670 5466
rect 7722 5414 7734 5466
rect 7786 5414 10856 5466
rect 1104 5392 10856 5414
rect 2498 5312 2504 5364
rect 2556 5361 2562 5364
rect 2556 5355 2575 5361
rect 2563 5321 2575 5355
rect 2682 5352 2688 5364
rect 2643 5324 2688 5352
rect 2556 5315 2575 5321
rect 2556 5312 2562 5315
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 3160 5324 5120 5352
rect 2317 5287 2375 5293
rect 2317 5253 2329 5287
rect 2363 5284 2375 5287
rect 2774 5284 2780 5296
rect 2363 5256 2780 5284
rect 2363 5253 2375 5256
rect 2317 5247 2375 5253
rect 2774 5244 2780 5256
rect 2832 5244 2838 5296
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5216 1639 5219
rect 1627 5188 2084 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 1854 5148 1860 5160
rect 1815 5120 1860 5148
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 2056 5148 2084 5188
rect 3160 5214 3188 5324
rect 4246 5284 4252 5296
rect 4159 5256 4252 5284
rect 3236 5219 3294 5225
rect 3236 5214 3248 5219
rect 3160 5186 3248 5214
rect 3236 5185 3248 5186
rect 3282 5185 3294 5219
rect 3418 5216 3424 5228
rect 3379 5188 3424 5216
rect 3236 5179 3294 5185
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 4172 5225 4200 5256
rect 4246 5244 4252 5256
rect 4304 5284 4310 5296
rect 4982 5284 4988 5296
rect 4304 5256 4988 5284
rect 4304 5244 4310 5256
rect 4982 5244 4988 5256
rect 5040 5244 5046 5296
rect 5092 5284 5120 5324
rect 5258 5312 5264 5364
rect 5316 5352 5322 5364
rect 5537 5355 5595 5361
rect 5537 5352 5549 5355
rect 5316 5324 5549 5352
rect 5316 5312 5322 5324
rect 5537 5321 5549 5324
rect 5583 5321 5595 5355
rect 5537 5315 5595 5321
rect 6178 5312 6184 5364
rect 6236 5352 6242 5364
rect 7834 5352 7840 5364
rect 6236 5324 7840 5352
rect 6236 5312 6242 5324
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 7975 5324 8493 5352
rect 5350 5284 5356 5296
rect 5092 5256 5356 5284
rect 5350 5244 5356 5256
rect 5408 5244 5414 5296
rect 5626 5244 5632 5296
rect 5684 5284 5690 5296
rect 7975 5284 8003 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 8754 5352 8760 5364
rect 8715 5324 8760 5352
rect 8481 5315 8539 5321
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 8846 5312 8852 5364
rect 8904 5352 8910 5364
rect 9398 5352 9404 5364
rect 8904 5324 9404 5352
rect 8904 5312 8910 5324
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 5684 5256 8003 5284
rect 5684 5244 5690 5256
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4424 5219 4482 5225
rect 4424 5185 4436 5219
rect 4470 5216 4482 5219
rect 4706 5216 4712 5228
rect 4470 5188 4712 5216
rect 4470 5185 4482 5188
rect 4424 5179 4482 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 6362 5216 6368 5228
rect 6323 5188 6368 5216
rect 6362 5176 6368 5188
rect 6420 5176 6426 5228
rect 6638 5225 6644 5228
rect 6632 5179 6644 5225
rect 6696 5216 6702 5228
rect 6696 5188 6732 5216
rect 6638 5176 6644 5179
rect 6696 5176 6702 5188
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7190 5216 7196 5228
rect 6972 5188 7196 5216
rect 6972 5176 6978 5188
rect 7190 5176 7196 5188
rect 7248 5216 7254 5228
rect 8205 5219 8263 5225
rect 8205 5216 8217 5219
rect 7248 5188 7788 5216
rect 7248 5176 7254 5188
rect 2406 5148 2412 5160
rect 2056 5120 2412 5148
rect 2406 5108 2412 5120
rect 2464 5148 2470 5160
rect 3326 5148 3332 5160
rect 2464 5120 3332 5148
rect 2464 5108 2470 5120
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 3510 5108 3516 5160
rect 3568 5148 3574 5160
rect 3568 5120 3924 5148
rect 3568 5108 3574 5120
rect 1765 5083 1823 5089
rect 1765 5049 1777 5083
rect 1811 5080 1823 5083
rect 3602 5080 3608 5092
rect 1811 5052 3608 5080
rect 1811 5049 1823 5052
rect 1765 5043 1823 5049
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 1673 5015 1731 5021
rect 1673 4981 1685 5015
rect 1719 5012 1731 5015
rect 1946 5012 1952 5024
rect 1719 4984 1952 5012
rect 1719 4981 1731 4984
rect 1673 4975 1731 4981
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 2372 4984 2513 5012
rect 2372 4972 2378 4984
rect 2501 4981 2513 4984
rect 2547 4981 2559 5015
rect 2501 4975 2559 4981
rect 3697 5015 3755 5021
rect 3697 4981 3709 5015
rect 3743 5012 3755 5015
rect 3786 5012 3792 5024
rect 3743 4984 3792 5012
rect 3743 4981 3755 4984
rect 3697 4975 3755 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 3896 5012 3924 5120
rect 7760 5080 7788 5188
rect 8128 5188 8217 5216
rect 7834 5108 7840 5160
rect 7892 5148 7898 5160
rect 8128 5148 8156 5188
rect 8205 5185 8217 5188
rect 8251 5185 8263 5219
rect 8386 5216 8392 5228
rect 8347 5188 8392 5216
rect 8205 5179 8263 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 8573 5219 8631 5225
rect 8573 5216 8585 5219
rect 8496 5188 8585 5216
rect 7892 5120 8156 5148
rect 7892 5108 7898 5120
rect 8496 5080 8524 5188
rect 8573 5185 8585 5188
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 8996 5188 9413 5216
rect 8996 5176 9002 5188
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 9582 5216 9588 5228
rect 9543 5188 9588 5216
rect 9401 5179 9459 5185
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 7760 5052 8524 5080
rect 8570 5040 8576 5092
rect 8628 5080 8634 5092
rect 9122 5080 9128 5092
rect 8628 5052 9128 5080
rect 8628 5040 8634 5052
rect 9122 5040 9128 5052
rect 9180 5080 9186 5092
rect 9217 5083 9275 5089
rect 9217 5080 9229 5083
rect 9180 5052 9229 5080
rect 9180 5040 9186 5052
rect 9217 5049 9229 5052
rect 9263 5049 9275 5083
rect 9217 5043 9275 5049
rect 5166 5012 5172 5024
rect 3896 4984 5172 5012
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 7558 4972 7564 5024
rect 7616 5012 7622 5024
rect 7745 5015 7803 5021
rect 7745 5012 7757 5015
rect 7616 4984 7757 5012
rect 7616 4972 7622 4984
rect 7745 4981 7757 4984
rect 7791 4981 7803 5015
rect 7745 4975 7803 4981
rect 1104 4922 10856 4944
rect 1104 4870 2582 4922
rect 2634 4870 2646 4922
rect 2698 4870 2710 4922
rect 2762 4870 2774 4922
rect 2826 4870 2838 4922
rect 2890 4870 5846 4922
rect 5898 4870 5910 4922
rect 5962 4870 5974 4922
rect 6026 4870 6038 4922
rect 6090 4870 6102 4922
rect 6154 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 9238 4922
rect 9290 4870 9302 4922
rect 9354 4870 9366 4922
rect 9418 4870 10856 4922
rect 1104 4848 10856 4870
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 3145 4811 3203 4817
rect 3145 4808 3157 4811
rect 2556 4780 3157 4808
rect 2556 4768 2562 4780
rect 3145 4777 3157 4780
rect 3191 4777 3203 4811
rect 3145 4771 3203 4777
rect 3418 4768 3424 4820
rect 3476 4808 3482 4820
rect 5442 4808 5448 4820
rect 3476 4780 5448 4808
rect 3476 4768 3482 4780
rect 5442 4768 5448 4780
rect 5500 4808 5506 4820
rect 5629 4811 5687 4817
rect 5629 4808 5641 4811
rect 5500 4780 5641 4808
rect 5500 4768 5506 4780
rect 5629 4777 5641 4780
rect 5675 4777 5687 4811
rect 8202 4808 8208 4820
rect 8163 4780 8208 4808
rect 5629 4771 5687 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8386 4768 8392 4820
rect 8444 4808 8450 4820
rect 9217 4811 9275 4817
rect 9217 4808 9229 4811
rect 8444 4780 9229 4808
rect 8444 4768 8450 4780
rect 9217 4777 9229 4780
rect 9263 4777 9275 4811
rect 9217 4771 9275 4777
rect 1765 4743 1823 4749
rect 1765 4709 1777 4743
rect 1811 4740 1823 4743
rect 2038 4740 2044 4752
rect 1811 4712 2044 4740
rect 1811 4709 1823 4712
rect 1765 4703 1823 4709
rect 2038 4700 2044 4712
rect 2096 4740 2102 4752
rect 2317 4743 2375 4749
rect 2317 4740 2329 4743
rect 2096 4712 2329 4740
rect 2096 4700 2102 4712
rect 2317 4709 2329 4712
rect 2363 4740 2375 4743
rect 3510 4740 3516 4752
rect 2363 4712 3516 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 3510 4700 3516 4712
rect 3568 4700 3574 4752
rect 7374 4700 7380 4752
rect 7432 4740 7438 4752
rect 9769 4743 9827 4749
rect 9769 4740 9781 4743
rect 7432 4712 9781 4740
rect 7432 4700 7438 4712
rect 9769 4709 9781 4712
rect 9815 4709 9827 4743
rect 9769 4703 9827 4709
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4672 2559 4675
rect 2961 4675 3019 4681
rect 2961 4672 2973 4675
rect 2547 4644 2973 4672
rect 2547 4641 2559 4644
rect 2501 4635 2559 4641
rect 2961 4641 2973 4644
rect 3007 4672 3019 4675
rect 4246 4672 4252 4684
rect 3007 4644 3188 4672
rect 4207 4644 4252 4672
rect 3007 4641 3019 4644
rect 2961 4635 3019 4641
rect 1578 4604 1584 4616
rect 1539 4576 1584 4604
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 2130 4564 2136 4616
rect 2188 4604 2194 4616
rect 2225 4607 2283 4613
rect 2225 4604 2237 4607
rect 2188 4576 2237 4604
rect 2188 4564 2194 4576
rect 2225 4573 2237 4576
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2130 4428 2136 4480
rect 2188 4468 2194 4480
rect 2501 4471 2559 4477
rect 2501 4468 2513 4471
rect 2188 4440 2513 4468
rect 2188 4428 2194 4440
rect 2501 4437 2513 4440
rect 2547 4437 2559 4471
rect 2501 4431 2559 4437
rect 2961 4471 3019 4477
rect 2961 4437 2973 4471
rect 3007 4468 3019 4471
rect 3050 4468 3056 4480
rect 3007 4440 3056 4468
rect 3007 4437 3019 4440
rect 2961 4431 3019 4437
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 3160 4468 3188 4644
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8536 4644 9045 4672
rect 8536 4632 8542 4644
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4604 3295 4607
rect 4062 4604 4068 4616
rect 3283 4576 4068 4604
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 5592 4576 8401 4604
rect 5592 4564 5598 4576
rect 8389 4573 8401 4576
rect 8435 4573 8447 4607
rect 9306 4604 9312 4616
rect 9267 4576 9312 4604
rect 8389 4567 8447 4573
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9398 4564 9404 4616
rect 9456 4604 9462 4616
rect 10045 4607 10103 4613
rect 10045 4604 10057 4607
rect 9456 4576 10057 4604
rect 9456 4564 9462 4576
rect 10045 4573 10057 4576
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 4516 4539 4574 4545
rect 4516 4505 4528 4539
rect 4562 4536 4574 4539
rect 4614 4536 4620 4548
rect 4562 4508 4620 4536
rect 4562 4505 4574 4508
rect 4516 4499 4574 4505
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 6632 4539 6690 4545
rect 6632 4505 6644 4539
rect 6678 4536 6690 4539
rect 6914 4536 6920 4548
rect 6678 4508 6920 4536
rect 6678 4505 6690 4508
rect 6632 4499 6690 4505
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 7374 4536 7380 4548
rect 7156 4508 7380 4536
rect 7156 4496 7162 4508
rect 7374 4496 7380 4508
rect 7432 4496 7438 4548
rect 7558 4496 7564 4548
rect 7616 4496 7622 4548
rect 7834 4496 7840 4548
rect 7892 4536 7898 4548
rect 9769 4539 9827 4545
rect 9769 4536 9781 4539
rect 7892 4508 9781 4536
rect 7892 4496 7898 4508
rect 9769 4505 9781 4508
rect 9815 4505 9827 4539
rect 9769 4499 9827 4505
rect 4890 4468 4896 4480
rect 3160 4440 4896 4468
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 7190 4428 7196 4480
rect 7248 4468 7254 4480
rect 7576 4468 7604 4496
rect 7248 4440 7604 4468
rect 7745 4471 7803 4477
rect 7248 4428 7254 4440
rect 7745 4437 7757 4471
rect 7791 4468 7803 4471
rect 8846 4468 8852 4480
rect 7791 4440 8852 4468
rect 7791 4437 7803 4440
rect 7745 4431 7803 4437
rect 8846 4428 8852 4440
rect 8904 4428 8910 4480
rect 9030 4468 9036 4480
rect 8991 4440 9036 4468
rect 9030 4428 9036 4440
rect 9088 4428 9094 4480
rect 9122 4428 9128 4480
rect 9180 4468 9186 4480
rect 9953 4471 10011 4477
rect 9953 4468 9965 4471
rect 9180 4440 9965 4468
rect 9180 4428 9186 4440
rect 9953 4437 9965 4440
rect 9999 4437 10011 4471
rect 9953 4431 10011 4437
rect 1104 4378 10856 4400
rect 1104 4326 4214 4378
rect 4266 4326 4278 4378
rect 4330 4326 4342 4378
rect 4394 4326 4406 4378
rect 4458 4326 4470 4378
rect 4522 4326 7478 4378
rect 7530 4326 7542 4378
rect 7594 4326 7606 4378
rect 7658 4326 7670 4378
rect 7722 4326 7734 4378
rect 7786 4326 10856 4378
rect 1104 4304 10856 4326
rect 1670 4224 1676 4276
rect 1728 4264 1734 4276
rect 2803 4267 2861 4273
rect 2803 4264 2815 4267
rect 1728 4236 2815 4264
rect 1728 4224 1734 4236
rect 2803 4233 2815 4236
rect 2849 4264 2861 4267
rect 3418 4264 3424 4276
rect 2849 4236 3424 4264
rect 2849 4233 2861 4236
rect 2803 4227 2861 4233
rect 3418 4224 3424 4236
rect 3476 4224 3482 4276
rect 3973 4267 4031 4273
rect 3973 4233 3985 4267
rect 4019 4264 4031 4267
rect 5534 4264 5540 4276
rect 4019 4236 5540 4264
rect 4019 4233 4031 4236
rect 3973 4227 4031 4233
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 6822 4224 6828 4276
rect 6880 4264 6886 4276
rect 8386 4264 8392 4276
rect 6880 4236 8392 4264
rect 6880 4224 6886 4236
rect 1762 4156 1768 4208
rect 1820 4196 1826 4208
rect 2590 4196 2596 4208
rect 1820 4168 2596 4196
rect 1820 4156 1826 4168
rect 2590 4156 2596 4168
rect 2648 4156 2654 4208
rect 2958 4156 2964 4208
rect 3016 4196 3022 4208
rect 3789 4199 3847 4205
rect 3789 4196 3801 4199
rect 3016 4168 3801 4196
rect 3016 4156 3022 4168
rect 3789 4165 3801 4168
rect 3835 4196 3847 4199
rect 4246 4196 4252 4208
rect 3835 4168 4252 4196
rect 3835 4165 3847 4168
rect 3789 4159 3847 4165
rect 4246 4156 4252 4168
rect 4304 4156 4310 4208
rect 4982 4196 4988 4208
rect 4448 4168 4988 4196
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 4448 4137 4476 4168
rect 4982 4156 4988 4168
rect 5040 4156 5046 4208
rect 8036 4196 8064 4236
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 8938 4264 8944 4276
rect 8899 4236 8944 4264
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 8036 4168 8156 4196
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4522 4088 4528 4140
rect 4580 4088 4586 4140
rect 4700 4131 4758 4137
rect 4700 4097 4712 4131
rect 4746 4128 4758 4131
rect 6362 4128 6368 4140
rect 4746 4100 6368 4128
rect 4746 4097 4758 4100
rect 4700 4091 4758 4097
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 8128 4137 8156 4168
rect 8113 4131 8171 4137
rect 7116 4100 8064 4128
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4060 2099 4063
rect 4540 4060 4568 4088
rect 2087 4032 4568 4060
rect 2087 4029 2099 4032
rect 2041 4023 2099 4029
rect 3142 3992 3148 4004
rect 2792 3964 3148 3992
rect 2792 3933 2820 3964
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 3421 3995 3479 4001
rect 3421 3961 3433 3995
rect 3467 3992 3479 3995
rect 3970 3992 3976 4004
rect 3467 3964 3976 3992
rect 3467 3961 3479 3964
rect 3421 3955 3479 3961
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 5813 3995 5871 4001
rect 5813 3961 5825 3995
rect 5859 3992 5871 3995
rect 7116 3992 7144 4100
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4060 7527 4063
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7515 4032 7941 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 8036 4060 8064 4100
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 8754 4128 8760 4140
rect 8715 4100 8760 4128
rect 8113 4091 8171 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8996 4100 9045 4128
rect 8996 4088 9002 4100
rect 9033 4097 9045 4100
rect 9079 4128 9091 4131
rect 9398 4128 9404 4140
rect 9079 4100 9404 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 9858 4128 9864 4140
rect 9819 4100 9864 4128
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 8036 4032 8309 4060
rect 7929 4023 7987 4029
rect 8297 4029 8309 4032
rect 8343 4060 8355 4063
rect 9306 4060 9312 4072
rect 8343 4032 9312 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 5859 3964 7144 3992
rect 7208 3992 7236 4023
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 7650 3992 7656 4004
rect 7208 3964 7656 3992
rect 5859 3961 5871 3964
rect 5813 3955 5871 3961
rect 7650 3952 7656 3964
rect 7708 3952 7714 4004
rect 10042 3992 10048 4004
rect 10003 3964 10048 3992
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 2777 3927 2835 3933
rect 2777 3893 2789 3927
rect 2823 3893 2835 3927
rect 2958 3924 2964 3936
rect 2919 3896 2964 3924
rect 2777 3887 2835 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 3786 3924 3792 3936
rect 3747 3896 3792 3924
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 5718 3924 5724 3936
rect 4120 3896 5724 3924
rect 4120 3884 4126 3896
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 7340 3896 8769 3924
rect 7340 3884 7346 3896
rect 8757 3893 8769 3896
rect 8803 3893 8815 3927
rect 8757 3887 8815 3893
rect 1104 3834 10856 3856
rect 1104 3782 2582 3834
rect 2634 3782 2646 3834
rect 2698 3782 2710 3834
rect 2762 3782 2774 3834
rect 2826 3782 2838 3834
rect 2890 3782 5846 3834
rect 5898 3782 5910 3834
rect 5962 3782 5974 3834
rect 6026 3782 6038 3834
rect 6090 3782 6102 3834
rect 6154 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 9238 3834
rect 9290 3782 9302 3834
rect 9354 3782 9366 3834
rect 9418 3782 10856 3834
rect 1104 3760 10856 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 2222 3720 2228 3732
rect 2179 3692 2228 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 2958 3720 2964 3732
rect 2915 3692 2964 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3142 3680 3148 3732
rect 3200 3720 3206 3732
rect 5534 3720 5540 3732
rect 3200 3692 5540 3720
rect 3200 3680 3206 3692
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 6454 3720 6460 3732
rect 6415 3692 6460 3720
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 7098 3720 7104 3732
rect 7059 3692 7104 3720
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 7282 3720 7288 3732
rect 7243 3692 7288 3720
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 8812 3692 9137 3720
rect 8812 3680 8818 3692
rect 9125 3689 9137 3692
rect 9171 3689 9183 3723
rect 9125 3683 9183 3689
rect 5074 3652 5080 3664
rect 2148 3624 5080 3652
rect 2148 3525 2176 3624
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 5350 3612 5356 3664
rect 5408 3612 5414 3664
rect 5629 3655 5687 3661
rect 5629 3621 5641 3655
rect 5675 3652 5687 3655
rect 7190 3652 7196 3664
rect 5675 3624 7196 3652
rect 5675 3621 5687 3624
rect 5629 3615 5687 3621
rect 7190 3612 7196 3624
rect 7248 3612 7254 3664
rect 7558 3652 7564 3664
rect 7392 3624 7564 3652
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 4249 3587 4307 3593
rect 3384 3556 4016 3584
rect 3384 3544 3390 3556
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3485 2375 3519
rect 2317 3479 2375 3485
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3516 3019 3519
rect 3878 3516 3884 3528
rect 3007 3488 3884 3516
rect 3007 3485 3019 3488
rect 2961 3479 3019 3485
rect 2332 3448 2360 3479
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 3988 3516 4016 3556
rect 4249 3553 4261 3587
rect 4295 3584 4307 3587
rect 5368 3584 5396 3612
rect 4295 3556 5396 3584
rect 6089 3587 6147 3593
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 6089 3553 6101 3587
rect 6135 3584 6147 3587
rect 6270 3584 6276 3596
rect 6135 3556 6276 3584
rect 6135 3553 6147 3556
rect 6089 3547 6147 3553
rect 6270 3544 6276 3556
rect 6328 3584 6334 3596
rect 7392 3584 7420 3624
rect 7558 3612 7564 3624
rect 7616 3612 7622 3664
rect 8110 3612 8116 3664
rect 8168 3652 8174 3664
rect 8297 3655 8355 3661
rect 8297 3652 8309 3655
rect 8168 3624 8309 3652
rect 8168 3612 8174 3624
rect 8297 3621 8309 3624
rect 8343 3621 8355 3655
rect 8297 3615 8355 3621
rect 7650 3584 7656 3596
rect 6328 3556 7420 3584
rect 7484 3556 7656 3584
rect 6328 3544 6334 3556
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 3988 3488 4445 3516
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 4890 3476 4896 3528
rect 4948 3516 4954 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 4948 3488 5365 3516
rect 4948 3476 4954 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5500 3488 5545 3516
rect 5500 3476 5506 3488
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 6730 3516 6736 3528
rect 5684 3488 6736 3516
rect 5684 3476 5690 3488
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 7484 3525 7512 3556
rect 7650 3544 7656 3556
rect 7708 3584 7714 3596
rect 8202 3584 8208 3596
rect 7708 3556 8208 3584
rect 7708 3544 7714 3556
rect 8202 3544 8208 3556
rect 8260 3584 8266 3596
rect 8260 3556 8984 3584
rect 8260 3544 8266 3556
rect 8956 3528 8984 3556
rect 7193 3519 7251 3525
rect 7193 3516 7205 3519
rect 7064 3488 7205 3516
rect 7064 3476 7070 3488
rect 7193 3485 7205 3488
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 7800 3488 8033 3516
rect 7800 3476 7806 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 8294 3516 8300 3528
rect 8255 3488 8300 3516
rect 8021 3479 8079 3485
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 8938 3516 8944 3528
rect 8899 3488 8944 3516
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 9088 3488 9137 3516
rect 9088 3476 9094 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 4617 3451 4675 3457
rect 2332 3420 4568 3448
rect 4540 3380 4568 3420
rect 4617 3417 4629 3451
rect 4663 3448 4675 3451
rect 4706 3448 4712 3460
rect 4663 3420 4712 3448
rect 4663 3417 4675 3420
rect 4617 3411 4675 3417
rect 4706 3408 4712 3420
rect 4764 3448 4770 3460
rect 5261 3451 5319 3457
rect 5261 3448 5273 3451
rect 4764 3420 5273 3448
rect 4764 3408 4770 3420
rect 5261 3417 5273 3420
rect 5307 3417 5319 3451
rect 6822 3448 6828 3460
rect 5261 3411 5319 3417
rect 5368 3420 6828 3448
rect 4798 3380 4804 3392
rect 4540 3352 4804 3380
rect 4798 3340 4804 3352
rect 4856 3340 4862 3392
rect 4890 3340 4896 3392
rect 4948 3380 4954 3392
rect 5077 3383 5135 3389
rect 5077 3380 5089 3383
rect 4948 3352 5089 3380
rect 4948 3340 4954 3352
rect 5077 3349 5089 3352
rect 5123 3380 5135 3383
rect 5368 3380 5396 3420
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 7098 3408 7104 3460
rect 7156 3448 7162 3460
rect 7561 3451 7619 3457
rect 7156 3420 7512 3448
rect 7156 3408 7162 3420
rect 6454 3380 6460 3392
rect 5123 3352 5396 3380
rect 6415 3352 6460 3380
rect 5123 3349 5135 3352
rect 5077 3343 5135 3349
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 6641 3383 6699 3389
rect 6641 3349 6653 3383
rect 6687 3380 6699 3383
rect 7374 3380 7380 3392
rect 6687 3352 7380 3380
rect 6687 3349 6699 3352
rect 6641 3343 6699 3349
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 7484 3380 7512 3420
rect 7561 3417 7573 3451
rect 7607 3448 7619 3451
rect 8570 3448 8576 3460
rect 7607 3420 8576 3448
rect 7607 3417 7619 3420
rect 7561 3411 7619 3417
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 8113 3383 8171 3389
rect 8113 3380 8125 3383
rect 7484 3352 8125 3380
rect 8113 3349 8125 3352
rect 8159 3349 8171 3383
rect 8113 3343 8171 3349
rect 1104 3290 10856 3312
rect 1104 3238 4214 3290
rect 4266 3238 4278 3290
rect 4330 3238 4342 3290
rect 4394 3238 4406 3290
rect 4458 3238 4470 3290
rect 4522 3238 7478 3290
rect 7530 3238 7542 3290
rect 7594 3238 7606 3290
rect 7658 3238 7670 3290
rect 7722 3238 7734 3290
rect 7786 3238 10856 3290
rect 1104 3216 10856 3238
rect 3237 3179 3295 3185
rect 3237 3145 3249 3179
rect 3283 3176 3295 3179
rect 4614 3176 4620 3188
rect 3283 3148 4620 3176
rect 3283 3145 3295 3148
rect 3237 3139 3295 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 4706 3136 4712 3188
rect 4764 3185 4770 3188
rect 4764 3179 4783 3185
rect 4771 3145 4783 3179
rect 4764 3139 4783 3145
rect 4764 3136 4770 3139
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 5534 3176 5540 3188
rect 5408 3148 5540 3176
rect 5408 3136 5414 3148
rect 5534 3136 5540 3148
rect 5592 3176 5598 3188
rect 7653 3179 7711 3185
rect 5592 3148 5672 3176
rect 5592 3136 5598 3148
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 4525 3111 4583 3117
rect 2004 3080 4108 3108
rect 2004 3068 2010 3080
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3040 3111 3043
rect 3234 3040 3240 3052
rect 3099 3012 3240 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3602 3000 3608 3052
rect 3660 3040 3666 3052
rect 4080 3049 4108 3080
rect 4525 3077 4537 3111
rect 4571 3108 4583 3111
rect 5442 3108 5448 3120
rect 4571 3080 5448 3108
rect 4571 3077 4583 3080
rect 4525 3071 4583 3077
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 3789 3043 3847 3049
rect 3789 3040 3801 3043
rect 3660 3012 3801 3040
rect 3660 3000 3666 3012
rect 3789 3009 3801 3012
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 3326 2932 3332 2984
rect 3384 2972 3390 2984
rect 3988 2972 4016 3003
rect 4798 3000 4804 3052
rect 4856 3040 4862 3052
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 4856 3012 5365 3040
rect 4856 3000 4862 3012
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5534 3040 5540 3052
rect 5495 3012 5540 3040
rect 5353 3003 5411 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5644 3049 5672 3148
rect 7653 3145 7665 3179
rect 7699 3176 7711 3179
rect 7834 3176 7840 3188
rect 7699 3148 7840 3176
rect 7699 3145 7711 3148
rect 7653 3139 7711 3145
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8386 3176 8392 3188
rect 7943 3148 8392 3176
rect 6454 3068 6460 3120
rect 6512 3108 6518 3120
rect 7943 3108 7971 3148
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 8573 3179 8631 3185
rect 8573 3176 8585 3179
rect 8536 3148 8585 3176
rect 8536 3136 8542 3148
rect 8573 3145 8585 3148
rect 8619 3145 8631 3179
rect 8573 3139 8631 3145
rect 8846 3108 8852 3120
rect 6512 3080 7971 3108
rect 8222 3080 8852 3108
rect 6512 3068 6518 3080
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3009 5687 3043
rect 7190 3040 7196 3052
rect 7151 3012 7196 3040
rect 5629 3003 5687 3009
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3038 7987 3043
rect 8222 3040 8250 3080
rect 8846 3068 8852 3080
rect 8904 3068 8910 3120
rect 8386 3040 8392 3052
rect 8036 3038 8250 3040
rect 7975 3012 8250 3038
rect 8347 3012 8392 3040
rect 7975 3010 8064 3012
rect 7975 3009 7987 3010
rect 7929 3003 7987 3009
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 3384 2944 4016 2972
rect 3384 2932 3390 2944
rect 4982 2932 4988 2984
rect 5040 2972 5046 2984
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 5040 2944 6929 2972
rect 5040 2932 5046 2944
rect 6917 2941 6929 2944
rect 6963 2972 6975 2975
rect 7650 2972 7656 2984
rect 6963 2944 7236 2972
rect 7611 2944 7656 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 3694 2864 3700 2916
rect 3752 2904 3758 2916
rect 3789 2907 3847 2913
rect 3789 2904 3801 2907
rect 3752 2876 3801 2904
rect 3752 2864 3758 2876
rect 3789 2873 3801 2876
rect 3835 2873 3847 2907
rect 3789 2867 3847 2873
rect 3970 2864 3976 2916
rect 4028 2904 4034 2916
rect 4893 2907 4951 2913
rect 4893 2904 4905 2907
rect 4028 2876 4905 2904
rect 4028 2864 4034 2876
rect 4893 2873 4905 2876
rect 4939 2904 4951 2907
rect 7101 2907 7159 2913
rect 7101 2904 7113 2907
rect 4939 2876 7113 2904
rect 4939 2873 4951 2876
rect 4893 2867 4951 2873
rect 7101 2873 7113 2876
rect 7147 2873 7159 2907
rect 7208 2904 7236 2944
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 8478 2972 8484 2984
rect 7760 2944 8484 2972
rect 7760 2904 7788 2944
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 7208 2876 7788 2904
rect 7837 2907 7895 2913
rect 7101 2867 7159 2873
rect 7837 2873 7849 2907
rect 7883 2904 7895 2907
rect 8202 2904 8208 2916
rect 7883 2876 8208 2904
rect 7883 2873 7895 2876
rect 7837 2867 7895 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 5166 2836 5172 2848
rect 4764 2808 5172 2836
rect 4764 2796 4770 2808
rect 5166 2796 5172 2808
rect 5224 2796 5230 2848
rect 7006 2836 7012 2848
rect 6967 2808 7012 2836
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 1104 2746 10856 2768
rect 1104 2694 2582 2746
rect 2634 2694 2646 2746
rect 2698 2694 2710 2746
rect 2762 2694 2774 2746
rect 2826 2694 2838 2746
rect 2890 2694 5846 2746
rect 5898 2694 5910 2746
rect 5962 2694 5974 2746
rect 6026 2694 6038 2746
rect 6090 2694 6102 2746
rect 6154 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 9238 2746
rect 9290 2694 9302 2746
rect 9354 2694 9366 2746
rect 9418 2694 10856 2746
rect 1104 2672 10856 2694
rect 4246 2632 4252 2644
rect 4207 2604 4252 2632
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2632 4399 2635
rect 4798 2632 4804 2644
rect 4387 2604 4804 2632
rect 4387 2601 4399 2604
rect 4341 2595 4399 2601
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 5074 2632 5080 2644
rect 5035 2604 5080 2632
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5169 2635 5227 2641
rect 5169 2601 5181 2635
rect 5215 2632 5227 2635
rect 5534 2632 5540 2644
rect 5215 2604 5540 2632
rect 5215 2601 5227 2604
rect 5169 2595 5227 2601
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 6270 2592 6276 2644
rect 6328 2632 6334 2644
rect 6549 2635 6607 2641
rect 6549 2632 6561 2635
rect 6328 2604 6561 2632
rect 6328 2592 6334 2604
rect 6549 2601 6561 2604
rect 6595 2601 6607 2635
rect 6549 2595 6607 2601
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 7101 2635 7159 2641
rect 7101 2632 7113 2635
rect 6972 2604 7113 2632
rect 6972 2592 6978 2604
rect 7101 2601 7113 2604
rect 7147 2601 7159 2635
rect 7101 2595 7159 2601
rect 7929 2635 7987 2641
rect 7929 2601 7941 2635
rect 7975 2632 7987 2635
rect 8662 2632 8668 2644
rect 7975 2604 8668 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 4890 2564 4896 2576
rect 2424 2536 4896 2564
rect 2424 2437 2452 2536
rect 4890 2524 4896 2536
rect 4948 2524 4954 2576
rect 5258 2524 5264 2576
rect 5316 2524 5322 2576
rect 6457 2567 6515 2573
rect 6457 2533 6469 2567
rect 6503 2564 6515 2567
rect 8018 2564 8024 2576
rect 6503 2536 8024 2564
rect 6503 2533 6515 2536
rect 6457 2527 6515 2533
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 4157 2499 4215 2505
rect 4157 2496 4169 2499
rect 2532 2468 4169 2496
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 1854 2320 1860 2372
rect 1912 2360 1918 2372
rect 2532 2360 2560 2468
rect 4157 2465 4169 2468
rect 4203 2465 4215 2499
rect 4982 2496 4988 2508
rect 4943 2468 4988 2496
rect 4157 2459 4215 2465
rect 4982 2456 4988 2468
rect 5040 2456 5046 2508
rect 5276 2496 5304 2524
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 5276 2468 6377 2496
rect 6365 2465 6377 2468
rect 6411 2496 6423 2499
rect 7650 2496 7656 2508
rect 6411 2468 7656 2496
rect 6411 2465 6423 2468
rect 6365 2459 6423 2465
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2397 2651 2431
rect 3050 2428 3056 2440
rect 3011 2400 3056 2428
rect 2593 2391 2651 2397
rect 1912 2332 2560 2360
rect 2608 2360 2636 2391
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 4246 2428 4252 2440
rect 3283 2400 4252 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 4430 2388 4436 2440
rect 4488 2428 4494 2440
rect 5261 2431 5319 2437
rect 4488 2400 4533 2428
rect 4488 2388 4494 2400
rect 5261 2397 5273 2431
rect 5307 2428 5319 2431
rect 5350 2428 5356 2440
rect 5307 2400 5356 2428
rect 5307 2397 5319 2400
rect 5261 2391 5319 2397
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 7098 2428 7104 2440
rect 6687 2400 7104 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7282 2428 7288 2440
rect 7243 2400 7288 2428
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 7524 2400 7757 2428
rect 7524 2388 7530 2400
rect 7745 2397 7757 2400
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 3145 2363 3203 2369
rect 2608 2332 2774 2360
rect 1912 2320 1918 2332
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 2746 2292 2774 2332
rect 3145 2329 3157 2363
rect 3191 2360 3203 2363
rect 6546 2360 6552 2372
rect 3191 2332 6552 2360
rect 3191 2329 3203 2332
rect 3145 2323 3203 2329
rect 6546 2320 6552 2332
rect 6604 2320 6610 2372
rect 7006 2292 7012 2304
rect 2746 2264 7012 2292
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 1104 2202 10856 2224
rect 1104 2150 4214 2202
rect 4266 2150 4278 2202
rect 4330 2150 4342 2202
rect 4394 2150 4406 2202
rect 4458 2150 4470 2202
rect 4522 2150 7478 2202
rect 7530 2150 7542 2202
rect 7594 2150 7606 2202
rect 7658 2150 7670 2202
rect 7722 2150 7734 2202
rect 7786 2150 10856 2202
rect 1104 2128 10856 2150
rect 2498 2048 2504 2100
rect 2556 2088 2562 2100
rect 6638 2088 6644 2100
rect 2556 2060 6644 2088
rect 2556 2048 2562 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
<< via1 >>
rect 5448 11500 5500 11552
rect 10140 11500 10192 11552
rect 2582 11398 2634 11450
rect 2646 11398 2698 11450
rect 2710 11398 2762 11450
rect 2774 11398 2826 11450
rect 2838 11398 2890 11450
rect 5846 11398 5898 11450
rect 5910 11398 5962 11450
rect 5974 11398 6026 11450
rect 6038 11398 6090 11450
rect 6102 11398 6154 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 9238 11398 9290 11450
rect 9302 11398 9354 11450
rect 9366 11398 9418 11450
rect 4804 11296 4856 11348
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 8116 11296 8168 11348
rect 3976 11271 4028 11280
rect 3976 11237 3985 11271
rect 3985 11237 4019 11271
rect 4019 11237 4028 11271
rect 3976 11228 4028 11237
rect 5172 11228 5224 11280
rect 9128 11228 9180 11280
rect 4528 11160 4580 11212
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 3240 11092 3292 11101
rect 3792 11135 3844 11144
rect 3792 11101 3801 11135
rect 3801 11101 3835 11135
rect 3835 11101 3844 11135
rect 3792 11092 3844 11101
rect 4160 11092 4212 11144
rect 4988 11092 5040 11144
rect 5356 11092 5408 11144
rect 6828 11160 6880 11212
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 8760 11160 8812 11212
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 3148 11067 3200 11076
rect 3148 11033 3157 11067
rect 3157 11033 3191 11067
rect 3191 11033 3200 11067
rect 3148 11024 3200 11033
rect 8484 11024 8536 11076
rect 1400 10999 1452 11008
rect 1400 10965 1409 10999
rect 1409 10965 1443 10999
rect 1443 10965 1452 10999
rect 1400 10956 1452 10965
rect 4896 10956 4948 11008
rect 5264 10999 5316 11008
rect 5264 10965 5289 10999
rect 5289 10965 5316 10999
rect 5264 10956 5316 10965
rect 6552 10956 6604 11008
rect 4214 10854 4266 10906
rect 4278 10854 4330 10906
rect 4342 10854 4394 10906
rect 4406 10854 4458 10906
rect 4470 10854 4522 10906
rect 7478 10854 7530 10906
rect 7542 10854 7594 10906
rect 7606 10854 7658 10906
rect 7670 10854 7722 10906
rect 7734 10854 7786 10906
rect 1768 10684 1820 10736
rect 5080 10727 5132 10736
rect 5080 10693 5089 10727
rect 5089 10693 5123 10727
rect 5123 10693 5132 10727
rect 5080 10684 5132 10693
rect 6368 10684 6420 10736
rect 8208 10752 8260 10804
rect 2504 10616 2556 10668
rect 4436 10616 4488 10668
rect 4528 10616 4580 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 3976 10591 4028 10600
rect 3332 10480 3384 10532
rect 3976 10557 3985 10591
rect 3985 10557 4019 10591
rect 4019 10557 4028 10591
rect 3976 10548 4028 10557
rect 4896 10616 4948 10668
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 8668 10684 8720 10736
rect 8024 10616 8076 10668
rect 9128 10659 9180 10668
rect 7104 10548 7156 10600
rect 4896 10480 4948 10532
rect 5264 10480 5316 10532
rect 6920 10523 6972 10532
rect 6920 10489 6929 10523
rect 6929 10489 6963 10523
rect 6963 10489 6972 10523
rect 6920 10480 6972 10489
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 3056 10412 3108 10464
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 4620 10412 4672 10464
rect 5540 10412 5592 10464
rect 6276 10412 6328 10464
rect 7472 10412 7524 10464
rect 8300 10412 8352 10464
rect 8944 10455 8996 10464
rect 8944 10421 8953 10455
rect 8953 10421 8987 10455
rect 8987 10421 8996 10455
rect 8944 10412 8996 10421
rect 2582 10310 2634 10362
rect 2646 10310 2698 10362
rect 2710 10310 2762 10362
rect 2774 10310 2826 10362
rect 2838 10310 2890 10362
rect 5846 10310 5898 10362
rect 5910 10310 5962 10362
rect 5974 10310 6026 10362
rect 6038 10310 6090 10362
rect 6102 10310 6154 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 9238 10310 9290 10362
rect 9302 10310 9354 10362
rect 9366 10310 9418 10362
rect 3516 10208 3568 10260
rect 2320 10140 2372 10192
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 4068 10072 4120 10124
rect 4160 10072 4212 10124
rect 5448 10208 5500 10260
rect 7932 10208 7984 10260
rect 8668 10208 8720 10260
rect 6736 10140 6788 10192
rect 4896 10072 4948 10124
rect 7104 10072 7156 10124
rect 7840 10072 7892 10124
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 2504 10004 2556 10056
rect 3424 10004 3476 10056
rect 3608 9936 3660 9988
rect 2596 9911 2648 9920
rect 2596 9877 2605 9911
rect 2605 9877 2639 9911
rect 2639 9877 2648 9911
rect 2596 9868 2648 9877
rect 3240 9868 3292 9920
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 7012 10004 7064 10056
rect 7472 10047 7524 10056
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 7564 10004 7616 10056
rect 8208 10072 8260 10124
rect 8576 10004 8628 10056
rect 4436 9936 4488 9988
rect 6184 9868 6236 9920
rect 9220 10004 9272 10056
rect 8392 9868 8444 9920
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 9588 9868 9640 9920
rect 4214 9766 4266 9818
rect 4278 9766 4330 9818
rect 4342 9766 4394 9818
rect 4406 9766 4458 9818
rect 4470 9766 4522 9818
rect 7478 9766 7530 9818
rect 7542 9766 7594 9818
rect 7606 9766 7658 9818
rect 7670 9766 7722 9818
rect 7734 9766 7786 9818
rect 2596 9664 2648 9716
rect 1676 9528 1728 9580
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 3332 9596 3384 9648
rect 2964 9528 3016 9580
rect 3516 9596 3568 9648
rect 5080 9664 5132 9716
rect 3700 9571 3752 9580
rect 3700 9537 3709 9571
rect 3709 9537 3743 9571
rect 3743 9537 3752 9571
rect 3700 9528 3752 9537
rect 3976 9571 4028 9580
rect 3976 9537 3985 9571
rect 3985 9537 4019 9571
rect 4019 9537 4028 9571
rect 3976 9528 4028 9537
rect 4160 9528 4212 9580
rect 4988 9596 5040 9648
rect 5264 9596 5316 9648
rect 6460 9664 6512 9716
rect 8576 9664 8628 9716
rect 8668 9664 8720 9716
rect 7104 9596 7156 9648
rect 8300 9596 8352 9648
rect 4528 9528 4580 9580
rect 6552 9528 6604 9580
rect 1952 9392 2004 9444
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 2320 9367 2372 9376
rect 2320 9333 2329 9367
rect 2329 9333 2363 9367
rect 2363 9333 2372 9367
rect 2320 9324 2372 9333
rect 3424 9460 3476 9512
rect 7748 9503 7800 9512
rect 7748 9469 7757 9503
rect 7757 9469 7791 9503
rect 7791 9469 7800 9503
rect 7748 9460 7800 9469
rect 8300 9460 8352 9512
rect 8852 9596 8904 9648
rect 9220 9639 9272 9648
rect 9220 9605 9229 9639
rect 9229 9605 9263 9639
rect 9263 9605 9272 9639
rect 9220 9596 9272 9605
rect 8576 9571 8628 9580
rect 8576 9537 8585 9571
rect 8585 9537 8619 9571
rect 8619 9537 8628 9571
rect 8576 9528 8628 9537
rect 8760 9528 8812 9580
rect 9128 9460 9180 9512
rect 9496 9392 9548 9444
rect 3424 9324 3476 9376
rect 3608 9324 3660 9376
rect 6184 9324 6236 9376
rect 6460 9324 6512 9376
rect 2582 9222 2634 9274
rect 2646 9222 2698 9274
rect 2710 9222 2762 9274
rect 2774 9222 2826 9274
rect 2838 9222 2890 9274
rect 5846 9222 5898 9274
rect 5910 9222 5962 9274
rect 5974 9222 6026 9274
rect 6038 9222 6090 9274
rect 6102 9222 6154 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 9238 9222 9290 9274
rect 9302 9222 9354 9274
rect 9366 9222 9418 9274
rect 2136 9120 2188 9172
rect 2780 8984 2832 9036
rect 1400 8916 1452 8968
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 2504 8916 2556 8968
rect 3792 9120 3844 9172
rect 4252 9120 4304 9172
rect 5632 9120 5684 9172
rect 8668 9120 8720 9172
rect 3332 9052 3384 9104
rect 4620 9052 4672 9104
rect 6828 9095 6880 9104
rect 6828 9061 6837 9095
rect 6837 9061 6871 9095
rect 6871 9061 6880 9095
rect 6828 9052 6880 9061
rect 8852 9052 8904 9104
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 8392 8984 8444 9036
rect 2964 8916 3016 8968
rect 5080 8916 5132 8968
rect 1584 8848 1636 8900
rect 1676 8780 1728 8832
rect 3516 8780 3568 8832
rect 4068 8780 4120 8832
rect 4620 8848 4672 8900
rect 5356 8848 5408 8900
rect 7748 8848 7800 8900
rect 8116 8916 8168 8968
rect 8300 8916 8352 8968
rect 9588 8984 9640 9036
rect 9496 8959 9548 8968
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 10140 8959 10192 8968
rect 9496 8916 9548 8925
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 8944 8848 8996 8900
rect 4896 8780 4948 8832
rect 7288 8780 7340 8832
rect 8484 8780 8536 8832
rect 4214 8678 4266 8730
rect 4278 8678 4330 8730
rect 4342 8678 4394 8730
rect 4406 8678 4458 8730
rect 4470 8678 4522 8730
rect 7478 8678 7530 8730
rect 7542 8678 7594 8730
rect 7606 8678 7658 8730
rect 7670 8678 7722 8730
rect 7734 8678 7786 8730
rect 1400 8576 1452 8628
rect 1768 8551 1820 8560
rect 1768 8517 1777 8551
rect 1777 8517 1811 8551
rect 1811 8517 1820 8551
rect 1768 8508 1820 8517
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 2320 8440 2372 8492
rect 1860 8236 1912 8288
rect 3424 8576 3476 8628
rect 3516 8576 3568 8628
rect 4712 8576 4764 8628
rect 4896 8576 4948 8628
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 4988 8508 5040 8560
rect 9036 8576 9088 8628
rect 8116 8508 8168 8560
rect 3792 8372 3844 8424
rect 4712 8440 4764 8492
rect 4896 8440 4948 8492
rect 5264 8440 5316 8492
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 9496 8440 9548 8492
rect 9588 8415 9640 8424
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 5724 8347 5776 8356
rect 5724 8313 5733 8347
rect 5733 8313 5767 8347
rect 5767 8313 5776 8347
rect 5724 8304 5776 8313
rect 7840 8304 7892 8356
rect 8392 8304 8444 8356
rect 4160 8236 4212 8288
rect 5448 8236 5500 8288
rect 8484 8236 8536 8288
rect 2582 8134 2634 8186
rect 2646 8134 2698 8186
rect 2710 8134 2762 8186
rect 2774 8134 2826 8186
rect 2838 8134 2890 8186
rect 5846 8134 5898 8186
rect 5910 8134 5962 8186
rect 5974 8134 6026 8186
rect 6038 8134 6090 8186
rect 6102 8134 6154 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 9238 8134 9290 8186
rect 9302 8134 9354 8186
rect 9366 8134 9418 8186
rect 2964 8032 3016 8084
rect 4160 8032 4212 8084
rect 5080 8032 5132 8084
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 1860 7896 1912 7948
rect 3240 7939 3292 7948
rect 3240 7905 3249 7939
rect 3249 7905 3283 7939
rect 3283 7905 3292 7939
rect 3240 7896 3292 7905
rect 7748 7896 7800 7948
rect 8484 7964 8536 8016
rect 2044 7828 2096 7880
rect 3332 7828 3384 7880
rect 7012 7871 7064 7880
rect 7012 7837 7030 7871
rect 7030 7837 7064 7871
rect 7012 7828 7064 7837
rect 9036 7828 9088 7880
rect 4620 7760 4672 7812
rect 4988 7760 5040 7812
rect 5172 7803 5224 7812
rect 5172 7769 5190 7803
rect 5190 7769 5224 7803
rect 5172 7760 5224 7769
rect 8852 7760 8904 7812
rect 7196 7692 7248 7744
rect 7840 7692 7892 7744
rect 8484 7692 8536 7744
rect 4214 7590 4266 7642
rect 4278 7590 4330 7642
rect 4342 7590 4394 7642
rect 4406 7590 4458 7642
rect 4470 7590 4522 7642
rect 7478 7590 7530 7642
rect 7542 7590 7594 7642
rect 7606 7590 7658 7642
rect 7670 7590 7722 7642
rect 7734 7590 7786 7642
rect 2044 7488 2096 7540
rect 5080 7488 5132 7540
rect 8208 7531 8260 7540
rect 8208 7497 8217 7531
rect 8217 7497 8251 7531
rect 8251 7497 8260 7531
rect 8208 7488 8260 7497
rect 1952 7420 2004 7472
rect 3148 7420 3200 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 4988 7420 5040 7472
rect 7840 7420 7892 7472
rect 8300 7420 8352 7472
rect 8668 7420 8720 7472
rect 7380 7352 7432 7404
rect 9588 7395 9640 7404
rect 9588 7361 9597 7395
rect 9597 7361 9631 7395
rect 9631 7361 9640 7395
rect 9588 7352 9640 7361
rect 6368 7327 6420 7336
rect 1768 7148 1820 7200
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 8944 7148 8996 7200
rect 2582 7046 2634 7098
rect 2646 7046 2698 7098
rect 2710 7046 2762 7098
rect 2774 7046 2826 7098
rect 2838 7046 2890 7098
rect 5846 7046 5898 7098
rect 5910 7046 5962 7098
rect 5974 7046 6026 7098
rect 6038 7046 6090 7098
rect 6102 7046 6154 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 9238 7046 9290 7098
rect 9302 7046 9354 7098
rect 9366 7046 9418 7098
rect 1860 6944 1912 6996
rect 4068 6944 4120 6996
rect 4160 6876 4212 6928
rect 4988 6944 5040 6996
rect 8300 6876 8352 6928
rect 9588 6876 9640 6928
rect 5632 6808 5684 6860
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 2228 6672 2280 6724
rect 3884 6672 3936 6724
rect 7840 6740 7892 6792
rect 3148 6604 3200 6656
rect 3332 6604 3384 6656
rect 3700 6604 3752 6656
rect 5724 6672 5776 6724
rect 9312 6808 9364 6860
rect 9404 6740 9456 6792
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 9588 6604 9640 6656
rect 4214 6502 4266 6554
rect 4278 6502 4330 6554
rect 4342 6502 4394 6554
rect 4406 6502 4458 6554
rect 4470 6502 4522 6554
rect 7478 6502 7530 6554
rect 7542 6502 7594 6554
rect 7606 6502 7658 6554
rect 7670 6502 7722 6554
rect 7734 6502 7786 6554
rect 2320 6400 2372 6452
rect 10140 6400 10192 6452
rect 2964 6332 3016 6384
rect 6368 6332 6420 6384
rect 3700 6307 3752 6316
rect 3700 6273 3718 6307
rect 3718 6273 3752 6307
rect 3700 6264 3752 6273
rect 4988 6264 5040 6316
rect 9588 6332 9640 6384
rect 6552 6264 6604 6316
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 1676 6128 1728 6180
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 2136 6103 2188 6112
rect 2136 6069 2145 6103
rect 2145 6069 2179 6103
rect 2179 6069 2188 6103
rect 2136 6060 2188 6069
rect 2412 6060 2464 6112
rect 3976 6060 4028 6112
rect 4712 6060 4764 6112
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 8576 6060 8628 6112
rect 9864 6060 9916 6112
rect 2582 5958 2634 6010
rect 2646 5958 2698 6010
rect 2710 5958 2762 6010
rect 2774 5958 2826 6010
rect 2838 5958 2890 6010
rect 5846 5958 5898 6010
rect 5910 5958 5962 6010
rect 5974 5958 6026 6010
rect 6038 5958 6090 6010
rect 6102 5958 6154 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 9238 5958 9290 6010
rect 9302 5958 9354 6010
rect 9366 5958 9418 6010
rect 3608 5856 3660 5908
rect 1952 5788 2004 5840
rect 9680 5856 9732 5908
rect 8208 5788 8260 5840
rect 8576 5788 8628 5840
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 3424 5720 3476 5772
rect 6368 5720 6420 5772
rect 8300 5720 8352 5772
rect 9404 5763 9456 5772
rect 9404 5729 9413 5763
rect 9413 5729 9447 5763
rect 9447 5729 9456 5763
rect 9404 5720 9456 5729
rect 2688 5695 2740 5704
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 5264 5652 5316 5704
rect 5540 5695 5592 5704
rect 5540 5661 5558 5695
rect 5558 5661 5592 5695
rect 5540 5652 5592 5661
rect 2780 5584 2832 5636
rect 3332 5584 3384 5636
rect 4068 5584 4120 5636
rect 7840 5652 7892 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 8208 5584 8260 5636
rect 8484 5584 8536 5636
rect 9496 5652 9548 5704
rect 10140 5695 10192 5704
rect 1952 5516 2004 5568
rect 2136 5516 2188 5568
rect 2964 5516 3016 5568
rect 3240 5559 3292 5568
rect 3240 5525 3249 5559
rect 3249 5525 3283 5559
rect 3283 5525 3292 5559
rect 3240 5516 3292 5525
rect 3884 5516 3936 5568
rect 5356 5516 5408 5568
rect 6644 5516 6696 5568
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 4214 5414 4266 5466
rect 4278 5414 4330 5466
rect 4342 5414 4394 5466
rect 4406 5414 4458 5466
rect 4470 5414 4522 5466
rect 7478 5414 7530 5466
rect 7542 5414 7594 5466
rect 7606 5414 7658 5466
rect 7670 5414 7722 5466
rect 7734 5414 7786 5466
rect 2504 5355 2556 5364
rect 2504 5321 2529 5355
rect 2529 5321 2556 5355
rect 2688 5355 2740 5364
rect 2504 5312 2556 5321
rect 2688 5321 2697 5355
rect 2697 5321 2731 5355
rect 2731 5321 2740 5355
rect 2688 5312 2740 5321
rect 2780 5244 2832 5296
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 4252 5244 4304 5296
rect 4988 5244 5040 5296
rect 5264 5312 5316 5364
rect 6184 5312 6236 5364
rect 7840 5312 7892 5364
rect 5356 5244 5408 5296
rect 5632 5244 5684 5296
rect 8760 5355 8812 5364
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 8852 5312 8904 5364
rect 9404 5312 9456 5364
rect 4712 5176 4764 5228
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 6644 5219 6696 5228
rect 6644 5185 6678 5219
rect 6678 5185 6696 5219
rect 6644 5176 6696 5185
rect 6920 5176 6972 5228
rect 7196 5176 7248 5228
rect 2412 5108 2464 5160
rect 3332 5151 3384 5160
rect 3332 5117 3341 5151
rect 3341 5117 3375 5151
rect 3375 5117 3384 5151
rect 3332 5108 3384 5117
rect 3516 5151 3568 5160
rect 3516 5117 3525 5151
rect 3525 5117 3559 5151
rect 3559 5117 3568 5151
rect 3516 5108 3568 5117
rect 3608 5040 3660 5092
rect 1952 4972 2004 5024
rect 2320 4972 2372 5024
rect 3792 4972 3844 5024
rect 7840 5108 7892 5160
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 8944 5176 8996 5228
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 8576 5040 8628 5092
rect 9128 5040 9180 5092
rect 5172 4972 5224 5024
rect 7564 4972 7616 5024
rect 2582 4870 2634 4922
rect 2646 4870 2698 4922
rect 2710 4870 2762 4922
rect 2774 4870 2826 4922
rect 2838 4870 2890 4922
rect 5846 4870 5898 4922
rect 5910 4870 5962 4922
rect 5974 4870 6026 4922
rect 6038 4870 6090 4922
rect 6102 4870 6154 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 9238 4870 9290 4922
rect 9302 4870 9354 4922
rect 9366 4870 9418 4922
rect 2504 4768 2556 4820
rect 3424 4768 3476 4820
rect 5448 4768 5500 4820
rect 8208 4811 8260 4820
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 8392 4768 8444 4820
rect 2044 4700 2096 4752
rect 3516 4700 3568 4752
rect 7380 4700 7432 4752
rect 4252 4675 4304 4684
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 2136 4564 2188 4616
rect 2136 4428 2188 4480
rect 3056 4428 3108 4480
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 8484 4632 8536 4684
rect 4068 4564 4120 4616
rect 5540 4564 5592 4616
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 9404 4564 9456 4616
rect 4620 4496 4672 4548
rect 6920 4496 6972 4548
rect 7104 4496 7156 4548
rect 7380 4496 7432 4548
rect 7564 4496 7616 4548
rect 7840 4496 7892 4548
rect 4896 4428 4948 4480
rect 7196 4428 7248 4480
rect 8852 4428 8904 4480
rect 9036 4471 9088 4480
rect 9036 4437 9045 4471
rect 9045 4437 9079 4471
rect 9079 4437 9088 4471
rect 9036 4428 9088 4437
rect 9128 4428 9180 4480
rect 4214 4326 4266 4378
rect 4278 4326 4330 4378
rect 4342 4326 4394 4378
rect 4406 4326 4458 4378
rect 4470 4326 4522 4378
rect 7478 4326 7530 4378
rect 7542 4326 7594 4378
rect 7606 4326 7658 4378
rect 7670 4326 7722 4378
rect 7734 4326 7786 4378
rect 1676 4224 1728 4276
rect 3424 4224 3476 4276
rect 5540 4224 5592 4276
rect 6828 4224 6880 4276
rect 1768 4156 1820 4208
rect 2596 4199 2648 4208
rect 2596 4165 2605 4199
rect 2605 4165 2639 4199
rect 2639 4165 2648 4199
rect 2596 4156 2648 4165
rect 2964 4156 3016 4208
rect 4252 4156 4304 4208
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 4988 4156 5040 4208
rect 8392 4224 8444 4276
rect 8944 4267 8996 4276
rect 8944 4233 8953 4267
rect 8953 4233 8987 4267
rect 8987 4233 8996 4267
rect 8944 4224 8996 4233
rect 4528 4088 4580 4140
rect 6368 4088 6420 4140
rect 3148 3952 3200 4004
rect 3976 3952 4028 4004
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 8944 4088 8996 4140
rect 9404 4088 9456 4140
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 9312 4020 9364 4072
rect 7656 3952 7708 4004
rect 10048 3995 10100 4004
rect 10048 3961 10057 3995
rect 10057 3961 10091 3995
rect 10091 3961 10100 3995
rect 10048 3952 10100 3961
rect 2964 3927 3016 3936
rect 2964 3893 2973 3927
rect 2973 3893 3007 3927
rect 3007 3893 3016 3927
rect 2964 3884 3016 3893
rect 3792 3927 3844 3936
rect 3792 3893 3801 3927
rect 3801 3893 3835 3927
rect 3835 3893 3844 3927
rect 3792 3884 3844 3893
rect 4068 3884 4120 3936
rect 5724 3884 5776 3936
rect 7288 3884 7340 3936
rect 2582 3782 2634 3834
rect 2646 3782 2698 3834
rect 2710 3782 2762 3834
rect 2774 3782 2826 3834
rect 2838 3782 2890 3834
rect 5846 3782 5898 3834
rect 5910 3782 5962 3834
rect 5974 3782 6026 3834
rect 6038 3782 6090 3834
rect 6102 3782 6154 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 9238 3782 9290 3834
rect 9302 3782 9354 3834
rect 9366 3782 9418 3834
rect 2228 3680 2280 3732
rect 2964 3680 3016 3732
rect 3148 3680 3200 3732
rect 5540 3680 5592 3732
rect 6460 3723 6512 3732
rect 6460 3689 6469 3723
rect 6469 3689 6503 3723
rect 6503 3689 6512 3723
rect 6460 3680 6512 3689
rect 7104 3723 7156 3732
rect 7104 3689 7113 3723
rect 7113 3689 7147 3723
rect 7147 3689 7156 3723
rect 7104 3680 7156 3689
rect 7288 3723 7340 3732
rect 7288 3689 7297 3723
rect 7297 3689 7331 3723
rect 7331 3689 7340 3723
rect 7288 3680 7340 3689
rect 8760 3680 8812 3732
rect 5080 3612 5132 3664
rect 5356 3612 5408 3664
rect 7196 3612 7248 3664
rect 3332 3544 3384 3596
rect 3884 3476 3936 3528
rect 6276 3544 6328 3596
rect 7564 3612 7616 3664
rect 8116 3612 8168 3664
rect 4896 3476 4948 3528
rect 5448 3519 5500 3528
rect 5448 3485 5457 3519
rect 5457 3485 5491 3519
rect 5491 3485 5500 3519
rect 5448 3476 5500 3485
rect 5632 3476 5684 3528
rect 6736 3476 6788 3528
rect 7012 3476 7064 3528
rect 7656 3544 7708 3596
rect 8208 3544 8260 3596
rect 7748 3476 7800 3528
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9036 3476 9088 3528
rect 4712 3408 4764 3460
rect 4804 3340 4856 3392
rect 4896 3340 4948 3392
rect 6828 3408 6880 3460
rect 7104 3408 7156 3460
rect 6460 3383 6512 3392
rect 6460 3349 6469 3383
rect 6469 3349 6503 3383
rect 6503 3349 6512 3383
rect 6460 3340 6512 3349
rect 7380 3340 7432 3392
rect 8576 3408 8628 3460
rect 4214 3238 4266 3290
rect 4278 3238 4330 3290
rect 4342 3238 4394 3290
rect 4406 3238 4458 3290
rect 4470 3238 4522 3290
rect 7478 3238 7530 3290
rect 7542 3238 7594 3290
rect 7606 3238 7658 3290
rect 7670 3238 7722 3290
rect 7734 3238 7786 3290
rect 4620 3136 4672 3188
rect 4712 3179 4764 3188
rect 4712 3145 4737 3179
rect 4737 3145 4764 3179
rect 4712 3136 4764 3145
rect 5356 3136 5408 3188
rect 5540 3136 5592 3188
rect 1952 3068 2004 3120
rect 3240 3000 3292 3052
rect 3608 3000 3660 3052
rect 5448 3068 5500 3120
rect 3332 2932 3384 2984
rect 4804 3000 4856 3052
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 7840 3136 7892 3188
rect 6460 3068 6512 3120
rect 8392 3136 8444 3188
rect 8484 3136 8536 3188
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 8852 3068 8904 3120
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 4988 2932 5040 2984
rect 7656 2975 7708 2984
rect 3700 2864 3752 2916
rect 3976 2864 4028 2916
rect 7656 2941 7665 2975
rect 7665 2941 7699 2975
rect 7699 2941 7708 2975
rect 7656 2932 7708 2941
rect 8484 2932 8536 2984
rect 8208 2864 8260 2916
rect 4712 2839 4764 2848
rect 4712 2805 4721 2839
rect 4721 2805 4755 2839
rect 4755 2805 4764 2839
rect 4712 2796 4764 2805
rect 5172 2796 5224 2848
rect 7012 2839 7064 2848
rect 7012 2805 7021 2839
rect 7021 2805 7055 2839
rect 7055 2805 7064 2839
rect 7012 2796 7064 2805
rect 2582 2694 2634 2746
rect 2646 2694 2698 2746
rect 2710 2694 2762 2746
rect 2774 2694 2826 2746
rect 2838 2694 2890 2746
rect 5846 2694 5898 2746
rect 5910 2694 5962 2746
rect 5974 2694 6026 2746
rect 6038 2694 6090 2746
rect 6102 2694 6154 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 9238 2694 9290 2746
rect 9302 2694 9354 2746
rect 9366 2694 9418 2746
rect 4252 2635 4304 2644
rect 4252 2601 4261 2635
rect 4261 2601 4295 2635
rect 4295 2601 4304 2635
rect 4252 2592 4304 2601
rect 4804 2592 4856 2644
rect 5080 2635 5132 2644
rect 5080 2601 5089 2635
rect 5089 2601 5123 2635
rect 5123 2601 5132 2635
rect 5080 2592 5132 2601
rect 5540 2592 5592 2644
rect 6276 2592 6328 2644
rect 6920 2592 6972 2644
rect 8668 2592 8720 2644
rect 4896 2524 4948 2576
rect 5264 2524 5316 2576
rect 8024 2524 8076 2576
rect 1860 2320 1912 2372
rect 4988 2499 5040 2508
rect 4988 2465 4997 2499
rect 4997 2465 5031 2499
rect 5031 2465 5040 2499
rect 4988 2456 5040 2465
rect 7656 2456 7708 2508
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 4252 2388 4304 2440
rect 4436 2431 4488 2440
rect 4436 2397 4445 2431
rect 4445 2397 4479 2431
rect 4479 2397 4488 2431
rect 4436 2388 4488 2397
rect 5356 2388 5408 2440
rect 7104 2388 7156 2440
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 7472 2388 7524 2440
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 6552 2320 6604 2372
rect 7012 2252 7064 2304
rect 4214 2150 4266 2202
rect 4278 2150 4330 2202
rect 4342 2150 4394 2202
rect 4406 2150 4458 2202
rect 4470 2150 4522 2202
rect 7478 2150 7530 2202
rect 7542 2150 7594 2202
rect 7606 2150 7658 2202
rect 7670 2150 7722 2202
rect 7734 2150 7786 2202
rect 2504 2048 2556 2100
rect 6644 2048 6696 2100
<< metal2 >>
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 2582 11452 2890 11472
rect 2582 11450 2588 11452
rect 2644 11450 2668 11452
rect 2724 11450 2748 11452
rect 2804 11450 2828 11452
rect 2884 11450 2890 11452
rect 2644 11398 2646 11450
rect 2826 11398 2828 11450
rect 2582 11396 2588 11398
rect 2644 11396 2668 11398
rect 2724 11396 2748 11398
rect 2804 11396 2828 11398
rect 2884 11396 2890 11398
rect 2582 11376 2890 11396
rect 5460 11354 5488 11494
rect 5846 11452 6154 11472
rect 5846 11450 5852 11452
rect 5908 11450 5932 11452
rect 5988 11450 6012 11452
rect 6068 11450 6092 11452
rect 6148 11450 6154 11452
rect 5908 11398 5910 11450
rect 6090 11398 6092 11450
rect 5846 11396 5852 11398
rect 5908 11396 5932 11398
rect 5988 11396 6012 11398
rect 6068 11396 6092 11398
rect 6148 11396 6154 11398
rect 5846 11376 6154 11396
rect 9110 11452 9418 11472
rect 9110 11450 9116 11452
rect 9172 11450 9196 11452
rect 9252 11450 9276 11452
rect 9332 11450 9356 11452
rect 9412 11450 9418 11452
rect 9172 11398 9174 11450
rect 9354 11398 9356 11450
rect 9110 11396 9116 11398
rect 9172 11396 9196 11398
rect 9252 11396 9276 11398
rect 9332 11396 9356 11398
rect 9412 11396 9418 11398
rect 9110 11376 9418 11396
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3240 11144 3292 11150
rect 3238 11112 3240 11121
rect 3792 11144 3844 11150
rect 3292 11112 3294 11121
rect 3148 11076 3200 11082
rect 3988 11121 4016 11222
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4160 11144 4212 11150
rect 3792 11086 3844 11092
rect 3974 11112 4030 11121
rect 3238 11047 3294 11056
rect 3148 11018 3200 11024
rect 1400 11008 1452 11014
rect 1400 10950 1452 10956
rect 1412 10606 1440 10950
rect 1768 10736 1820 10742
rect 1768 10678 1820 10684
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1412 10441 1440 10542
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 1688 9586 1716 10542
rect 1780 10062 1808 10678
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1766 9616 1822 9625
rect 1676 9580 1728 9586
rect 2332 9586 2360 10134
rect 2516 10062 2544 10610
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2582 10364 2890 10384
rect 2582 10362 2588 10364
rect 2644 10362 2668 10364
rect 2724 10362 2748 10364
rect 2804 10362 2828 10364
rect 2884 10362 2890 10364
rect 2644 10310 2646 10362
rect 2826 10310 2828 10362
rect 2582 10308 2588 10310
rect 2644 10308 2668 10310
rect 2724 10308 2748 10310
rect 2804 10308 2828 10310
rect 2884 10308 2890 10310
rect 2582 10288 2890 10308
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 1766 9551 1822 9560
rect 2136 9580 2188 9586
rect 1676 9522 1728 9528
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8634 1440 8910
rect 1584 8900 1636 8906
rect 1584 8842 1636 8848
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1412 7410 1440 8570
rect 1596 7954 1624 8842
rect 1688 8838 1716 9318
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1780 8566 1808 9551
rect 2136 9522 2188 9528
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 1768 8560 1820 8566
rect 1768 8502 1820 8508
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1872 7954 1900 8230
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1860 7948 1912 7954
rect 1860 7890 1912 7896
rect 1964 7478 1992 9386
rect 2148 9178 2176 9522
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2134 8936 2190 8945
rect 2056 7886 2084 8910
rect 2134 8871 2190 8880
rect 2148 8498 2176 8871
rect 2332 8498 2360 9318
rect 2424 8945 2452 9998
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2608 9722 2636 9862
rect 2596 9716 2648 9722
rect 2516 9664 2596 9674
rect 2516 9658 2648 9664
rect 2516 9646 2636 9658
rect 2516 8974 2544 9646
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2582 9276 2890 9296
rect 2582 9274 2588 9276
rect 2644 9274 2668 9276
rect 2724 9274 2748 9276
rect 2804 9274 2828 9276
rect 2884 9274 2890 9276
rect 2644 9222 2646 9274
rect 2826 9222 2828 9274
rect 2582 9220 2588 9222
rect 2644 9220 2668 9222
rect 2724 9220 2748 9222
rect 2804 9220 2828 9222
rect 2884 9220 2890 9222
rect 2582 9200 2890 9220
rect 2976 9058 3004 9522
rect 2792 9042 3004 9058
rect 2780 9036 3004 9042
rect 2832 9030 3004 9036
rect 2780 8978 2832 8984
rect 2504 8968 2556 8974
rect 2410 8936 2466 8945
rect 2504 8910 2556 8916
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2410 8871 2466 8880
rect 2516 8820 2544 8910
rect 2424 8792 2544 8820
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7546 2084 7822
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1596 3641 1624 4558
rect 1688 4282 1716 6122
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1780 4214 1808 7142
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1872 5166 1900 6938
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 1964 5846 1992 6054
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 2044 5704 2096 5710
rect 2148 5681 2176 6054
rect 2044 5646 2096 5652
rect 2134 5672 2190 5681
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1768 4208 1820 4214
rect 1768 4150 1820 4156
rect 1582 3632 1638 3641
rect 1582 3567 1638 3576
rect 1872 2378 1900 5102
rect 1964 5030 1992 5510
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1964 4146 1992 4966
rect 2056 4758 2084 5646
rect 2134 5607 2190 5616
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2044 4752 2096 4758
rect 2044 4694 2096 4700
rect 2148 4622 2176 5510
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2148 4146 2176 4422
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 1964 3126 1992 4082
rect 2240 3738 2268 6666
rect 2320 6452 2372 6458
rect 2424 6440 2452 8792
rect 2582 8188 2890 8208
rect 2582 8186 2588 8188
rect 2644 8186 2668 8188
rect 2724 8186 2748 8188
rect 2804 8186 2828 8188
rect 2884 8186 2890 8188
rect 2644 8134 2646 8186
rect 2826 8134 2828 8186
rect 2582 8132 2588 8134
rect 2644 8132 2668 8134
rect 2724 8132 2748 8134
rect 2804 8132 2828 8134
rect 2884 8132 2890 8134
rect 2582 8112 2890 8132
rect 2976 8090 3004 8910
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2582 7100 2890 7120
rect 2582 7098 2588 7100
rect 2644 7098 2668 7100
rect 2724 7098 2748 7100
rect 2804 7098 2828 7100
rect 2884 7098 2890 7100
rect 2644 7046 2646 7098
rect 2826 7046 2828 7098
rect 2582 7044 2588 7046
rect 2644 7044 2668 7046
rect 2724 7044 2748 7046
rect 2804 7044 2828 7046
rect 2884 7044 2890 7046
rect 2582 7024 2890 7044
rect 2502 6760 2558 6769
rect 2502 6695 2558 6704
rect 2372 6412 2452 6440
rect 2320 6394 2372 6400
rect 2332 5030 2360 6394
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5166 2452 6054
rect 2516 5370 2544 6695
rect 2964 6384 3016 6390
rect 3068 6372 3096 10406
rect 3160 7478 3188 11018
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3252 7954 3280 9862
rect 3344 9654 3372 10474
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3436 9518 3464 9998
rect 3528 9654 3556 10202
rect 3608 9988 3660 9994
rect 3608 9930 3660 9936
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3424 9512 3476 9518
rect 3620 9489 3648 9930
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3424 9454 3476 9460
rect 3606 9480 3662 9489
rect 3606 9415 3662 9424
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3344 7886 3372 9046
rect 3436 8634 3464 9318
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 8634 3556 8774
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3016 6344 3096 6372
rect 2964 6326 3016 6332
rect 2582 6012 2890 6032
rect 2582 6010 2588 6012
rect 2644 6010 2668 6012
rect 2724 6010 2748 6012
rect 2804 6010 2828 6012
rect 2884 6010 2890 6012
rect 2644 5958 2646 6010
rect 2826 5958 2828 6010
rect 2582 5956 2588 5958
rect 2644 5956 2668 5958
rect 2724 5956 2748 5958
rect 2804 5956 2828 5958
rect 2884 5956 2890 5958
rect 2582 5936 2890 5956
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2700 5370 2728 5646
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2412 5160 2464 5166
rect 2700 5114 2728 5306
rect 2792 5302 2820 5578
rect 2976 5574 3004 6326
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2412 5102 2464 5108
rect 2516 5086 2728 5114
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2516 4826 2544 5086
rect 2582 4924 2890 4944
rect 2582 4922 2588 4924
rect 2644 4922 2668 4924
rect 2724 4922 2748 4924
rect 2804 4922 2828 4924
rect 2884 4922 2890 4924
rect 2644 4870 2646 4922
rect 2826 4870 2828 4922
rect 2582 4868 2588 4870
rect 2644 4868 2668 4870
rect 2724 4868 2748 4870
rect 2804 4868 2828 4870
rect 2884 4868 2890 4870
rect 2582 4848 2890 4868
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2976 4214 3004 5510
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2596 4208 2648 4214
rect 2594 4176 2596 4185
rect 2964 4208 3016 4214
rect 2648 4176 2650 4185
rect 2964 4150 3016 4156
rect 2594 4111 2650 4120
rect 2962 4040 3018 4049
rect 2962 3975 3018 3984
rect 2976 3942 3004 3975
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2582 3836 2890 3856
rect 2582 3834 2588 3836
rect 2644 3834 2668 3836
rect 2724 3834 2748 3836
rect 2804 3834 2828 3836
rect 2884 3834 2890 3836
rect 2644 3782 2646 3834
rect 2826 3782 2828 3834
rect 2582 3780 2588 3782
rect 2644 3780 2668 3782
rect 2724 3780 2748 3782
rect 2804 3780 2828 3782
rect 2884 3780 2890 3782
rect 2582 3760 2890 3780
rect 2962 3768 3018 3777
rect 2228 3732 2280 3738
rect 2962 3703 2964 3712
rect 2228 3674 2280 3680
rect 3016 3703 3018 3712
rect 2964 3674 3016 3680
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 2582 2748 2890 2768
rect 2582 2746 2588 2748
rect 2644 2746 2668 2748
rect 2724 2746 2748 2748
rect 2804 2746 2828 2748
rect 2884 2746 2890 2748
rect 2644 2694 2646 2746
rect 2826 2694 2828 2746
rect 2582 2692 2588 2694
rect 2644 2692 2668 2694
rect 2724 2692 2748 2694
rect 2804 2692 2828 2694
rect 2884 2692 2890 2694
rect 2582 2672 2890 2692
rect 3068 2446 3096 4422
rect 3160 4010 3188 6598
rect 3344 5642 3372 6598
rect 3620 5914 3648 9318
rect 3712 6662 3740 9522
rect 3804 9178 3832 11086
rect 3974 11047 4030 11056
rect 4080 11092 4160 11098
rect 4080 11086 4212 11092
rect 4540 11098 4568 11154
rect 4080 11070 4200 11086
rect 4540 11070 4660 11098
rect 4080 10690 4108 11070
rect 4214 10908 4522 10928
rect 4214 10906 4220 10908
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4516 10906 4522 10908
rect 4276 10854 4278 10906
rect 4458 10854 4460 10906
rect 4214 10852 4220 10854
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4516 10852 4522 10854
rect 4214 10832 4522 10852
rect 4080 10662 4200 10690
rect 3976 10600 4028 10606
rect 3974 10568 3976 10577
rect 4028 10568 4030 10577
rect 3974 10503 4030 10512
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3974 10296 4030 10305
rect 3974 10231 4030 10240
rect 3988 9586 4016 10231
rect 4080 10130 4108 10406
rect 4172 10130 4200 10662
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4250 10568 4306 10577
rect 4250 10503 4306 10512
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4264 10010 4292 10503
rect 4080 9982 4292 10010
rect 4448 9994 4476 10610
rect 4436 9988 4488 9994
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 4080 8922 4108 9982
rect 4540 9976 4568 10610
rect 4632 10470 4660 11070
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 10044 4660 10406
rect 4632 10016 4752 10044
rect 4540 9948 4660 9976
rect 4436 9930 4488 9936
rect 4214 9820 4522 9840
rect 4214 9818 4220 9820
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4516 9818 4522 9820
rect 4276 9766 4278 9818
rect 4458 9766 4460 9818
rect 4214 9764 4220 9766
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4516 9764 4522 9766
rect 4214 9744 4522 9764
rect 4632 9761 4660 9948
rect 4618 9752 4674 9761
rect 4618 9687 4674 9696
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 3988 8894 4108 8922
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3804 8242 3832 8366
rect 3988 8344 4016 8894
rect 4068 8832 4120 8838
rect 4172 8820 4200 9522
rect 4540 9489 4568 9522
rect 4526 9480 4582 9489
rect 4526 9415 4582 9424
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4264 8945 4292 9114
rect 4632 9110 4660 9687
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4250 8936 4306 8945
rect 4724 8922 4752 10016
rect 4816 9625 4844 11290
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10674 4936 10950
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4908 10441 4936 10474
rect 4894 10432 4950 10441
rect 4894 10367 4950 10376
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4802 9616 4858 9625
rect 4802 9551 4858 9560
rect 4250 8871 4306 8880
rect 4620 8900 4672 8906
rect 4724 8894 4844 8922
rect 4620 8842 4672 8848
rect 4068 8774 4120 8780
rect 4152 8792 4200 8820
rect 4080 8514 4108 8774
rect 4152 8616 4180 8792
rect 4214 8732 4522 8752
rect 4214 8730 4220 8732
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4516 8730 4522 8732
rect 4276 8678 4278 8730
rect 4458 8678 4460 8730
rect 4214 8676 4220 8678
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4516 8676 4522 8678
rect 4214 8656 4522 8676
rect 4152 8588 4292 8616
rect 4080 8486 4200 8514
rect 3988 8316 4108 8344
rect 3804 8214 4016 8242
rect 3988 6798 4016 8214
rect 4080 7002 4108 8316
rect 4172 8294 4200 8486
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4172 8090 4200 8230
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4264 7732 4292 8588
rect 4632 7818 4660 8842
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4724 8498 4752 8570
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4152 7704 4292 7732
rect 4152 7528 4180 7704
rect 4214 7644 4522 7664
rect 4214 7642 4220 7644
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4516 7642 4522 7644
rect 4276 7590 4278 7642
rect 4458 7590 4460 7642
rect 4214 7588 4220 7590
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4516 7588 4522 7590
rect 4214 7568 4522 7588
rect 4152 7500 4200 7528
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4172 6934 4200 7500
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 3976 6792 4028 6798
rect 4172 6769 4200 6870
rect 3976 6734 4028 6740
rect 4158 6760 4214 6769
rect 3884 6724 3936 6730
rect 3884 6666 3936 6672
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3160 3738 3188 3946
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3252 3058 3280 5510
rect 3436 5234 3464 5714
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3344 3602 3372 5102
rect 3436 4826 3464 5170
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3528 4758 3556 5102
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3344 2990 3372 3538
rect 3436 3097 3464 4218
rect 3422 3088 3478 3097
rect 3620 3058 3648 5034
rect 3422 3023 3478 3032
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3712 2922 3740 6258
rect 3896 5574 3924 6666
rect 3988 6118 4016 6734
rect 4158 6695 4214 6704
rect 4214 6556 4522 6576
rect 4214 6554 4220 6556
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4516 6554 4522 6556
rect 4276 6502 4278 6554
rect 4458 6502 4460 6554
rect 4214 6500 4220 6502
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4516 6500 4522 6502
rect 4214 6480 4522 6500
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3804 3942 3832 4966
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3896 3534 3924 5510
rect 4080 4622 4108 5578
rect 4724 5545 4752 6054
rect 4710 5536 4766 5545
rect 4214 5468 4522 5488
rect 4710 5471 4766 5480
rect 4214 5466 4220 5468
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4516 5466 4522 5468
rect 4276 5414 4278 5466
rect 4458 5414 4460 5466
rect 4214 5412 4220 5414
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4516 5412 4522 5414
rect 4214 5392 4522 5412
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4264 4690 4292 5238
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4214 4380 4522 4400
rect 4214 4378 4220 4380
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4516 4378 4522 4380
rect 4276 4326 4278 4378
rect 4458 4326 4460 4378
rect 4214 4324 4220 4326
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4516 4324 4522 4326
rect 4214 4304 4522 4324
rect 4252 4208 4304 4214
rect 4632 4162 4660 4490
rect 4252 4150 4304 4156
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3988 2922 4016 3946
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3505 4108 3878
rect 4264 3505 4292 4150
rect 4540 4146 4660 4162
rect 4528 4140 4660 4146
rect 4580 4134 4660 4140
rect 4528 4082 4580 4088
rect 4724 3618 4752 5170
rect 4816 4049 4844 8894
rect 4908 8838 4936 10066
rect 5000 9761 5028 11086
rect 5080 10736 5132 10742
rect 5080 10678 5132 10684
rect 4986 9752 5042 9761
rect 5092 9722 5120 10678
rect 4986 9687 5042 9696
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 5000 9042 5028 9590
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8634 4936 8774
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5000 8566 5028 8978
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4908 4593 4936 8434
rect 5000 7818 5028 8502
rect 5092 8090 5120 8910
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 5000 7478 5028 7754
rect 5092 7546 5120 8026
rect 5184 7818 5212 11222
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 5264 11008 5316 11014
rect 5262 10976 5264 10985
rect 5316 10976 5318 10985
rect 5262 10911 5318 10920
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5276 10305 5304 10474
rect 5262 10296 5318 10305
rect 5262 10231 5318 10240
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5276 9654 5304 9998
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 5368 9466 5396 11086
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6368 10736 6420 10742
rect 6368 10678 6420 10684
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5276 9438 5396 9466
rect 5276 8498 5304 9438
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5368 8401 5396 8842
rect 5354 8392 5410 8401
rect 5354 8327 5410 8336
rect 5460 8294 5488 10202
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 5000 7002 5028 7414
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5000 6322 5028 6938
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5000 5302 5028 6258
rect 5262 6216 5318 6225
rect 5262 6151 5318 6160
rect 5078 5808 5134 5817
rect 5078 5743 5134 5752
rect 4988 5296 5040 5302
rect 4988 5238 5040 5244
rect 4894 4584 4950 4593
rect 4894 4519 4950 4528
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4802 4040 4858 4049
rect 4908 4026 4936 4422
rect 5000 4214 5028 5238
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 4908 3998 5028 4026
rect 4802 3975 4858 3984
rect 4894 3768 4950 3777
rect 4894 3703 4950 3712
rect 4632 3590 4752 3618
rect 4066 3496 4122 3505
rect 4066 3431 4122 3440
rect 4250 3496 4306 3505
rect 4250 3431 4306 3440
rect 4214 3292 4522 3312
rect 4214 3290 4220 3292
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4516 3290 4522 3292
rect 4276 3238 4278 3290
rect 4458 3238 4460 3290
rect 4214 3236 4220 3238
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4516 3236 4522 3238
rect 4214 3216 4522 3236
rect 4632 3194 4660 3590
rect 4908 3534 4936 3703
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4724 3194 4752 3402
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4816 3058 4844 3334
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 3700 2916 3752 2922
rect 3700 2858 3752 2864
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 4356 2910 4752 2938
rect 4250 2680 4306 2689
rect 4250 2615 4252 2624
rect 4304 2615 4306 2624
rect 4252 2586 4304 2592
rect 4356 2530 4384 2910
rect 4724 2854 4752 2910
rect 4712 2848 4764 2854
rect 4434 2816 4490 2825
rect 4712 2790 4764 2796
rect 4434 2751 4490 2760
rect 4264 2502 4384 2530
rect 4264 2446 4292 2502
rect 4448 2446 4476 2751
rect 4816 2650 4844 2994
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4908 2582 4936 3334
rect 5000 2990 5028 3998
rect 5092 3777 5120 5743
rect 5276 5710 5304 6151
rect 5552 5710 5580 10406
rect 5846 10364 6154 10384
rect 5846 10362 5852 10364
rect 5908 10362 5932 10364
rect 5988 10362 6012 10364
rect 6068 10362 6092 10364
rect 6148 10362 6154 10364
rect 5908 10310 5910 10362
rect 6090 10310 6092 10362
rect 5846 10308 5852 10310
rect 5908 10308 5932 10310
rect 5988 10308 6012 10310
rect 6068 10308 6092 10310
rect 6148 10308 6154 10310
rect 5846 10288 6154 10308
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6196 9382 6224 9862
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 5846 9276 6154 9296
rect 5846 9274 5852 9276
rect 5908 9274 5932 9276
rect 5988 9274 6012 9276
rect 6068 9274 6092 9276
rect 6148 9274 6154 9276
rect 5908 9222 5910 9274
rect 6090 9222 6092 9274
rect 5846 9220 5852 9222
rect 5908 9220 5932 9222
rect 5988 9220 6012 9222
rect 6068 9220 6092 9222
rect 6148 9220 6154 9222
rect 5846 9200 6154 9220
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5644 6866 5672 9114
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5736 6730 5764 8298
rect 5846 8188 6154 8208
rect 5846 8186 5852 8188
rect 5908 8186 5932 8188
rect 5988 8186 6012 8188
rect 6068 8186 6092 8188
rect 6148 8186 6154 8188
rect 5908 8134 5910 8186
rect 6090 8134 6092 8186
rect 5846 8132 5852 8134
rect 5908 8132 5932 8134
rect 5988 8132 6012 8134
rect 6068 8132 6092 8134
rect 6148 8132 6154 8134
rect 5846 8112 6154 8132
rect 5846 7100 6154 7120
rect 5846 7098 5852 7100
rect 5908 7098 5932 7100
rect 5988 7098 6012 7100
rect 6068 7098 6092 7100
rect 6148 7098 6154 7100
rect 5908 7046 5910 7098
rect 6090 7046 6092 7098
rect 5846 7044 5852 7046
rect 5908 7044 5932 7046
rect 5988 7044 6012 7046
rect 6068 7044 6092 7046
rect 6148 7044 6154 7046
rect 5846 7024 6154 7044
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5276 5370 5304 5646
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5368 5302 5396 5510
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5262 5128 5318 5137
rect 5262 5063 5318 5072
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5078 3768 5134 3777
rect 5078 3703 5134 3712
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5000 2514 5028 2926
rect 5092 2650 5120 3606
rect 5184 2854 5212 4966
rect 5276 4185 5304 5063
rect 5262 4176 5318 4185
rect 5262 4111 5318 4120
rect 5276 2961 5304 4111
rect 5368 3670 5396 5238
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5460 3534 5488 4762
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5552 4282 5580 4558
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5540 3732 5592 3738
rect 5644 3720 5672 5238
rect 5736 3942 5764 6666
rect 5846 6012 6154 6032
rect 5846 6010 5852 6012
rect 5908 6010 5932 6012
rect 5988 6010 6012 6012
rect 6068 6010 6092 6012
rect 6148 6010 6154 6012
rect 5908 5958 5910 6010
rect 6090 5958 6092 6010
rect 5846 5956 5852 5958
rect 5908 5956 5932 5958
rect 5988 5956 6012 5958
rect 6068 5956 6092 5958
rect 6148 5956 6154 5958
rect 5846 5936 6154 5956
rect 6196 5370 6224 9318
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 5846 4924 6154 4944
rect 5846 4922 5852 4924
rect 5908 4922 5932 4924
rect 5988 4922 6012 4924
rect 6068 4922 6092 4924
rect 6148 4922 6154 4924
rect 5908 4870 5910 4922
rect 6090 4870 6092 4922
rect 5846 4868 5852 4870
rect 5908 4868 5932 4870
rect 5988 4868 6012 4870
rect 6068 4868 6092 4870
rect 6148 4868 6154 4870
rect 5846 4848 6154 4868
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5846 3836 6154 3856
rect 5846 3834 5852 3836
rect 5908 3834 5932 3836
rect 5988 3834 6012 3836
rect 6068 3834 6092 3836
rect 6148 3834 6154 3836
rect 5908 3782 5910 3834
rect 6090 3782 6092 3834
rect 5846 3780 5852 3782
rect 5908 3780 5932 3782
rect 5988 3780 6012 3782
rect 6068 3780 6092 3782
rect 6148 3780 6154 3782
rect 5846 3760 6154 3780
rect 5592 3692 5672 3720
rect 5540 3674 5592 3680
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5262 2952 5318 2961
rect 5262 2887 5318 2896
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5262 2816 5318 2825
rect 5262 2751 5318 2760
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5276 2582 5304 2751
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 5368 2446 5396 3130
rect 5460 3126 5488 3470
rect 5552 3194 5580 3674
rect 6288 3602 6316 10406
rect 6380 9738 6408 10678
rect 6564 10674 6592 10950
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6380 9722 6500 9738
rect 6380 9716 6512 9722
rect 6380 9710 6460 9716
rect 6380 8634 6408 9710
rect 6460 9658 6512 9664
rect 6564 9586 6592 10610
rect 6748 10198 6776 11086
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6380 6390 6408 7278
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 6380 5778 6408 6326
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6380 5234 6408 5714
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6380 4690 6408 5170
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6380 3777 6408 4082
rect 6366 3768 6422 3777
rect 6472 3738 6500 9318
rect 6840 9110 6868 11154
rect 7478 10908 7786 10928
rect 7478 10906 7484 10908
rect 7540 10906 7564 10908
rect 7620 10906 7644 10908
rect 7700 10906 7724 10908
rect 7780 10906 7786 10908
rect 7540 10854 7542 10906
rect 7722 10854 7724 10906
rect 7478 10852 7484 10854
rect 7540 10852 7564 10854
rect 7620 10852 7644 10854
rect 7700 10852 7724 10854
rect 7780 10852 7786 10854
rect 7478 10832 7786 10852
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7562 10568 7618 10577
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6932 9625 6960 10474
rect 7116 10130 7144 10542
rect 7562 10503 7618 10512
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 7024 9761 7052 9998
rect 7010 9752 7066 9761
rect 7010 9687 7066 9696
rect 6918 9616 6974 9625
rect 6918 9551 6974 9560
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 7024 8945 7052 9687
rect 7116 9654 7144 10066
rect 7484 10062 7512 10406
rect 7576 10062 7604 10503
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7478 9820 7786 9840
rect 7478 9818 7484 9820
rect 7540 9818 7564 9820
rect 7620 9818 7644 9820
rect 7700 9818 7724 9820
rect 7780 9818 7786 9820
rect 7540 9766 7542 9818
rect 7722 9766 7724 9818
rect 7478 9764 7484 9766
rect 7540 9764 7564 9766
rect 7620 9764 7644 9766
rect 7700 9764 7724 9766
rect 7780 9764 7786 9766
rect 7478 9744 7786 9764
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7010 8936 7066 8945
rect 7010 8871 7066 8880
rect 7024 8129 7052 8871
rect 7010 8120 7066 8129
rect 7010 8055 7066 8064
rect 7010 7984 7066 7993
rect 7010 7919 7066 7928
rect 7024 7886 7052 7919
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7116 7698 7144 9590
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7760 8906 7788 9454
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7024 7670 7144 7698
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6366 3703 6422 3712
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5538 3088 5594 3097
rect 5644 3040 5672 3470
rect 5594 3032 5672 3040
rect 5538 3023 5540 3032
rect 5592 3012 5672 3032
rect 5540 2994 5592 3000
rect 5552 2650 5580 2994
rect 5846 2748 6154 2768
rect 5846 2746 5852 2748
rect 5908 2746 5932 2748
rect 5988 2746 6012 2748
rect 6068 2746 6092 2748
rect 6148 2746 6154 2748
rect 5908 2694 5910 2746
rect 6090 2694 6092 2746
rect 5846 2692 5852 2694
rect 5908 2692 5932 2694
rect 5988 2692 6012 2694
rect 6068 2692 6092 2694
rect 6148 2692 6154 2694
rect 5846 2672 6154 2692
rect 6288 2650 6316 3538
rect 6458 3496 6514 3505
rect 6458 3431 6514 3440
rect 6472 3398 6500 3431
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 3126 6500 3334
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 6564 2378 6592 6258
rect 6644 5568 6696 5574
rect 6642 5536 6644 5545
rect 6696 5536 6698 5545
rect 6642 5471 6698 5480
rect 6644 5228 6696 5234
rect 6920 5228 6972 5234
rect 6644 5170 6696 5176
rect 6748 5188 6920 5216
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 2106 2544 2246
rect 4214 2204 4522 2224
rect 4214 2202 4220 2204
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4516 2202 4522 2204
rect 4276 2150 4278 2202
rect 4458 2150 4460 2202
rect 4214 2148 4220 2150
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4516 2148 4522 2150
rect 4214 2128 4522 2148
rect 6656 2106 6684 5170
rect 6748 3534 6776 5188
rect 6920 5170 6972 5176
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6840 3466 6868 4218
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6932 2650 6960 4490
rect 7024 3618 7052 7670
rect 7102 5672 7158 5681
rect 7102 5607 7158 5616
rect 7116 4554 7144 5607
rect 7208 5234 7236 7686
rect 7300 5273 7328 8774
rect 7478 8732 7786 8752
rect 7478 8730 7484 8732
rect 7540 8730 7564 8732
rect 7620 8730 7644 8732
rect 7700 8730 7724 8732
rect 7780 8730 7786 8732
rect 7540 8678 7542 8730
rect 7722 8678 7724 8730
rect 7478 8676 7484 8678
rect 7540 8676 7564 8678
rect 7620 8676 7644 8678
rect 7700 8676 7724 8678
rect 7780 8676 7786 8678
rect 7478 8656 7786 8676
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7760 7954 7788 8434
rect 7852 8362 7880 10066
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7478 7644 7786 7664
rect 7478 7642 7484 7644
rect 7540 7642 7564 7644
rect 7620 7642 7644 7644
rect 7700 7642 7724 7644
rect 7780 7642 7786 7644
rect 7540 7590 7542 7642
rect 7722 7590 7724 7642
rect 7478 7588 7484 7590
rect 7540 7588 7564 7590
rect 7620 7588 7644 7590
rect 7700 7588 7724 7590
rect 7780 7588 7786 7590
rect 7478 7568 7786 7588
rect 7852 7478 7880 7686
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7286 5264 7342 5273
rect 7196 5228 7248 5234
rect 7286 5199 7342 5208
rect 7196 5170 7248 5176
rect 7392 4758 7420 7346
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7478 6556 7786 6576
rect 7478 6554 7484 6556
rect 7540 6554 7564 6556
rect 7620 6554 7644 6556
rect 7700 6554 7724 6556
rect 7780 6554 7786 6556
rect 7540 6502 7542 6554
rect 7722 6502 7724 6554
rect 7478 6500 7484 6502
rect 7540 6500 7564 6502
rect 7620 6500 7644 6502
rect 7700 6500 7724 6502
rect 7780 6500 7786 6502
rect 7478 6480 7786 6500
rect 7852 6118 7880 6734
rect 7944 6497 7972 10202
rect 7930 6488 7986 6497
rect 7930 6423 7986 6432
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5710 7880 6054
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7478 5468 7786 5488
rect 7478 5466 7484 5468
rect 7540 5466 7564 5468
rect 7620 5466 7644 5468
rect 7700 5466 7724 5468
rect 7780 5466 7786 5468
rect 7540 5414 7542 5466
rect 7722 5414 7724 5466
rect 7478 5412 7484 5414
rect 7540 5412 7564 5414
rect 7620 5412 7644 5414
rect 7700 5412 7724 5414
rect 7780 5412 7786 5414
rect 7478 5392 7786 5412
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7852 5166 7880 5306
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 7576 4554 7604 4966
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7380 4548 7432 4554
rect 7380 4490 7432 4496
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7102 4040 7158 4049
rect 7102 3975 7158 3984
rect 7116 3738 7144 3975
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7208 3670 7236 4422
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7300 3738 7328 3878
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7196 3664 7248 3670
rect 7024 3590 7144 3618
rect 7392 3618 7420 4490
rect 7478 4380 7786 4400
rect 7478 4378 7484 4380
rect 7540 4378 7564 4380
rect 7620 4378 7644 4380
rect 7700 4378 7724 4380
rect 7780 4378 7786 4380
rect 7540 4326 7542 4378
rect 7722 4326 7724 4378
rect 7478 4324 7484 4326
rect 7540 4324 7564 4326
rect 7620 4324 7644 4326
rect 7700 4324 7724 4326
rect 7780 4324 7786 4326
rect 7478 4304 7786 4324
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7196 3606 7248 3612
rect 7012 3528 7064 3534
rect 7010 3496 7012 3505
rect 7064 3496 7066 3505
rect 7116 3466 7144 3590
rect 7010 3431 7066 3440
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7024 2310 7052 2790
rect 7116 2446 7144 3402
rect 7208 3058 7236 3606
rect 7300 3590 7420 3618
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7300 2446 7328 3590
rect 7576 3482 7604 3606
rect 7668 3602 7696 3946
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7748 3528 7800 3534
rect 7576 3476 7748 3482
rect 7576 3470 7800 3476
rect 7576 3454 7788 3470
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 2774 7420 3334
rect 7478 3292 7786 3312
rect 7478 3290 7484 3292
rect 7540 3290 7564 3292
rect 7620 3290 7644 3292
rect 7700 3290 7724 3292
rect 7780 3290 7786 3292
rect 7540 3238 7542 3290
rect 7722 3238 7724 3290
rect 7478 3236 7484 3238
rect 7540 3236 7564 3238
rect 7620 3236 7644 3238
rect 7700 3236 7724 3238
rect 7780 3236 7786 3238
rect 7478 3216 7786 3236
rect 7852 3194 7880 4490
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7392 2746 7512 2774
rect 7484 2446 7512 2746
rect 7668 2514 7696 2926
rect 8036 2582 8064 10610
rect 8128 9489 8156 11290
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8220 10810 8248 11086
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8220 10130 8248 10746
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8312 9654 8340 10406
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 9648 8352 9654
rect 8206 9616 8262 9625
rect 8300 9590 8352 9596
rect 8206 9551 8262 9560
rect 8114 9480 8170 9489
rect 8114 9415 8170 9424
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8128 8566 8156 8910
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8220 7546 8248 9551
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8312 8974 8340 9454
rect 8404 9042 8432 9862
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8496 8838 8524 11018
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 8680 10266 8708 10678
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9722 8616 9998
rect 8680 9722 8708 10202
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8588 9586 8616 9658
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8680 9330 8708 9658
rect 8772 9586 8800 11154
rect 9140 10674 9168 11222
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8680 9302 8800 9330
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8312 7018 8340 7414
rect 8220 6990 8340 7018
rect 8114 6760 8170 6769
rect 8114 6695 8170 6704
rect 8128 3670 8156 6695
rect 8220 5846 8248 6990
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8312 6322 8340 6870
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8312 5778 8340 6258
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8404 5658 8432 8298
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 8022 8524 8230
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8312 5630 8432 5658
rect 8496 5642 8524 7686
rect 8680 7562 8708 9114
rect 8588 7534 8708 7562
rect 8588 6118 8616 7534
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8484 5636 8536 5642
rect 8220 4826 8248 5578
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8220 2922 8248 3538
rect 8312 3534 8340 5630
rect 8484 5578 8536 5584
rect 8588 5522 8616 5782
rect 8496 5494 8616 5522
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8404 5137 8432 5170
rect 8390 5128 8446 5137
rect 8390 5063 8446 5072
rect 8392 4820 8444 4826
rect 8496 4808 8524 5494
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 8444 4780 8524 4808
rect 8392 4762 8444 4768
rect 8404 4282 8432 4762
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8496 3194 8524 4626
rect 8588 3466 8616 5034
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8404 3058 8432 3130
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8496 2990 8524 3130
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 8680 2650 8708 7414
rect 8772 5370 8800 9302
rect 8864 9110 8892 9590
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 8956 8906 8984 10406
rect 9110 10364 9418 10384
rect 9110 10362 9116 10364
rect 9172 10362 9196 10364
rect 9252 10362 9276 10364
rect 9332 10362 9356 10364
rect 9412 10362 9418 10364
rect 9172 10310 9174 10362
rect 9354 10310 9356 10362
rect 9110 10308 9116 10310
rect 9172 10308 9196 10310
rect 9252 10308 9276 10310
rect 9332 10308 9356 10310
rect 9412 10308 9418 10310
rect 9110 10288 9418 10308
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 9048 8634 9076 9862
rect 9232 9654 9260 9998
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9220 9648 9272 9654
rect 9126 9616 9182 9625
rect 9220 9590 9272 9596
rect 9126 9551 9182 9560
rect 9140 9518 9168 9551
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9494 9480 9550 9489
rect 9494 9415 9496 9424
rect 9548 9415 9550 9424
rect 9496 9386 9548 9392
rect 9110 9276 9418 9296
rect 9110 9274 9116 9276
rect 9172 9274 9196 9276
rect 9252 9274 9276 9276
rect 9332 9274 9356 9276
rect 9412 9274 9418 9276
rect 9172 9222 9174 9274
rect 9354 9222 9356 9274
rect 9110 9220 9116 9222
rect 9172 9220 9196 9222
rect 9252 9220 9276 9222
rect 9332 9220 9356 9222
rect 9412 9220 9418 9222
rect 9110 9200 9418 9220
rect 9600 9042 9628 9862
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 10152 8974 10180 11494
rect 9496 8968 9548 8974
rect 9494 8936 9496 8945
rect 10140 8968 10192 8974
rect 9548 8936 9550 8945
rect 10140 8910 10192 8916
rect 9494 8871 9550 8880
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9110 8188 9418 8208
rect 9110 8186 9116 8188
rect 9172 8186 9196 8188
rect 9252 8186 9276 8188
rect 9332 8186 9356 8188
rect 9412 8186 9418 8188
rect 9172 8134 9174 8186
rect 9354 8134 9356 8186
rect 9110 8132 9116 8134
rect 9172 8132 9196 8134
rect 9252 8132 9276 8134
rect 9332 8132 9356 8134
rect 9412 8132 9418 8134
rect 9110 8112 9418 8132
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8864 5370 8892 7754
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8758 5264 8814 5273
rect 8758 5199 8814 5208
rect 8772 4146 8800 5199
rect 8864 4486 8892 5306
rect 8956 5234 8984 7142
rect 9048 5692 9076 7822
rect 9110 7100 9418 7120
rect 9110 7098 9116 7100
rect 9172 7098 9196 7100
rect 9252 7098 9276 7100
rect 9332 7098 9356 7100
rect 9412 7098 9418 7100
rect 9172 7046 9174 7098
rect 9354 7046 9356 7098
rect 9110 7044 9116 7046
rect 9172 7044 9196 7046
rect 9252 7044 9276 7046
rect 9332 7044 9356 7046
rect 9412 7044 9418 7046
rect 9110 7024 9418 7044
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9324 6769 9352 6802
rect 9404 6792 9456 6798
rect 9310 6760 9366 6769
rect 9404 6734 9456 6740
rect 9508 6746 9536 8434
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9600 7410 9628 8366
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9600 6934 9628 7346
rect 10046 7032 10102 7041
rect 10046 6967 10102 6976
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9678 6896 9734 6905
rect 9678 6831 9734 6840
rect 9310 6695 9366 6704
rect 9128 6656 9180 6662
rect 9312 6656 9364 6662
rect 9128 6598 9180 6604
rect 9310 6624 9312 6633
rect 9364 6624 9366 6633
rect 9140 6225 9168 6598
rect 9310 6559 9366 6568
rect 9416 6497 9444 6734
rect 9508 6718 9628 6746
rect 9600 6662 9628 6718
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9402 6488 9458 6497
rect 9402 6423 9458 6432
rect 9126 6216 9182 6225
rect 9126 6151 9182 6160
rect 9110 6012 9418 6032
rect 9110 6010 9116 6012
rect 9172 6010 9196 6012
rect 9252 6010 9276 6012
rect 9332 6010 9356 6012
rect 9412 6010 9418 6012
rect 9172 5958 9174 6010
rect 9354 5958 9356 6010
rect 9110 5956 9116 5958
rect 9172 5956 9196 5958
rect 9252 5956 9276 5958
rect 9332 5956 9356 5958
rect 9412 5956 9418 5958
rect 9110 5936 9418 5956
rect 9508 5817 9536 6598
rect 9600 6390 9628 6598
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9692 5914 9720 6831
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9494 5808 9550 5817
rect 9404 5772 9456 5778
rect 9494 5743 9550 5752
rect 9404 5714 9456 5720
rect 9128 5704 9180 5710
rect 9048 5664 9128 5692
rect 9128 5646 9180 5652
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8956 4570 8984 5170
rect 9140 5098 9168 5646
rect 9416 5370 9444 5714
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9110 4924 9418 4944
rect 9110 4922 9116 4924
rect 9172 4922 9196 4924
rect 9252 4922 9276 4924
rect 9332 4922 9356 4924
rect 9412 4922 9418 4924
rect 9172 4870 9174 4922
rect 9354 4870 9356 4922
rect 9110 4868 9116 4870
rect 9172 4868 9196 4870
rect 9252 4868 9276 4870
rect 9332 4868 9356 4870
rect 9412 4868 9418 4870
rect 9110 4848 9418 4868
rect 9508 4808 9536 5646
rect 9586 5264 9642 5273
rect 9586 5199 9588 5208
rect 9640 5199 9642 5208
rect 9588 5170 9640 5176
rect 9324 4780 9536 4808
rect 9324 4622 9352 4780
rect 9312 4616 9364 4622
rect 8956 4542 9168 4570
rect 9312 4558 9364 4564
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8956 4282 8984 4542
rect 9140 4486 9168 4542
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 8944 4276 8996 4282
rect 8864 4236 8944 4264
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8758 3768 8814 3777
rect 8758 3703 8760 3712
rect 8812 3703 8814 3712
rect 8760 3674 8812 3680
rect 8864 3126 8892 4236
rect 8944 4218 8996 4224
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8956 3534 8984 4082
rect 9048 3534 9076 4422
rect 9324 4078 9352 4558
rect 9416 4146 9444 4558
rect 9876 4146 9904 6054
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 10060 4010 10088 6967
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10152 5710 10180 6394
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9110 3836 9418 3856
rect 9110 3834 9116 3836
rect 9172 3834 9196 3836
rect 9252 3834 9276 3836
rect 9332 3834 9356 3836
rect 9412 3834 9418 3836
rect 9172 3782 9174 3834
rect 9354 3782 9356 3834
rect 9110 3780 9116 3782
rect 9172 3780 9196 3782
rect 9252 3780 9276 3782
rect 9332 3780 9356 3782
rect 9412 3780 9418 3782
rect 9110 3760 9418 3780
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 9110 2748 9418 2768
rect 9110 2746 9116 2748
rect 9172 2746 9196 2748
rect 9252 2746 9276 2748
rect 9332 2746 9356 2748
rect 9412 2746 9418 2748
rect 9172 2694 9174 2746
rect 9354 2694 9356 2746
rect 9110 2692 9116 2694
rect 9172 2692 9196 2694
rect 9252 2692 9276 2694
rect 9332 2692 9356 2694
rect 9412 2692 9418 2694
rect 9110 2672 9418 2692
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7478 2204 7786 2224
rect 7478 2202 7484 2204
rect 7540 2202 7564 2204
rect 7620 2202 7644 2204
rect 7700 2202 7724 2204
rect 7780 2202 7786 2204
rect 7540 2150 7542 2202
rect 7722 2150 7724 2202
rect 7478 2148 7484 2150
rect 7540 2148 7564 2150
rect 7620 2148 7644 2150
rect 7700 2148 7724 2150
rect 7780 2148 7786 2150
rect 7478 2128 7786 2148
rect 2504 2100 2556 2106
rect 2504 2042 2556 2048
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
<< via2 >>
rect 2588 11450 2644 11452
rect 2668 11450 2724 11452
rect 2748 11450 2804 11452
rect 2828 11450 2884 11452
rect 2588 11398 2634 11450
rect 2634 11398 2644 11450
rect 2668 11398 2698 11450
rect 2698 11398 2710 11450
rect 2710 11398 2724 11450
rect 2748 11398 2762 11450
rect 2762 11398 2774 11450
rect 2774 11398 2804 11450
rect 2828 11398 2838 11450
rect 2838 11398 2884 11450
rect 2588 11396 2644 11398
rect 2668 11396 2724 11398
rect 2748 11396 2804 11398
rect 2828 11396 2884 11398
rect 5852 11450 5908 11452
rect 5932 11450 5988 11452
rect 6012 11450 6068 11452
rect 6092 11450 6148 11452
rect 5852 11398 5898 11450
rect 5898 11398 5908 11450
rect 5932 11398 5962 11450
rect 5962 11398 5974 11450
rect 5974 11398 5988 11450
rect 6012 11398 6026 11450
rect 6026 11398 6038 11450
rect 6038 11398 6068 11450
rect 6092 11398 6102 11450
rect 6102 11398 6148 11450
rect 5852 11396 5908 11398
rect 5932 11396 5988 11398
rect 6012 11396 6068 11398
rect 6092 11396 6148 11398
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 9276 11450 9332 11452
rect 9356 11450 9412 11452
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9238 11450
rect 9238 11398 9252 11450
rect 9276 11398 9290 11450
rect 9290 11398 9302 11450
rect 9302 11398 9332 11450
rect 9356 11398 9366 11450
rect 9366 11398 9412 11450
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 9276 11396 9332 11398
rect 9356 11396 9412 11398
rect 3238 11092 3240 11112
rect 3240 11092 3292 11112
rect 3292 11092 3294 11112
rect 3238 11056 3294 11092
rect 1398 10376 1454 10432
rect 1766 9560 1822 9616
rect 2588 10362 2644 10364
rect 2668 10362 2724 10364
rect 2748 10362 2804 10364
rect 2828 10362 2884 10364
rect 2588 10310 2634 10362
rect 2634 10310 2644 10362
rect 2668 10310 2698 10362
rect 2698 10310 2710 10362
rect 2710 10310 2724 10362
rect 2748 10310 2762 10362
rect 2762 10310 2774 10362
rect 2774 10310 2804 10362
rect 2828 10310 2838 10362
rect 2838 10310 2884 10362
rect 2588 10308 2644 10310
rect 2668 10308 2724 10310
rect 2748 10308 2804 10310
rect 2828 10308 2884 10310
rect 2134 8880 2190 8936
rect 2588 9274 2644 9276
rect 2668 9274 2724 9276
rect 2748 9274 2804 9276
rect 2828 9274 2884 9276
rect 2588 9222 2634 9274
rect 2634 9222 2644 9274
rect 2668 9222 2698 9274
rect 2698 9222 2710 9274
rect 2710 9222 2724 9274
rect 2748 9222 2762 9274
rect 2762 9222 2774 9274
rect 2774 9222 2804 9274
rect 2828 9222 2838 9274
rect 2838 9222 2884 9274
rect 2588 9220 2644 9222
rect 2668 9220 2724 9222
rect 2748 9220 2804 9222
rect 2828 9220 2884 9222
rect 2410 8880 2466 8936
rect 1582 3576 1638 3632
rect 2134 5616 2190 5672
rect 2588 8186 2644 8188
rect 2668 8186 2724 8188
rect 2748 8186 2804 8188
rect 2828 8186 2884 8188
rect 2588 8134 2634 8186
rect 2634 8134 2644 8186
rect 2668 8134 2698 8186
rect 2698 8134 2710 8186
rect 2710 8134 2724 8186
rect 2748 8134 2762 8186
rect 2762 8134 2774 8186
rect 2774 8134 2804 8186
rect 2828 8134 2838 8186
rect 2838 8134 2884 8186
rect 2588 8132 2644 8134
rect 2668 8132 2724 8134
rect 2748 8132 2804 8134
rect 2828 8132 2884 8134
rect 2588 7098 2644 7100
rect 2668 7098 2724 7100
rect 2748 7098 2804 7100
rect 2828 7098 2884 7100
rect 2588 7046 2634 7098
rect 2634 7046 2644 7098
rect 2668 7046 2698 7098
rect 2698 7046 2710 7098
rect 2710 7046 2724 7098
rect 2748 7046 2762 7098
rect 2762 7046 2774 7098
rect 2774 7046 2804 7098
rect 2828 7046 2838 7098
rect 2838 7046 2884 7098
rect 2588 7044 2644 7046
rect 2668 7044 2724 7046
rect 2748 7044 2804 7046
rect 2828 7044 2884 7046
rect 2502 6704 2558 6760
rect 3606 9424 3662 9480
rect 2588 6010 2644 6012
rect 2668 6010 2724 6012
rect 2748 6010 2804 6012
rect 2828 6010 2884 6012
rect 2588 5958 2634 6010
rect 2634 5958 2644 6010
rect 2668 5958 2698 6010
rect 2698 5958 2710 6010
rect 2710 5958 2724 6010
rect 2748 5958 2762 6010
rect 2762 5958 2774 6010
rect 2774 5958 2804 6010
rect 2828 5958 2838 6010
rect 2838 5958 2884 6010
rect 2588 5956 2644 5958
rect 2668 5956 2724 5958
rect 2748 5956 2804 5958
rect 2828 5956 2884 5958
rect 2588 4922 2644 4924
rect 2668 4922 2724 4924
rect 2748 4922 2804 4924
rect 2828 4922 2884 4924
rect 2588 4870 2634 4922
rect 2634 4870 2644 4922
rect 2668 4870 2698 4922
rect 2698 4870 2710 4922
rect 2710 4870 2724 4922
rect 2748 4870 2762 4922
rect 2762 4870 2774 4922
rect 2774 4870 2804 4922
rect 2828 4870 2838 4922
rect 2838 4870 2884 4922
rect 2588 4868 2644 4870
rect 2668 4868 2724 4870
rect 2748 4868 2804 4870
rect 2828 4868 2884 4870
rect 2594 4156 2596 4176
rect 2596 4156 2648 4176
rect 2648 4156 2650 4176
rect 2594 4120 2650 4156
rect 2962 3984 3018 4040
rect 2588 3834 2644 3836
rect 2668 3834 2724 3836
rect 2748 3834 2804 3836
rect 2828 3834 2884 3836
rect 2588 3782 2634 3834
rect 2634 3782 2644 3834
rect 2668 3782 2698 3834
rect 2698 3782 2710 3834
rect 2710 3782 2724 3834
rect 2748 3782 2762 3834
rect 2762 3782 2774 3834
rect 2774 3782 2804 3834
rect 2828 3782 2838 3834
rect 2838 3782 2884 3834
rect 2588 3780 2644 3782
rect 2668 3780 2724 3782
rect 2748 3780 2804 3782
rect 2828 3780 2884 3782
rect 2962 3732 3018 3768
rect 2962 3712 2964 3732
rect 2964 3712 3016 3732
rect 3016 3712 3018 3732
rect 2588 2746 2644 2748
rect 2668 2746 2724 2748
rect 2748 2746 2804 2748
rect 2828 2746 2884 2748
rect 2588 2694 2634 2746
rect 2634 2694 2644 2746
rect 2668 2694 2698 2746
rect 2698 2694 2710 2746
rect 2710 2694 2724 2746
rect 2748 2694 2762 2746
rect 2762 2694 2774 2746
rect 2774 2694 2804 2746
rect 2828 2694 2838 2746
rect 2838 2694 2884 2746
rect 2588 2692 2644 2694
rect 2668 2692 2724 2694
rect 2748 2692 2804 2694
rect 2828 2692 2884 2694
rect 3974 11056 4030 11112
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4266 10906
rect 4266 10854 4276 10906
rect 4300 10854 4330 10906
rect 4330 10854 4342 10906
rect 4342 10854 4356 10906
rect 4380 10854 4394 10906
rect 4394 10854 4406 10906
rect 4406 10854 4436 10906
rect 4460 10854 4470 10906
rect 4470 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 3974 10548 3976 10568
rect 3976 10548 4028 10568
rect 4028 10548 4030 10568
rect 3974 10512 4030 10548
rect 3974 10240 4030 10296
rect 4250 10512 4306 10568
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4266 9818
rect 4266 9766 4276 9818
rect 4300 9766 4330 9818
rect 4330 9766 4342 9818
rect 4342 9766 4356 9818
rect 4380 9766 4394 9818
rect 4394 9766 4406 9818
rect 4406 9766 4436 9818
rect 4460 9766 4470 9818
rect 4470 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4618 9696 4674 9752
rect 4526 9424 4582 9480
rect 4250 8880 4306 8936
rect 4894 10376 4950 10432
rect 4802 9560 4858 9616
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4266 8730
rect 4266 8678 4276 8730
rect 4300 8678 4330 8730
rect 4330 8678 4342 8730
rect 4342 8678 4356 8730
rect 4380 8678 4394 8730
rect 4394 8678 4406 8730
rect 4406 8678 4436 8730
rect 4460 8678 4470 8730
rect 4470 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4266 7642
rect 4266 7590 4276 7642
rect 4300 7590 4330 7642
rect 4330 7590 4342 7642
rect 4342 7590 4356 7642
rect 4380 7590 4394 7642
rect 4394 7590 4406 7642
rect 4406 7590 4436 7642
rect 4460 7590 4470 7642
rect 4470 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 3422 3032 3478 3088
rect 4158 6704 4214 6760
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4266 6554
rect 4266 6502 4276 6554
rect 4300 6502 4330 6554
rect 4330 6502 4342 6554
rect 4342 6502 4356 6554
rect 4380 6502 4394 6554
rect 4394 6502 4406 6554
rect 4406 6502 4436 6554
rect 4460 6502 4470 6554
rect 4470 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4710 5480 4766 5536
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4266 5466
rect 4266 5414 4276 5466
rect 4300 5414 4330 5466
rect 4330 5414 4342 5466
rect 4342 5414 4356 5466
rect 4380 5414 4394 5466
rect 4394 5414 4406 5466
rect 4406 5414 4436 5466
rect 4460 5414 4470 5466
rect 4470 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4266 4378
rect 4266 4326 4276 4378
rect 4300 4326 4330 4378
rect 4330 4326 4342 4378
rect 4342 4326 4356 4378
rect 4380 4326 4394 4378
rect 4394 4326 4406 4378
rect 4406 4326 4436 4378
rect 4460 4326 4470 4378
rect 4470 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4986 9696 5042 9752
rect 5262 10956 5264 10976
rect 5264 10956 5316 10976
rect 5316 10956 5318 10976
rect 5262 10920 5318 10956
rect 5262 10240 5318 10296
rect 5354 8336 5410 8392
rect 5262 6160 5318 6216
rect 5078 5752 5134 5808
rect 4894 4528 4950 4584
rect 4802 3984 4858 4040
rect 4894 3712 4950 3768
rect 4066 3440 4122 3496
rect 4250 3440 4306 3496
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4266 3290
rect 4266 3238 4276 3290
rect 4300 3238 4330 3290
rect 4330 3238 4342 3290
rect 4342 3238 4356 3290
rect 4380 3238 4394 3290
rect 4394 3238 4406 3290
rect 4406 3238 4436 3290
rect 4460 3238 4470 3290
rect 4470 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4250 2644 4306 2680
rect 4250 2624 4252 2644
rect 4252 2624 4304 2644
rect 4304 2624 4306 2644
rect 4434 2760 4490 2816
rect 5852 10362 5908 10364
rect 5932 10362 5988 10364
rect 6012 10362 6068 10364
rect 6092 10362 6148 10364
rect 5852 10310 5898 10362
rect 5898 10310 5908 10362
rect 5932 10310 5962 10362
rect 5962 10310 5974 10362
rect 5974 10310 5988 10362
rect 6012 10310 6026 10362
rect 6026 10310 6038 10362
rect 6038 10310 6068 10362
rect 6092 10310 6102 10362
rect 6102 10310 6148 10362
rect 5852 10308 5908 10310
rect 5932 10308 5988 10310
rect 6012 10308 6068 10310
rect 6092 10308 6148 10310
rect 5852 9274 5908 9276
rect 5932 9274 5988 9276
rect 6012 9274 6068 9276
rect 6092 9274 6148 9276
rect 5852 9222 5898 9274
rect 5898 9222 5908 9274
rect 5932 9222 5962 9274
rect 5962 9222 5974 9274
rect 5974 9222 5988 9274
rect 6012 9222 6026 9274
rect 6026 9222 6038 9274
rect 6038 9222 6068 9274
rect 6092 9222 6102 9274
rect 6102 9222 6148 9274
rect 5852 9220 5908 9222
rect 5932 9220 5988 9222
rect 6012 9220 6068 9222
rect 6092 9220 6148 9222
rect 5852 8186 5908 8188
rect 5932 8186 5988 8188
rect 6012 8186 6068 8188
rect 6092 8186 6148 8188
rect 5852 8134 5898 8186
rect 5898 8134 5908 8186
rect 5932 8134 5962 8186
rect 5962 8134 5974 8186
rect 5974 8134 5988 8186
rect 6012 8134 6026 8186
rect 6026 8134 6038 8186
rect 6038 8134 6068 8186
rect 6092 8134 6102 8186
rect 6102 8134 6148 8186
rect 5852 8132 5908 8134
rect 5932 8132 5988 8134
rect 6012 8132 6068 8134
rect 6092 8132 6148 8134
rect 5852 7098 5908 7100
rect 5932 7098 5988 7100
rect 6012 7098 6068 7100
rect 6092 7098 6148 7100
rect 5852 7046 5898 7098
rect 5898 7046 5908 7098
rect 5932 7046 5962 7098
rect 5962 7046 5974 7098
rect 5974 7046 5988 7098
rect 6012 7046 6026 7098
rect 6026 7046 6038 7098
rect 6038 7046 6068 7098
rect 6092 7046 6102 7098
rect 6102 7046 6148 7098
rect 5852 7044 5908 7046
rect 5932 7044 5988 7046
rect 6012 7044 6068 7046
rect 6092 7044 6148 7046
rect 5262 5072 5318 5128
rect 5078 3712 5134 3768
rect 5262 4120 5318 4176
rect 5852 6010 5908 6012
rect 5932 6010 5988 6012
rect 6012 6010 6068 6012
rect 6092 6010 6148 6012
rect 5852 5958 5898 6010
rect 5898 5958 5908 6010
rect 5932 5958 5962 6010
rect 5962 5958 5974 6010
rect 5974 5958 5988 6010
rect 6012 5958 6026 6010
rect 6026 5958 6038 6010
rect 6038 5958 6068 6010
rect 6092 5958 6102 6010
rect 6102 5958 6148 6010
rect 5852 5956 5908 5958
rect 5932 5956 5988 5958
rect 6012 5956 6068 5958
rect 6092 5956 6148 5958
rect 5852 4922 5908 4924
rect 5932 4922 5988 4924
rect 6012 4922 6068 4924
rect 6092 4922 6148 4924
rect 5852 4870 5898 4922
rect 5898 4870 5908 4922
rect 5932 4870 5962 4922
rect 5962 4870 5974 4922
rect 5974 4870 5988 4922
rect 6012 4870 6026 4922
rect 6026 4870 6038 4922
rect 6038 4870 6068 4922
rect 6092 4870 6102 4922
rect 6102 4870 6148 4922
rect 5852 4868 5908 4870
rect 5932 4868 5988 4870
rect 6012 4868 6068 4870
rect 6092 4868 6148 4870
rect 5852 3834 5908 3836
rect 5932 3834 5988 3836
rect 6012 3834 6068 3836
rect 6092 3834 6148 3836
rect 5852 3782 5898 3834
rect 5898 3782 5908 3834
rect 5932 3782 5962 3834
rect 5962 3782 5974 3834
rect 5974 3782 5988 3834
rect 6012 3782 6026 3834
rect 6026 3782 6038 3834
rect 6038 3782 6068 3834
rect 6092 3782 6102 3834
rect 6102 3782 6148 3834
rect 5852 3780 5908 3782
rect 5932 3780 5988 3782
rect 6012 3780 6068 3782
rect 6092 3780 6148 3782
rect 5262 2896 5318 2952
rect 5262 2760 5318 2816
rect 6366 3712 6422 3768
rect 7484 10906 7540 10908
rect 7564 10906 7620 10908
rect 7644 10906 7700 10908
rect 7724 10906 7780 10908
rect 7484 10854 7530 10906
rect 7530 10854 7540 10906
rect 7564 10854 7594 10906
rect 7594 10854 7606 10906
rect 7606 10854 7620 10906
rect 7644 10854 7658 10906
rect 7658 10854 7670 10906
rect 7670 10854 7700 10906
rect 7724 10854 7734 10906
rect 7734 10854 7780 10906
rect 7484 10852 7540 10854
rect 7564 10852 7620 10854
rect 7644 10852 7700 10854
rect 7724 10852 7780 10854
rect 7562 10512 7618 10568
rect 7010 9696 7066 9752
rect 6918 9560 6974 9616
rect 7484 9818 7540 9820
rect 7564 9818 7620 9820
rect 7644 9818 7700 9820
rect 7724 9818 7780 9820
rect 7484 9766 7530 9818
rect 7530 9766 7540 9818
rect 7564 9766 7594 9818
rect 7594 9766 7606 9818
rect 7606 9766 7620 9818
rect 7644 9766 7658 9818
rect 7658 9766 7670 9818
rect 7670 9766 7700 9818
rect 7724 9766 7734 9818
rect 7734 9766 7780 9818
rect 7484 9764 7540 9766
rect 7564 9764 7620 9766
rect 7644 9764 7700 9766
rect 7724 9764 7780 9766
rect 7010 8880 7066 8936
rect 7010 8064 7066 8120
rect 7010 7928 7066 7984
rect 5538 3052 5594 3088
rect 5538 3032 5540 3052
rect 5540 3032 5592 3052
rect 5592 3032 5594 3052
rect 5852 2746 5908 2748
rect 5932 2746 5988 2748
rect 6012 2746 6068 2748
rect 6092 2746 6148 2748
rect 5852 2694 5898 2746
rect 5898 2694 5908 2746
rect 5932 2694 5962 2746
rect 5962 2694 5974 2746
rect 5974 2694 5988 2746
rect 6012 2694 6026 2746
rect 6026 2694 6038 2746
rect 6038 2694 6068 2746
rect 6092 2694 6102 2746
rect 6102 2694 6148 2746
rect 5852 2692 5908 2694
rect 5932 2692 5988 2694
rect 6012 2692 6068 2694
rect 6092 2692 6148 2694
rect 6458 3440 6514 3496
rect 6642 5516 6644 5536
rect 6644 5516 6696 5536
rect 6696 5516 6698 5536
rect 6642 5480 6698 5516
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4266 2202
rect 4266 2150 4276 2202
rect 4300 2150 4330 2202
rect 4330 2150 4342 2202
rect 4342 2150 4356 2202
rect 4380 2150 4394 2202
rect 4394 2150 4406 2202
rect 4406 2150 4436 2202
rect 4460 2150 4470 2202
rect 4470 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 7102 5616 7158 5672
rect 7484 8730 7540 8732
rect 7564 8730 7620 8732
rect 7644 8730 7700 8732
rect 7724 8730 7780 8732
rect 7484 8678 7530 8730
rect 7530 8678 7540 8730
rect 7564 8678 7594 8730
rect 7594 8678 7606 8730
rect 7606 8678 7620 8730
rect 7644 8678 7658 8730
rect 7658 8678 7670 8730
rect 7670 8678 7700 8730
rect 7724 8678 7734 8730
rect 7734 8678 7780 8730
rect 7484 8676 7540 8678
rect 7564 8676 7620 8678
rect 7644 8676 7700 8678
rect 7724 8676 7780 8678
rect 7484 7642 7540 7644
rect 7564 7642 7620 7644
rect 7644 7642 7700 7644
rect 7724 7642 7780 7644
rect 7484 7590 7530 7642
rect 7530 7590 7540 7642
rect 7564 7590 7594 7642
rect 7594 7590 7606 7642
rect 7606 7590 7620 7642
rect 7644 7590 7658 7642
rect 7658 7590 7670 7642
rect 7670 7590 7700 7642
rect 7724 7590 7734 7642
rect 7734 7590 7780 7642
rect 7484 7588 7540 7590
rect 7564 7588 7620 7590
rect 7644 7588 7700 7590
rect 7724 7588 7780 7590
rect 7286 5208 7342 5264
rect 7484 6554 7540 6556
rect 7564 6554 7620 6556
rect 7644 6554 7700 6556
rect 7724 6554 7780 6556
rect 7484 6502 7530 6554
rect 7530 6502 7540 6554
rect 7564 6502 7594 6554
rect 7594 6502 7606 6554
rect 7606 6502 7620 6554
rect 7644 6502 7658 6554
rect 7658 6502 7670 6554
rect 7670 6502 7700 6554
rect 7724 6502 7734 6554
rect 7734 6502 7780 6554
rect 7484 6500 7540 6502
rect 7564 6500 7620 6502
rect 7644 6500 7700 6502
rect 7724 6500 7780 6502
rect 7930 6432 7986 6488
rect 7484 5466 7540 5468
rect 7564 5466 7620 5468
rect 7644 5466 7700 5468
rect 7724 5466 7780 5468
rect 7484 5414 7530 5466
rect 7530 5414 7540 5466
rect 7564 5414 7594 5466
rect 7594 5414 7606 5466
rect 7606 5414 7620 5466
rect 7644 5414 7658 5466
rect 7658 5414 7670 5466
rect 7670 5414 7700 5466
rect 7724 5414 7734 5466
rect 7734 5414 7780 5466
rect 7484 5412 7540 5414
rect 7564 5412 7620 5414
rect 7644 5412 7700 5414
rect 7724 5412 7780 5414
rect 7102 3984 7158 4040
rect 7484 4378 7540 4380
rect 7564 4378 7620 4380
rect 7644 4378 7700 4380
rect 7724 4378 7780 4380
rect 7484 4326 7530 4378
rect 7530 4326 7540 4378
rect 7564 4326 7594 4378
rect 7594 4326 7606 4378
rect 7606 4326 7620 4378
rect 7644 4326 7658 4378
rect 7658 4326 7670 4378
rect 7670 4326 7700 4378
rect 7724 4326 7734 4378
rect 7734 4326 7780 4378
rect 7484 4324 7540 4326
rect 7564 4324 7620 4326
rect 7644 4324 7700 4326
rect 7724 4324 7780 4326
rect 7010 3476 7012 3496
rect 7012 3476 7064 3496
rect 7064 3476 7066 3496
rect 7010 3440 7066 3476
rect 7484 3290 7540 3292
rect 7564 3290 7620 3292
rect 7644 3290 7700 3292
rect 7724 3290 7780 3292
rect 7484 3238 7530 3290
rect 7530 3238 7540 3290
rect 7564 3238 7594 3290
rect 7594 3238 7606 3290
rect 7606 3238 7620 3290
rect 7644 3238 7658 3290
rect 7658 3238 7670 3290
rect 7670 3238 7700 3290
rect 7724 3238 7734 3290
rect 7734 3238 7780 3290
rect 7484 3236 7540 3238
rect 7564 3236 7620 3238
rect 7644 3236 7700 3238
rect 7724 3236 7780 3238
rect 8206 9560 8262 9616
rect 8114 9424 8170 9480
rect 8114 6704 8170 6760
rect 8390 5072 8446 5128
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 9276 10362 9332 10364
rect 9356 10362 9412 10364
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9238 10362
rect 9238 10310 9252 10362
rect 9276 10310 9290 10362
rect 9290 10310 9302 10362
rect 9302 10310 9332 10362
rect 9356 10310 9366 10362
rect 9366 10310 9412 10362
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 9276 10308 9332 10310
rect 9356 10308 9412 10310
rect 9126 9560 9182 9616
rect 9494 9444 9550 9480
rect 9494 9424 9496 9444
rect 9496 9424 9548 9444
rect 9548 9424 9550 9444
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 9276 9274 9332 9276
rect 9356 9274 9412 9276
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9238 9274
rect 9238 9222 9252 9274
rect 9276 9222 9290 9274
rect 9290 9222 9302 9274
rect 9302 9222 9332 9274
rect 9356 9222 9366 9274
rect 9366 9222 9412 9274
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 9276 9220 9332 9222
rect 9356 9220 9412 9222
rect 9494 8916 9496 8936
rect 9496 8916 9548 8936
rect 9548 8916 9550 8936
rect 9494 8880 9550 8916
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 9276 8186 9332 8188
rect 9356 8186 9412 8188
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9238 8186
rect 9238 8134 9252 8186
rect 9276 8134 9290 8186
rect 9290 8134 9302 8186
rect 9302 8134 9332 8186
rect 9356 8134 9366 8186
rect 9366 8134 9412 8186
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 9276 8132 9332 8134
rect 9356 8132 9412 8134
rect 8758 5208 8814 5264
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 9276 7098 9332 7100
rect 9356 7098 9412 7100
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9238 7098
rect 9238 7046 9252 7098
rect 9276 7046 9290 7098
rect 9290 7046 9302 7098
rect 9302 7046 9332 7098
rect 9356 7046 9366 7098
rect 9366 7046 9412 7098
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 9276 7044 9332 7046
rect 9356 7044 9412 7046
rect 9310 6704 9366 6760
rect 10046 6976 10102 7032
rect 9678 6840 9734 6896
rect 9310 6604 9312 6624
rect 9312 6604 9364 6624
rect 9364 6604 9366 6624
rect 9310 6568 9366 6604
rect 9402 6432 9458 6488
rect 9126 6160 9182 6216
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 9276 6010 9332 6012
rect 9356 6010 9412 6012
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9238 6010
rect 9238 5958 9252 6010
rect 9276 5958 9290 6010
rect 9290 5958 9302 6010
rect 9302 5958 9332 6010
rect 9356 5958 9366 6010
rect 9366 5958 9412 6010
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 9276 5956 9332 5958
rect 9356 5956 9412 5958
rect 9494 5752 9550 5808
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 9276 4922 9332 4924
rect 9356 4922 9412 4924
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9238 4922
rect 9238 4870 9252 4922
rect 9276 4870 9290 4922
rect 9290 4870 9302 4922
rect 9302 4870 9332 4922
rect 9356 4870 9366 4922
rect 9366 4870 9412 4922
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 9276 4868 9332 4870
rect 9356 4868 9412 4870
rect 9586 5228 9642 5264
rect 9586 5208 9588 5228
rect 9588 5208 9640 5228
rect 9640 5208 9642 5228
rect 8758 3732 8814 3768
rect 8758 3712 8760 3732
rect 8760 3712 8812 3732
rect 8812 3712 8814 3732
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 9276 3834 9332 3836
rect 9356 3834 9412 3836
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9238 3834
rect 9238 3782 9252 3834
rect 9276 3782 9290 3834
rect 9290 3782 9302 3834
rect 9302 3782 9332 3834
rect 9356 3782 9366 3834
rect 9366 3782 9412 3834
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 9276 3780 9332 3782
rect 9356 3780 9412 3782
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 9276 2746 9332 2748
rect 9356 2746 9412 2748
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9238 2746
rect 9238 2694 9252 2746
rect 9276 2694 9290 2746
rect 9290 2694 9302 2746
rect 9302 2694 9332 2746
rect 9356 2694 9366 2746
rect 9366 2694 9412 2746
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 9276 2692 9332 2694
rect 9356 2692 9412 2694
rect 7484 2202 7540 2204
rect 7564 2202 7620 2204
rect 7644 2202 7700 2204
rect 7724 2202 7780 2204
rect 7484 2150 7530 2202
rect 7530 2150 7540 2202
rect 7564 2150 7594 2202
rect 7594 2150 7606 2202
rect 7606 2150 7620 2202
rect 7644 2150 7658 2202
rect 7658 2150 7670 2202
rect 7670 2150 7700 2202
rect 7724 2150 7734 2202
rect 7734 2150 7780 2202
rect 7484 2148 7540 2150
rect 7564 2148 7620 2150
rect 7644 2148 7700 2150
rect 7724 2148 7780 2150
<< metal3 >>
rect 2576 11456 2896 11457
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 11391 2896 11392
rect 5840 11456 6160 11457
rect 5840 11392 5848 11456
rect 5912 11392 5928 11456
rect 5992 11392 6008 11456
rect 6072 11392 6088 11456
rect 6152 11392 6160 11456
rect 5840 11391 6160 11392
rect 9104 11456 9424 11457
rect 9104 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9272 11456
rect 9336 11392 9352 11456
rect 9416 11392 9424 11456
rect 9104 11391 9424 11392
rect 3233 11114 3299 11117
rect 3969 11116 4035 11117
rect 3366 11114 3372 11116
rect 3233 11112 3372 11114
rect 3233 11056 3238 11112
rect 3294 11056 3372 11112
rect 3233 11054 3372 11056
rect 3233 11051 3299 11054
rect 3366 11052 3372 11054
rect 3436 11052 3442 11116
rect 3918 11114 3924 11116
rect 3878 11054 3924 11114
rect 3988 11112 4035 11116
rect 4030 11056 4035 11112
rect 3918 11052 3924 11054
rect 3988 11052 4035 11056
rect 3969 11051 4035 11052
rect 5257 10980 5323 10981
rect 5206 10916 5212 10980
rect 5276 10978 5323 10980
rect 5276 10976 5368 10978
rect 5318 10920 5368 10976
rect 5276 10918 5368 10920
rect 5276 10916 5323 10918
rect 5257 10915 5323 10916
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 7472 10912 7792 10913
rect 7472 10848 7480 10912
rect 7544 10848 7560 10912
rect 7624 10848 7640 10912
rect 7704 10848 7720 10912
rect 7784 10848 7792 10912
rect 7472 10847 7792 10848
rect 3969 10570 4035 10573
rect 4245 10570 4311 10573
rect 7557 10570 7623 10573
rect 3969 10568 7623 10570
rect 3969 10512 3974 10568
rect 4030 10512 4250 10568
rect 4306 10512 7562 10568
rect 7618 10512 7623 10568
rect 3969 10510 7623 10512
rect 3969 10507 4035 10510
rect 4245 10507 4311 10510
rect 7557 10507 7623 10510
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4654 10372 4660 10436
rect 4724 10434 4730 10436
rect 4889 10434 4955 10437
rect 4724 10432 4955 10434
rect 4724 10376 4894 10432
rect 4950 10376 4955 10432
rect 4724 10374 4955 10376
rect 4724 10372 4730 10374
rect 4889 10371 4955 10374
rect 2576 10368 2896 10369
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 10303 2896 10304
rect 5840 10368 6160 10369
rect 5840 10304 5848 10368
rect 5912 10304 5928 10368
rect 5992 10304 6008 10368
rect 6072 10304 6088 10368
rect 6152 10304 6160 10368
rect 5840 10303 6160 10304
rect 9104 10368 9424 10369
rect 9104 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9272 10368
rect 9336 10304 9352 10368
rect 9416 10304 9424 10368
rect 9104 10303 9424 10304
rect 3969 10298 4035 10301
rect 5257 10298 5323 10301
rect 3969 10296 5323 10298
rect 3969 10240 3974 10296
rect 4030 10240 5262 10296
rect 5318 10240 5323 10296
rect 3969 10238 5323 10240
rect 3969 10235 4035 10238
rect 5257 10235 5323 10238
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 7472 9824 7792 9825
rect 7472 9760 7480 9824
rect 7544 9760 7560 9824
rect 7624 9760 7640 9824
rect 7704 9760 7720 9824
rect 7784 9760 7792 9824
rect 7472 9759 7792 9760
rect 4613 9754 4679 9757
rect 4981 9754 5047 9757
rect 7005 9754 7071 9757
rect 4613 9752 7071 9754
rect 4613 9696 4618 9752
rect 4674 9696 4986 9752
rect 5042 9696 7010 9752
rect 7066 9696 7071 9752
rect 4613 9694 7071 9696
rect 4613 9691 4679 9694
rect 4981 9691 5047 9694
rect 7005 9691 7071 9694
rect 1761 9618 1827 9621
rect 4797 9618 4863 9621
rect 1761 9616 4863 9618
rect 1761 9560 1766 9616
rect 1822 9560 4802 9616
rect 4858 9560 4863 9616
rect 1761 9558 4863 9560
rect 1761 9555 1827 9558
rect 4797 9555 4863 9558
rect 6913 9618 6979 9621
rect 8201 9618 8267 9621
rect 9121 9618 9187 9621
rect 6913 9616 9187 9618
rect 6913 9560 6918 9616
rect 6974 9560 8206 9616
rect 8262 9560 9126 9616
rect 9182 9560 9187 9616
rect 6913 9558 9187 9560
rect 6913 9555 6979 9558
rect 8201 9555 8267 9558
rect 9121 9555 9187 9558
rect 3601 9482 3667 9485
rect 4521 9482 4587 9485
rect 3601 9480 4587 9482
rect 3601 9424 3606 9480
rect 3662 9424 4526 9480
rect 4582 9424 4587 9480
rect 3601 9422 4587 9424
rect 3601 9419 3667 9422
rect 4521 9419 4587 9422
rect 8109 9482 8175 9485
rect 9489 9482 9555 9485
rect 8109 9480 9555 9482
rect 8109 9424 8114 9480
rect 8170 9424 9494 9480
rect 9550 9424 9555 9480
rect 8109 9422 9555 9424
rect 8109 9419 8175 9422
rect 9489 9419 9555 9422
rect 2576 9280 2896 9281
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 9215 2896 9216
rect 5840 9280 6160 9281
rect 5840 9216 5848 9280
rect 5912 9216 5928 9280
rect 5992 9216 6008 9280
rect 6072 9216 6088 9280
rect 6152 9216 6160 9280
rect 5840 9215 6160 9216
rect 9104 9280 9424 9281
rect 9104 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9272 9280
rect 9336 9216 9352 9280
rect 9416 9216 9424 9280
rect 9104 9215 9424 9216
rect 2129 8938 2195 8941
rect 2405 8938 2471 8941
rect 4245 8938 4311 8941
rect 2129 8936 4311 8938
rect 2129 8880 2134 8936
rect 2190 8880 2410 8936
rect 2466 8880 4250 8936
rect 4306 8880 4311 8936
rect 2129 8878 4311 8880
rect 2129 8875 2195 8878
rect 2405 8875 2471 8878
rect 4245 8875 4311 8878
rect 7005 8938 7071 8941
rect 9489 8938 9555 8941
rect 7005 8936 9555 8938
rect 7005 8880 7010 8936
rect 7066 8880 9494 8936
rect 9550 8880 9555 8936
rect 7005 8878 9555 8880
rect 7005 8875 7071 8878
rect 9489 8875 9555 8878
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 7472 8736 7792 8737
rect 7472 8672 7480 8736
rect 7544 8672 7560 8736
rect 7624 8672 7640 8736
rect 7704 8672 7720 8736
rect 7784 8672 7792 8736
rect 7472 8671 7792 8672
rect 5349 8396 5415 8397
rect 5349 8392 5396 8396
rect 5460 8394 5466 8396
rect 5349 8336 5354 8392
rect 5349 8332 5396 8336
rect 5460 8334 5506 8394
rect 5460 8332 5466 8334
rect 5349 8331 5415 8332
rect 2576 8192 2896 8193
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 8127 2896 8128
rect 5840 8192 6160 8193
rect 5840 8128 5848 8192
rect 5912 8128 5928 8192
rect 5992 8128 6008 8192
rect 6072 8128 6088 8192
rect 6152 8128 6160 8192
rect 5840 8127 6160 8128
rect 9104 8192 9424 8193
rect 9104 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9272 8192
rect 9336 8128 9352 8192
rect 9416 8128 9424 8192
rect 9104 8127 9424 8128
rect 7005 8124 7071 8125
rect 7005 8122 7052 8124
rect 6960 8120 7052 8122
rect 6960 8064 7010 8120
rect 6960 8062 7052 8064
rect 7005 8060 7052 8062
rect 7116 8060 7122 8124
rect 7005 8059 7071 8060
rect 3918 7924 3924 7988
rect 3988 7986 3994 7988
rect 7005 7986 7071 7989
rect 3988 7984 7071 7986
rect 3988 7928 7010 7984
rect 7066 7928 7071 7984
rect 3988 7926 7071 7928
rect 3988 7924 3994 7926
rect 7005 7923 7071 7926
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 7472 7648 7792 7649
rect 7472 7584 7480 7648
rect 7544 7584 7560 7648
rect 7624 7584 7640 7648
rect 7704 7584 7720 7648
rect 7784 7584 7792 7648
rect 7472 7583 7792 7584
rect 2576 7104 2896 7105
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2576 7039 2896 7040
rect 5840 7104 6160 7105
rect 5840 7040 5848 7104
rect 5912 7040 5928 7104
rect 5992 7040 6008 7104
rect 6072 7040 6088 7104
rect 6152 7040 6160 7104
rect 5840 7039 6160 7040
rect 9104 7104 9424 7105
rect 9104 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9272 7104
rect 9336 7040 9352 7104
rect 9416 7040 9424 7104
rect 9104 7039 9424 7040
rect 10041 7034 10107 7037
rect 11200 7034 12000 7064
rect 10041 7032 12000 7034
rect 10041 6976 10046 7032
rect 10102 6976 12000 7032
rect 10041 6974 12000 6976
rect 10041 6971 10107 6974
rect 11200 6944 12000 6974
rect 5206 6836 5212 6900
rect 5276 6898 5282 6900
rect 9673 6898 9739 6901
rect 5276 6896 9739 6898
rect 5276 6840 9678 6896
rect 9734 6840 9739 6896
rect 5276 6838 9739 6840
rect 5276 6836 5282 6838
rect 9673 6835 9739 6838
rect 2497 6762 2563 6765
rect 4153 6762 4219 6765
rect 8109 6762 8175 6765
rect 9305 6762 9371 6765
rect 2497 6760 7988 6762
rect 2497 6704 2502 6760
rect 2558 6704 4158 6760
rect 4214 6704 7988 6760
rect 2497 6702 7988 6704
rect 2497 6699 2563 6702
rect 4153 6699 4219 6702
rect 7928 6626 7988 6702
rect 8109 6760 9371 6762
rect 8109 6704 8114 6760
rect 8170 6704 9310 6760
rect 9366 6704 9371 6760
rect 8109 6702 9371 6704
rect 8109 6699 8175 6702
rect 9305 6699 9371 6702
rect 9305 6626 9371 6629
rect 7928 6624 9371 6626
rect 7928 6568 9310 6624
rect 9366 6568 9371 6624
rect 7928 6566 9371 6568
rect 9305 6563 9371 6566
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 7472 6560 7792 6561
rect 7472 6496 7480 6560
rect 7544 6496 7560 6560
rect 7624 6496 7640 6560
rect 7704 6496 7720 6560
rect 7784 6496 7792 6560
rect 7472 6495 7792 6496
rect 7925 6490 7991 6493
rect 9397 6490 9463 6493
rect 7925 6488 9463 6490
rect 7925 6432 7930 6488
rect 7986 6432 9402 6488
rect 9458 6432 9463 6488
rect 7925 6430 9463 6432
rect 7925 6427 7991 6430
rect 9397 6427 9463 6430
rect 5257 6218 5323 6221
rect 9121 6218 9187 6221
rect 5257 6216 9187 6218
rect 5257 6160 5262 6216
rect 5318 6160 9126 6216
rect 9182 6160 9187 6216
rect 5257 6158 9187 6160
rect 5257 6155 5323 6158
rect 9121 6155 9187 6158
rect 2576 6016 2896 6017
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 5951 2896 5952
rect 5840 6016 6160 6017
rect 5840 5952 5848 6016
rect 5912 5952 5928 6016
rect 5992 5952 6008 6016
rect 6072 5952 6088 6016
rect 6152 5952 6160 6016
rect 5840 5951 6160 5952
rect 9104 6016 9424 6017
rect 9104 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9272 6016
rect 9336 5952 9352 6016
rect 9416 5952 9424 6016
rect 9104 5951 9424 5952
rect 5073 5810 5139 5813
rect 9489 5810 9555 5813
rect 5073 5808 9555 5810
rect 5073 5752 5078 5808
rect 5134 5752 9494 5808
rect 9550 5752 9555 5808
rect 5073 5750 9555 5752
rect 5073 5747 5139 5750
rect 9489 5747 9555 5750
rect 2129 5674 2195 5677
rect 7097 5674 7163 5677
rect 2129 5672 7163 5674
rect 2129 5616 2134 5672
rect 2190 5616 7102 5672
rect 7158 5616 7163 5672
rect 2129 5614 7163 5616
rect 2129 5611 2195 5614
rect 7097 5611 7163 5614
rect 4705 5538 4771 5541
rect 6637 5538 6703 5541
rect 4705 5536 6703 5538
rect 4705 5480 4710 5536
rect 4766 5480 6642 5536
rect 6698 5480 6703 5536
rect 4705 5478 6703 5480
rect 4705 5475 4771 5478
rect 6637 5475 6703 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 7472 5472 7792 5473
rect 7472 5408 7480 5472
rect 7544 5408 7560 5472
rect 7624 5408 7640 5472
rect 7704 5408 7720 5472
rect 7784 5408 7792 5472
rect 7472 5407 7792 5408
rect 7281 5266 7347 5269
rect 8753 5266 8819 5269
rect 9581 5266 9647 5269
rect 7281 5264 9647 5266
rect 7281 5208 7286 5264
rect 7342 5208 8758 5264
rect 8814 5208 9586 5264
rect 9642 5208 9647 5264
rect 7281 5206 9647 5208
rect 7281 5203 7347 5206
rect 8753 5203 8819 5206
rect 9581 5203 9647 5206
rect 5257 5130 5323 5133
rect 8385 5130 8451 5133
rect 5257 5128 8451 5130
rect 5257 5072 5262 5128
rect 5318 5072 8390 5128
rect 8446 5072 8451 5128
rect 5257 5070 8451 5072
rect 5257 5067 5323 5070
rect 8385 5067 8451 5070
rect 2576 4928 2896 4929
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 4863 2896 4864
rect 5840 4928 6160 4929
rect 5840 4864 5848 4928
rect 5912 4864 5928 4928
rect 5992 4864 6008 4928
rect 6072 4864 6088 4928
rect 6152 4864 6160 4928
rect 5840 4863 6160 4864
rect 9104 4928 9424 4929
rect 9104 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9272 4928
rect 9336 4864 9352 4928
rect 9416 4864 9424 4928
rect 9104 4863 9424 4864
rect 4889 4586 4955 4589
rect 5206 4586 5212 4588
rect 4889 4584 5212 4586
rect 4889 4528 4894 4584
rect 4950 4528 5212 4584
rect 4889 4526 5212 4528
rect 4889 4523 4955 4526
rect 5206 4524 5212 4526
rect 5276 4524 5282 4588
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 7472 4384 7792 4385
rect 7472 4320 7480 4384
rect 7544 4320 7560 4384
rect 7624 4320 7640 4384
rect 7704 4320 7720 4384
rect 7784 4320 7792 4384
rect 7472 4319 7792 4320
rect 2589 4178 2655 4181
rect 5257 4178 5323 4181
rect 2589 4176 5323 4178
rect 2589 4120 2594 4176
rect 2650 4120 5262 4176
rect 5318 4120 5323 4176
rect 2589 4118 5323 4120
rect 2589 4115 2655 4118
rect 5257 4115 5323 4118
rect 2957 4042 3023 4045
rect 4797 4042 4863 4045
rect 2957 4040 4863 4042
rect 2957 3984 2962 4040
rect 3018 3984 4802 4040
rect 4858 3984 4863 4040
rect 2957 3982 4863 3984
rect 2957 3979 3023 3982
rect 4797 3979 4863 3982
rect 5390 3980 5396 4044
rect 5460 4042 5466 4044
rect 7097 4042 7163 4045
rect 5460 4040 7163 4042
rect 5460 3984 7102 4040
rect 7158 3984 7163 4040
rect 5460 3982 7163 3984
rect 5460 3980 5466 3982
rect 7097 3979 7163 3982
rect 2576 3840 2896 3841
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 3775 2896 3776
rect 5840 3840 6160 3841
rect 5840 3776 5848 3840
rect 5912 3776 5928 3840
rect 5992 3776 6008 3840
rect 6072 3776 6088 3840
rect 6152 3776 6160 3840
rect 5840 3775 6160 3776
rect 9104 3840 9424 3841
rect 9104 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9272 3840
rect 9336 3776 9352 3840
rect 9416 3776 9424 3840
rect 9104 3775 9424 3776
rect 2957 3770 3023 3773
rect 4654 3770 4660 3772
rect 2957 3768 4660 3770
rect 2957 3712 2962 3768
rect 3018 3712 4660 3768
rect 2957 3710 4660 3712
rect 2957 3707 3023 3710
rect 4654 3708 4660 3710
rect 4724 3708 4730 3772
rect 4889 3770 4955 3773
rect 5073 3770 5139 3773
rect 4846 3768 5139 3770
rect 4846 3712 4894 3768
rect 4950 3712 5078 3768
rect 5134 3712 5139 3768
rect 4846 3710 5139 3712
rect 4846 3707 4955 3710
rect 5073 3707 5139 3710
rect 6361 3770 6427 3773
rect 8753 3770 8819 3773
rect 6361 3768 8819 3770
rect 6361 3712 6366 3768
rect 6422 3712 8758 3768
rect 8814 3712 8819 3768
rect 6361 3710 8819 3712
rect 6361 3707 6427 3710
rect 8753 3707 8819 3710
rect 1577 3634 1643 3637
rect 4846 3634 4906 3707
rect 1577 3632 4906 3634
rect 1577 3576 1582 3632
rect 1638 3576 4906 3632
rect 1577 3574 4906 3576
rect 1577 3571 1643 3574
rect 0 3498 800 3528
rect 4061 3498 4127 3501
rect 0 3496 4127 3498
rect 0 3440 4066 3496
rect 4122 3440 4127 3496
rect 0 3438 4127 3440
rect 0 3408 800 3438
rect 4061 3435 4127 3438
rect 4245 3498 4311 3501
rect 6453 3498 6519 3501
rect 4245 3496 6519 3498
rect 4245 3440 4250 3496
rect 4306 3440 6458 3496
rect 6514 3440 6519 3496
rect 4245 3438 6519 3440
rect 4245 3435 4311 3438
rect 6453 3435 6519 3438
rect 7005 3500 7071 3501
rect 7005 3496 7052 3500
rect 7116 3498 7122 3500
rect 7005 3440 7010 3496
rect 7005 3436 7052 3440
rect 7116 3438 7162 3498
rect 7116 3436 7122 3438
rect 7005 3435 7071 3436
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 7472 3296 7792 3297
rect 7472 3232 7480 3296
rect 7544 3232 7560 3296
rect 7624 3232 7640 3296
rect 7704 3232 7720 3296
rect 7784 3232 7792 3296
rect 7472 3231 7792 3232
rect 3417 3090 3483 3093
rect 5533 3090 5599 3093
rect 3417 3088 5599 3090
rect 3417 3032 3422 3088
rect 3478 3032 5538 3088
rect 5594 3032 5599 3088
rect 3417 3030 5599 3032
rect 3417 3027 3483 3030
rect 5533 3027 5599 3030
rect 5257 2954 5323 2957
rect 4662 2952 5323 2954
rect 4662 2896 5262 2952
rect 5318 2896 5323 2952
rect 4662 2894 5323 2896
rect 4429 2818 4495 2821
rect 4662 2818 4722 2894
rect 5257 2891 5323 2894
rect 5257 2820 5323 2821
rect 5206 2818 5212 2820
rect 4429 2816 4722 2818
rect 4429 2760 4434 2816
rect 4490 2760 4722 2816
rect 4429 2758 4722 2760
rect 5166 2758 5212 2818
rect 5276 2816 5323 2820
rect 5318 2760 5323 2816
rect 4429 2755 4495 2758
rect 5206 2756 5212 2758
rect 5276 2756 5323 2760
rect 5257 2755 5323 2756
rect 2576 2752 2896 2753
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2687 2896 2688
rect 5840 2752 6160 2753
rect 5840 2688 5848 2752
rect 5912 2688 5928 2752
rect 5992 2688 6008 2752
rect 6072 2688 6088 2752
rect 6152 2688 6160 2752
rect 5840 2687 6160 2688
rect 9104 2752 9424 2753
rect 9104 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9272 2752
rect 9336 2688 9352 2752
rect 9416 2688 9424 2752
rect 9104 2687 9424 2688
rect 3366 2620 3372 2684
rect 3436 2682 3442 2684
rect 4245 2682 4311 2685
rect 3436 2680 4311 2682
rect 3436 2624 4250 2680
rect 4306 2624 4311 2680
rect 3436 2622 4311 2624
rect 3436 2620 3442 2622
rect 4245 2619 4311 2622
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 7472 2208 7792 2209
rect 7472 2144 7480 2208
rect 7544 2144 7560 2208
rect 7624 2144 7640 2208
rect 7704 2144 7720 2208
rect 7784 2144 7792 2208
rect 7472 2143 7792 2144
<< via3 >>
rect 2584 11452 2648 11456
rect 2584 11396 2588 11452
rect 2588 11396 2644 11452
rect 2644 11396 2648 11452
rect 2584 11392 2648 11396
rect 2664 11452 2728 11456
rect 2664 11396 2668 11452
rect 2668 11396 2724 11452
rect 2724 11396 2728 11452
rect 2664 11392 2728 11396
rect 2744 11452 2808 11456
rect 2744 11396 2748 11452
rect 2748 11396 2804 11452
rect 2804 11396 2808 11452
rect 2744 11392 2808 11396
rect 2824 11452 2888 11456
rect 2824 11396 2828 11452
rect 2828 11396 2884 11452
rect 2884 11396 2888 11452
rect 2824 11392 2888 11396
rect 5848 11452 5912 11456
rect 5848 11396 5852 11452
rect 5852 11396 5908 11452
rect 5908 11396 5912 11452
rect 5848 11392 5912 11396
rect 5928 11452 5992 11456
rect 5928 11396 5932 11452
rect 5932 11396 5988 11452
rect 5988 11396 5992 11452
rect 5928 11392 5992 11396
rect 6008 11452 6072 11456
rect 6008 11396 6012 11452
rect 6012 11396 6068 11452
rect 6068 11396 6072 11452
rect 6008 11392 6072 11396
rect 6088 11452 6152 11456
rect 6088 11396 6092 11452
rect 6092 11396 6148 11452
rect 6148 11396 6152 11452
rect 6088 11392 6152 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 9272 11452 9336 11456
rect 9272 11396 9276 11452
rect 9276 11396 9332 11452
rect 9332 11396 9336 11452
rect 9272 11392 9336 11396
rect 9352 11452 9416 11456
rect 9352 11396 9356 11452
rect 9356 11396 9412 11452
rect 9412 11396 9416 11452
rect 9352 11392 9416 11396
rect 3372 11052 3436 11116
rect 3924 11112 3988 11116
rect 3924 11056 3974 11112
rect 3974 11056 3988 11112
rect 3924 11052 3988 11056
rect 5212 10976 5276 10980
rect 5212 10920 5262 10976
rect 5262 10920 5276 10976
rect 5212 10916 5276 10920
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 7480 10908 7544 10912
rect 7480 10852 7484 10908
rect 7484 10852 7540 10908
rect 7540 10852 7544 10908
rect 7480 10848 7544 10852
rect 7560 10908 7624 10912
rect 7560 10852 7564 10908
rect 7564 10852 7620 10908
rect 7620 10852 7624 10908
rect 7560 10848 7624 10852
rect 7640 10908 7704 10912
rect 7640 10852 7644 10908
rect 7644 10852 7700 10908
rect 7700 10852 7704 10908
rect 7640 10848 7704 10852
rect 7720 10908 7784 10912
rect 7720 10852 7724 10908
rect 7724 10852 7780 10908
rect 7780 10852 7784 10908
rect 7720 10848 7784 10852
rect 4660 10372 4724 10436
rect 2584 10364 2648 10368
rect 2584 10308 2588 10364
rect 2588 10308 2644 10364
rect 2644 10308 2648 10364
rect 2584 10304 2648 10308
rect 2664 10364 2728 10368
rect 2664 10308 2668 10364
rect 2668 10308 2724 10364
rect 2724 10308 2728 10364
rect 2664 10304 2728 10308
rect 2744 10364 2808 10368
rect 2744 10308 2748 10364
rect 2748 10308 2804 10364
rect 2804 10308 2808 10364
rect 2744 10304 2808 10308
rect 2824 10364 2888 10368
rect 2824 10308 2828 10364
rect 2828 10308 2884 10364
rect 2884 10308 2888 10364
rect 2824 10304 2888 10308
rect 5848 10364 5912 10368
rect 5848 10308 5852 10364
rect 5852 10308 5908 10364
rect 5908 10308 5912 10364
rect 5848 10304 5912 10308
rect 5928 10364 5992 10368
rect 5928 10308 5932 10364
rect 5932 10308 5988 10364
rect 5988 10308 5992 10364
rect 5928 10304 5992 10308
rect 6008 10364 6072 10368
rect 6008 10308 6012 10364
rect 6012 10308 6068 10364
rect 6068 10308 6072 10364
rect 6008 10304 6072 10308
rect 6088 10364 6152 10368
rect 6088 10308 6092 10364
rect 6092 10308 6148 10364
rect 6148 10308 6152 10364
rect 6088 10304 6152 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 9272 10364 9336 10368
rect 9272 10308 9276 10364
rect 9276 10308 9332 10364
rect 9332 10308 9336 10364
rect 9272 10304 9336 10308
rect 9352 10364 9416 10368
rect 9352 10308 9356 10364
rect 9356 10308 9412 10364
rect 9412 10308 9416 10364
rect 9352 10304 9416 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 7480 9820 7544 9824
rect 7480 9764 7484 9820
rect 7484 9764 7540 9820
rect 7540 9764 7544 9820
rect 7480 9760 7544 9764
rect 7560 9820 7624 9824
rect 7560 9764 7564 9820
rect 7564 9764 7620 9820
rect 7620 9764 7624 9820
rect 7560 9760 7624 9764
rect 7640 9820 7704 9824
rect 7640 9764 7644 9820
rect 7644 9764 7700 9820
rect 7700 9764 7704 9820
rect 7640 9760 7704 9764
rect 7720 9820 7784 9824
rect 7720 9764 7724 9820
rect 7724 9764 7780 9820
rect 7780 9764 7784 9820
rect 7720 9760 7784 9764
rect 2584 9276 2648 9280
rect 2584 9220 2588 9276
rect 2588 9220 2644 9276
rect 2644 9220 2648 9276
rect 2584 9216 2648 9220
rect 2664 9276 2728 9280
rect 2664 9220 2668 9276
rect 2668 9220 2724 9276
rect 2724 9220 2728 9276
rect 2664 9216 2728 9220
rect 2744 9276 2808 9280
rect 2744 9220 2748 9276
rect 2748 9220 2804 9276
rect 2804 9220 2808 9276
rect 2744 9216 2808 9220
rect 2824 9276 2888 9280
rect 2824 9220 2828 9276
rect 2828 9220 2884 9276
rect 2884 9220 2888 9276
rect 2824 9216 2888 9220
rect 5848 9276 5912 9280
rect 5848 9220 5852 9276
rect 5852 9220 5908 9276
rect 5908 9220 5912 9276
rect 5848 9216 5912 9220
rect 5928 9276 5992 9280
rect 5928 9220 5932 9276
rect 5932 9220 5988 9276
rect 5988 9220 5992 9276
rect 5928 9216 5992 9220
rect 6008 9276 6072 9280
rect 6008 9220 6012 9276
rect 6012 9220 6068 9276
rect 6068 9220 6072 9276
rect 6008 9216 6072 9220
rect 6088 9276 6152 9280
rect 6088 9220 6092 9276
rect 6092 9220 6148 9276
rect 6148 9220 6152 9276
rect 6088 9216 6152 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 9272 9276 9336 9280
rect 9272 9220 9276 9276
rect 9276 9220 9332 9276
rect 9332 9220 9336 9276
rect 9272 9216 9336 9220
rect 9352 9276 9416 9280
rect 9352 9220 9356 9276
rect 9356 9220 9412 9276
rect 9412 9220 9416 9276
rect 9352 9216 9416 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 7480 8732 7544 8736
rect 7480 8676 7484 8732
rect 7484 8676 7540 8732
rect 7540 8676 7544 8732
rect 7480 8672 7544 8676
rect 7560 8732 7624 8736
rect 7560 8676 7564 8732
rect 7564 8676 7620 8732
rect 7620 8676 7624 8732
rect 7560 8672 7624 8676
rect 7640 8732 7704 8736
rect 7640 8676 7644 8732
rect 7644 8676 7700 8732
rect 7700 8676 7704 8732
rect 7640 8672 7704 8676
rect 7720 8732 7784 8736
rect 7720 8676 7724 8732
rect 7724 8676 7780 8732
rect 7780 8676 7784 8732
rect 7720 8672 7784 8676
rect 5396 8392 5460 8396
rect 5396 8336 5410 8392
rect 5410 8336 5460 8392
rect 5396 8332 5460 8336
rect 2584 8188 2648 8192
rect 2584 8132 2588 8188
rect 2588 8132 2644 8188
rect 2644 8132 2648 8188
rect 2584 8128 2648 8132
rect 2664 8188 2728 8192
rect 2664 8132 2668 8188
rect 2668 8132 2724 8188
rect 2724 8132 2728 8188
rect 2664 8128 2728 8132
rect 2744 8188 2808 8192
rect 2744 8132 2748 8188
rect 2748 8132 2804 8188
rect 2804 8132 2808 8188
rect 2744 8128 2808 8132
rect 2824 8188 2888 8192
rect 2824 8132 2828 8188
rect 2828 8132 2884 8188
rect 2884 8132 2888 8188
rect 2824 8128 2888 8132
rect 5848 8188 5912 8192
rect 5848 8132 5852 8188
rect 5852 8132 5908 8188
rect 5908 8132 5912 8188
rect 5848 8128 5912 8132
rect 5928 8188 5992 8192
rect 5928 8132 5932 8188
rect 5932 8132 5988 8188
rect 5988 8132 5992 8188
rect 5928 8128 5992 8132
rect 6008 8188 6072 8192
rect 6008 8132 6012 8188
rect 6012 8132 6068 8188
rect 6068 8132 6072 8188
rect 6008 8128 6072 8132
rect 6088 8188 6152 8192
rect 6088 8132 6092 8188
rect 6092 8132 6148 8188
rect 6148 8132 6152 8188
rect 6088 8128 6152 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 9272 8188 9336 8192
rect 9272 8132 9276 8188
rect 9276 8132 9332 8188
rect 9332 8132 9336 8188
rect 9272 8128 9336 8132
rect 9352 8188 9416 8192
rect 9352 8132 9356 8188
rect 9356 8132 9412 8188
rect 9412 8132 9416 8188
rect 9352 8128 9416 8132
rect 7052 8120 7116 8124
rect 7052 8064 7066 8120
rect 7066 8064 7116 8120
rect 7052 8060 7116 8064
rect 3924 7924 3988 7988
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 7480 7644 7544 7648
rect 7480 7588 7484 7644
rect 7484 7588 7540 7644
rect 7540 7588 7544 7644
rect 7480 7584 7544 7588
rect 7560 7644 7624 7648
rect 7560 7588 7564 7644
rect 7564 7588 7620 7644
rect 7620 7588 7624 7644
rect 7560 7584 7624 7588
rect 7640 7644 7704 7648
rect 7640 7588 7644 7644
rect 7644 7588 7700 7644
rect 7700 7588 7704 7644
rect 7640 7584 7704 7588
rect 7720 7644 7784 7648
rect 7720 7588 7724 7644
rect 7724 7588 7780 7644
rect 7780 7588 7784 7644
rect 7720 7584 7784 7588
rect 2584 7100 2648 7104
rect 2584 7044 2588 7100
rect 2588 7044 2644 7100
rect 2644 7044 2648 7100
rect 2584 7040 2648 7044
rect 2664 7100 2728 7104
rect 2664 7044 2668 7100
rect 2668 7044 2724 7100
rect 2724 7044 2728 7100
rect 2664 7040 2728 7044
rect 2744 7100 2808 7104
rect 2744 7044 2748 7100
rect 2748 7044 2804 7100
rect 2804 7044 2808 7100
rect 2744 7040 2808 7044
rect 2824 7100 2888 7104
rect 2824 7044 2828 7100
rect 2828 7044 2884 7100
rect 2884 7044 2888 7100
rect 2824 7040 2888 7044
rect 5848 7100 5912 7104
rect 5848 7044 5852 7100
rect 5852 7044 5908 7100
rect 5908 7044 5912 7100
rect 5848 7040 5912 7044
rect 5928 7100 5992 7104
rect 5928 7044 5932 7100
rect 5932 7044 5988 7100
rect 5988 7044 5992 7100
rect 5928 7040 5992 7044
rect 6008 7100 6072 7104
rect 6008 7044 6012 7100
rect 6012 7044 6068 7100
rect 6068 7044 6072 7100
rect 6008 7040 6072 7044
rect 6088 7100 6152 7104
rect 6088 7044 6092 7100
rect 6092 7044 6148 7100
rect 6148 7044 6152 7100
rect 6088 7040 6152 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 9272 7100 9336 7104
rect 9272 7044 9276 7100
rect 9276 7044 9332 7100
rect 9332 7044 9336 7100
rect 9272 7040 9336 7044
rect 9352 7100 9416 7104
rect 9352 7044 9356 7100
rect 9356 7044 9412 7100
rect 9412 7044 9416 7100
rect 9352 7040 9416 7044
rect 5212 6836 5276 6900
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 7480 6556 7544 6560
rect 7480 6500 7484 6556
rect 7484 6500 7540 6556
rect 7540 6500 7544 6556
rect 7480 6496 7544 6500
rect 7560 6556 7624 6560
rect 7560 6500 7564 6556
rect 7564 6500 7620 6556
rect 7620 6500 7624 6556
rect 7560 6496 7624 6500
rect 7640 6556 7704 6560
rect 7640 6500 7644 6556
rect 7644 6500 7700 6556
rect 7700 6500 7704 6556
rect 7640 6496 7704 6500
rect 7720 6556 7784 6560
rect 7720 6500 7724 6556
rect 7724 6500 7780 6556
rect 7780 6500 7784 6556
rect 7720 6496 7784 6500
rect 2584 6012 2648 6016
rect 2584 5956 2588 6012
rect 2588 5956 2644 6012
rect 2644 5956 2648 6012
rect 2584 5952 2648 5956
rect 2664 6012 2728 6016
rect 2664 5956 2668 6012
rect 2668 5956 2724 6012
rect 2724 5956 2728 6012
rect 2664 5952 2728 5956
rect 2744 6012 2808 6016
rect 2744 5956 2748 6012
rect 2748 5956 2804 6012
rect 2804 5956 2808 6012
rect 2744 5952 2808 5956
rect 2824 6012 2888 6016
rect 2824 5956 2828 6012
rect 2828 5956 2884 6012
rect 2884 5956 2888 6012
rect 2824 5952 2888 5956
rect 5848 6012 5912 6016
rect 5848 5956 5852 6012
rect 5852 5956 5908 6012
rect 5908 5956 5912 6012
rect 5848 5952 5912 5956
rect 5928 6012 5992 6016
rect 5928 5956 5932 6012
rect 5932 5956 5988 6012
rect 5988 5956 5992 6012
rect 5928 5952 5992 5956
rect 6008 6012 6072 6016
rect 6008 5956 6012 6012
rect 6012 5956 6068 6012
rect 6068 5956 6072 6012
rect 6008 5952 6072 5956
rect 6088 6012 6152 6016
rect 6088 5956 6092 6012
rect 6092 5956 6148 6012
rect 6148 5956 6152 6012
rect 6088 5952 6152 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 9272 6012 9336 6016
rect 9272 5956 9276 6012
rect 9276 5956 9332 6012
rect 9332 5956 9336 6012
rect 9272 5952 9336 5956
rect 9352 6012 9416 6016
rect 9352 5956 9356 6012
rect 9356 5956 9412 6012
rect 9412 5956 9416 6012
rect 9352 5952 9416 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 7480 5468 7544 5472
rect 7480 5412 7484 5468
rect 7484 5412 7540 5468
rect 7540 5412 7544 5468
rect 7480 5408 7544 5412
rect 7560 5468 7624 5472
rect 7560 5412 7564 5468
rect 7564 5412 7620 5468
rect 7620 5412 7624 5468
rect 7560 5408 7624 5412
rect 7640 5468 7704 5472
rect 7640 5412 7644 5468
rect 7644 5412 7700 5468
rect 7700 5412 7704 5468
rect 7640 5408 7704 5412
rect 7720 5468 7784 5472
rect 7720 5412 7724 5468
rect 7724 5412 7780 5468
rect 7780 5412 7784 5468
rect 7720 5408 7784 5412
rect 2584 4924 2648 4928
rect 2584 4868 2588 4924
rect 2588 4868 2644 4924
rect 2644 4868 2648 4924
rect 2584 4864 2648 4868
rect 2664 4924 2728 4928
rect 2664 4868 2668 4924
rect 2668 4868 2724 4924
rect 2724 4868 2728 4924
rect 2664 4864 2728 4868
rect 2744 4924 2808 4928
rect 2744 4868 2748 4924
rect 2748 4868 2804 4924
rect 2804 4868 2808 4924
rect 2744 4864 2808 4868
rect 2824 4924 2888 4928
rect 2824 4868 2828 4924
rect 2828 4868 2884 4924
rect 2884 4868 2888 4924
rect 2824 4864 2888 4868
rect 5848 4924 5912 4928
rect 5848 4868 5852 4924
rect 5852 4868 5908 4924
rect 5908 4868 5912 4924
rect 5848 4864 5912 4868
rect 5928 4924 5992 4928
rect 5928 4868 5932 4924
rect 5932 4868 5988 4924
rect 5988 4868 5992 4924
rect 5928 4864 5992 4868
rect 6008 4924 6072 4928
rect 6008 4868 6012 4924
rect 6012 4868 6068 4924
rect 6068 4868 6072 4924
rect 6008 4864 6072 4868
rect 6088 4924 6152 4928
rect 6088 4868 6092 4924
rect 6092 4868 6148 4924
rect 6148 4868 6152 4924
rect 6088 4864 6152 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 9272 4924 9336 4928
rect 9272 4868 9276 4924
rect 9276 4868 9332 4924
rect 9332 4868 9336 4924
rect 9272 4864 9336 4868
rect 9352 4924 9416 4928
rect 9352 4868 9356 4924
rect 9356 4868 9412 4924
rect 9412 4868 9416 4924
rect 9352 4864 9416 4868
rect 5212 4524 5276 4588
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 7480 4380 7544 4384
rect 7480 4324 7484 4380
rect 7484 4324 7540 4380
rect 7540 4324 7544 4380
rect 7480 4320 7544 4324
rect 7560 4380 7624 4384
rect 7560 4324 7564 4380
rect 7564 4324 7620 4380
rect 7620 4324 7624 4380
rect 7560 4320 7624 4324
rect 7640 4380 7704 4384
rect 7640 4324 7644 4380
rect 7644 4324 7700 4380
rect 7700 4324 7704 4380
rect 7640 4320 7704 4324
rect 7720 4380 7784 4384
rect 7720 4324 7724 4380
rect 7724 4324 7780 4380
rect 7780 4324 7784 4380
rect 7720 4320 7784 4324
rect 5396 3980 5460 4044
rect 2584 3836 2648 3840
rect 2584 3780 2588 3836
rect 2588 3780 2644 3836
rect 2644 3780 2648 3836
rect 2584 3776 2648 3780
rect 2664 3836 2728 3840
rect 2664 3780 2668 3836
rect 2668 3780 2724 3836
rect 2724 3780 2728 3836
rect 2664 3776 2728 3780
rect 2744 3836 2808 3840
rect 2744 3780 2748 3836
rect 2748 3780 2804 3836
rect 2804 3780 2808 3836
rect 2744 3776 2808 3780
rect 2824 3836 2888 3840
rect 2824 3780 2828 3836
rect 2828 3780 2884 3836
rect 2884 3780 2888 3836
rect 2824 3776 2888 3780
rect 5848 3836 5912 3840
rect 5848 3780 5852 3836
rect 5852 3780 5908 3836
rect 5908 3780 5912 3836
rect 5848 3776 5912 3780
rect 5928 3836 5992 3840
rect 5928 3780 5932 3836
rect 5932 3780 5988 3836
rect 5988 3780 5992 3836
rect 5928 3776 5992 3780
rect 6008 3836 6072 3840
rect 6008 3780 6012 3836
rect 6012 3780 6068 3836
rect 6068 3780 6072 3836
rect 6008 3776 6072 3780
rect 6088 3836 6152 3840
rect 6088 3780 6092 3836
rect 6092 3780 6148 3836
rect 6148 3780 6152 3836
rect 6088 3776 6152 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 9272 3836 9336 3840
rect 9272 3780 9276 3836
rect 9276 3780 9332 3836
rect 9332 3780 9336 3836
rect 9272 3776 9336 3780
rect 9352 3836 9416 3840
rect 9352 3780 9356 3836
rect 9356 3780 9412 3836
rect 9412 3780 9416 3836
rect 9352 3776 9416 3780
rect 4660 3708 4724 3772
rect 7052 3496 7116 3500
rect 7052 3440 7066 3496
rect 7066 3440 7116 3496
rect 7052 3436 7116 3440
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 7480 3292 7544 3296
rect 7480 3236 7484 3292
rect 7484 3236 7540 3292
rect 7540 3236 7544 3292
rect 7480 3232 7544 3236
rect 7560 3292 7624 3296
rect 7560 3236 7564 3292
rect 7564 3236 7620 3292
rect 7620 3236 7624 3292
rect 7560 3232 7624 3236
rect 7640 3292 7704 3296
rect 7640 3236 7644 3292
rect 7644 3236 7700 3292
rect 7700 3236 7704 3292
rect 7640 3232 7704 3236
rect 7720 3292 7784 3296
rect 7720 3236 7724 3292
rect 7724 3236 7780 3292
rect 7780 3236 7784 3292
rect 7720 3232 7784 3236
rect 5212 2816 5276 2820
rect 5212 2760 5262 2816
rect 5262 2760 5276 2816
rect 5212 2756 5276 2760
rect 2584 2748 2648 2752
rect 2584 2692 2588 2748
rect 2588 2692 2644 2748
rect 2644 2692 2648 2748
rect 2584 2688 2648 2692
rect 2664 2748 2728 2752
rect 2664 2692 2668 2748
rect 2668 2692 2724 2748
rect 2724 2692 2728 2748
rect 2664 2688 2728 2692
rect 2744 2748 2808 2752
rect 2744 2692 2748 2748
rect 2748 2692 2804 2748
rect 2804 2692 2808 2748
rect 2744 2688 2808 2692
rect 2824 2748 2888 2752
rect 2824 2692 2828 2748
rect 2828 2692 2884 2748
rect 2884 2692 2888 2748
rect 2824 2688 2888 2692
rect 5848 2748 5912 2752
rect 5848 2692 5852 2748
rect 5852 2692 5908 2748
rect 5908 2692 5912 2748
rect 5848 2688 5912 2692
rect 5928 2748 5992 2752
rect 5928 2692 5932 2748
rect 5932 2692 5988 2748
rect 5988 2692 5992 2748
rect 5928 2688 5992 2692
rect 6008 2748 6072 2752
rect 6008 2692 6012 2748
rect 6012 2692 6068 2748
rect 6068 2692 6072 2748
rect 6008 2688 6072 2692
rect 6088 2748 6152 2752
rect 6088 2692 6092 2748
rect 6092 2692 6148 2748
rect 6148 2692 6152 2748
rect 6088 2688 6152 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 9272 2748 9336 2752
rect 9272 2692 9276 2748
rect 9276 2692 9332 2748
rect 9332 2692 9336 2748
rect 9272 2688 9336 2692
rect 9352 2748 9416 2752
rect 9352 2692 9356 2748
rect 9356 2692 9412 2748
rect 9412 2692 9416 2748
rect 9352 2688 9416 2692
rect 3372 2620 3436 2684
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 7480 2204 7544 2208
rect 7480 2148 7484 2204
rect 7484 2148 7540 2204
rect 7540 2148 7544 2204
rect 7480 2144 7544 2148
rect 7560 2204 7624 2208
rect 7560 2148 7564 2204
rect 7564 2148 7620 2204
rect 7620 2148 7624 2204
rect 7560 2144 7624 2148
rect 7640 2204 7704 2208
rect 7640 2148 7644 2204
rect 7644 2148 7700 2204
rect 7700 2148 7704 2204
rect 7640 2144 7704 2148
rect 7720 2204 7784 2208
rect 7720 2148 7724 2204
rect 7724 2148 7780 2204
rect 7780 2148 7784 2204
rect 7720 2144 7784 2148
<< metal4 >>
rect 2576 11456 2896 11472
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 10368 2896 11392
rect 3371 11116 3437 11117
rect 3371 11052 3372 11116
rect 3436 11052 3437 11116
rect 3371 11051 3437 11052
rect 3923 11116 3989 11117
rect 3923 11052 3924 11116
rect 3988 11052 3989 11116
rect 3923 11051 3989 11052
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 9280 2896 10304
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 8192 2896 9216
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 7104 2896 8128
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2576 6016 2896 7040
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 4928 2896 5952
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 3840 2896 4864
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 2752 2896 3776
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2128 2896 2688
rect 3374 2685 3434 11051
rect 3926 7989 3986 11051
rect 4208 10912 4528 11472
rect 5840 11456 6160 11472
rect 5840 11392 5848 11456
rect 5912 11392 5928 11456
rect 5992 11392 6008 11456
rect 6072 11392 6088 11456
rect 6152 11392 6160 11456
rect 5211 10980 5277 10981
rect 5211 10916 5212 10980
rect 5276 10916 5277 10980
rect 5211 10915 5277 10916
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4659 10436 4725 10437
rect 4659 10372 4660 10436
rect 4724 10372 4725 10436
rect 4659 10371 4725 10372
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 3923 7988 3989 7989
rect 3923 7924 3924 7988
rect 3988 7924 3989 7988
rect 3923 7923 3989 7924
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4662 3773 4722 10371
rect 5214 6901 5274 10915
rect 5840 10368 6160 11392
rect 5840 10304 5848 10368
rect 5912 10304 5928 10368
rect 5992 10304 6008 10368
rect 6072 10304 6088 10368
rect 6152 10304 6160 10368
rect 5840 9280 6160 10304
rect 5840 9216 5848 9280
rect 5912 9216 5928 9280
rect 5992 9216 6008 9280
rect 6072 9216 6088 9280
rect 6152 9216 6160 9280
rect 5395 8396 5461 8397
rect 5395 8332 5396 8396
rect 5460 8332 5461 8396
rect 5395 8331 5461 8332
rect 5211 6900 5277 6901
rect 5211 6836 5212 6900
rect 5276 6836 5277 6900
rect 5211 6835 5277 6836
rect 5211 4588 5277 4589
rect 5211 4524 5212 4588
rect 5276 4524 5277 4588
rect 5211 4523 5277 4524
rect 4659 3772 4725 3773
rect 4659 3708 4660 3772
rect 4724 3708 4725 3772
rect 4659 3707 4725 3708
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 3371 2684 3437 2685
rect 3371 2620 3372 2684
rect 3436 2620 3437 2684
rect 3371 2619 3437 2620
rect 4208 2208 4528 3232
rect 5214 2821 5274 4523
rect 5398 4045 5458 8331
rect 5840 8192 6160 9216
rect 5840 8128 5848 8192
rect 5912 8128 5928 8192
rect 5992 8128 6008 8192
rect 6072 8128 6088 8192
rect 6152 8128 6160 8192
rect 5840 7104 6160 8128
rect 7472 10912 7792 11472
rect 7472 10848 7480 10912
rect 7544 10848 7560 10912
rect 7624 10848 7640 10912
rect 7704 10848 7720 10912
rect 7784 10848 7792 10912
rect 7472 9824 7792 10848
rect 7472 9760 7480 9824
rect 7544 9760 7560 9824
rect 7624 9760 7640 9824
rect 7704 9760 7720 9824
rect 7784 9760 7792 9824
rect 7472 8736 7792 9760
rect 7472 8672 7480 8736
rect 7544 8672 7560 8736
rect 7624 8672 7640 8736
rect 7704 8672 7720 8736
rect 7784 8672 7792 8736
rect 7051 8124 7117 8125
rect 7051 8060 7052 8124
rect 7116 8060 7117 8124
rect 7051 8059 7117 8060
rect 5840 7040 5848 7104
rect 5912 7040 5928 7104
rect 5992 7040 6008 7104
rect 6072 7040 6088 7104
rect 6152 7040 6160 7104
rect 5840 6016 6160 7040
rect 5840 5952 5848 6016
rect 5912 5952 5928 6016
rect 5992 5952 6008 6016
rect 6072 5952 6088 6016
rect 6152 5952 6160 6016
rect 5840 4928 6160 5952
rect 5840 4864 5848 4928
rect 5912 4864 5928 4928
rect 5992 4864 6008 4928
rect 6072 4864 6088 4928
rect 6152 4864 6160 4928
rect 5395 4044 5461 4045
rect 5395 3980 5396 4044
rect 5460 3980 5461 4044
rect 5395 3979 5461 3980
rect 5840 3840 6160 4864
rect 5840 3776 5848 3840
rect 5912 3776 5928 3840
rect 5992 3776 6008 3840
rect 6072 3776 6088 3840
rect 6152 3776 6160 3840
rect 5211 2820 5277 2821
rect 5211 2756 5212 2820
rect 5276 2756 5277 2820
rect 5211 2755 5277 2756
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 5840 2752 6160 3776
rect 7054 3501 7114 8059
rect 7472 7648 7792 8672
rect 7472 7584 7480 7648
rect 7544 7584 7560 7648
rect 7624 7584 7640 7648
rect 7704 7584 7720 7648
rect 7784 7584 7792 7648
rect 7472 6560 7792 7584
rect 7472 6496 7480 6560
rect 7544 6496 7560 6560
rect 7624 6496 7640 6560
rect 7704 6496 7720 6560
rect 7784 6496 7792 6560
rect 7472 5472 7792 6496
rect 7472 5408 7480 5472
rect 7544 5408 7560 5472
rect 7624 5408 7640 5472
rect 7704 5408 7720 5472
rect 7784 5408 7792 5472
rect 7472 4384 7792 5408
rect 7472 4320 7480 4384
rect 7544 4320 7560 4384
rect 7624 4320 7640 4384
rect 7704 4320 7720 4384
rect 7784 4320 7792 4384
rect 7051 3500 7117 3501
rect 7051 3436 7052 3500
rect 7116 3436 7117 3500
rect 7051 3435 7117 3436
rect 5840 2688 5848 2752
rect 5912 2688 5928 2752
rect 5992 2688 6008 2752
rect 6072 2688 6088 2752
rect 6152 2688 6160 2752
rect 5840 2128 6160 2688
rect 7472 3296 7792 4320
rect 7472 3232 7480 3296
rect 7544 3232 7560 3296
rect 7624 3232 7640 3296
rect 7704 3232 7720 3296
rect 7784 3232 7792 3296
rect 7472 2208 7792 3232
rect 7472 2144 7480 2208
rect 7544 2144 7560 2208
rect 7624 2144 7640 2208
rect 7704 2144 7720 2208
rect 7784 2144 7792 2208
rect 7472 2128 7792 2144
rect 9104 11456 9424 11472
rect 9104 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9272 11456
rect 9336 11392 9352 11456
rect 9416 11392 9424 11456
rect 9104 10368 9424 11392
rect 9104 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9272 10368
rect 9336 10304 9352 10368
rect 9416 10304 9424 10368
rect 9104 9280 9424 10304
rect 9104 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9272 9280
rect 9336 9216 9352 9280
rect 9416 9216 9424 9280
rect 9104 8192 9424 9216
rect 9104 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9272 8192
rect 9336 8128 9352 8192
rect 9416 8128 9424 8192
rect 9104 7104 9424 8128
rect 9104 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9272 7104
rect 9336 7040 9352 7104
rect 9416 7040 9424 7104
rect 9104 6016 9424 7040
rect 9104 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9272 6016
rect 9336 5952 9352 6016
rect 9416 5952 9424 6016
rect 9104 4928 9424 5952
rect 9104 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9272 4928
rect 9336 4864 9352 4928
rect 9416 4864 9424 4928
rect 9104 3840 9424 4864
rect 9104 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9272 3840
rect 9336 3776 9352 3840
rect 9416 3776 9424 3840
rect 9104 2752 9424 3776
rect 9104 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9272 2752
rect 9336 2688 9352 2752
rect 9416 2688 9424 2752
rect 9104 2128 9424 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46
timestamp 1644511149
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1644511149
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1644511149
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_33
timestamp 1644511149
transform 1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_42
timestamp 1644511149
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_67
timestamp 1644511149
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1644511149
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1644511149
transform 1 0 8648 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_94
timestamp 1644511149
transform 1 0 9752 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_102
timestamp 1644511149
transform 1 0 10488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1644511149
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_39
timestamp 1644511149
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1644511149
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1644511149
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_71
timestamp 1644511149
transform 1 0 7636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1644511149
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_88
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_100
timestamp 1644511149
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_12
timestamp 1644511149
transform 1 0 2208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_21
timestamp 1644511149
transform 1 0 3036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_32
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_70
timestamp 1644511149
transform 1 0 7544 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_79
timestamp 1644511149
transform 1 0 8372 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_87
timestamp 1644511149
transform 1 0 9108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1644511149
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_8
timestamp 1644511149
transform 1 0 1840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_16
timestamp 1644511149
transform 1 0 2576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1644511149
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_50
timestamp 1644511149
transform 1 0 5704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_56
timestamp 1644511149
transform 1 0 6256 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_73
timestamp 1644511149
transform 1 0 7820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1644511149
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1644511149
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_98
timestamp 1644511149
transform 1 0 10120 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_102
timestamp 1644511149
transform 1 0 10488 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1644511149
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_18
timestamp 1644511149
transform 1 0 2760 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_29
timestamp 1644511149
transform 1 0 3772 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_73
timestamp 1644511149
transform 1 0 7820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_84
timestamp 1644511149
transform 1 0 8832 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1644511149
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1644511149
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp 1644511149
transform 1 0 4324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1644511149
transform 1 0 5888 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_56
timestamp 1644511149
transform 1 0 6256 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_73
timestamp 1644511149
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1644511149
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_92
timestamp 1644511149
transform 1 0 9568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1644511149
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1644511149
transform 1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_32
timestamp 1644511149
transform 1 0 4048 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1644511149
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1644511149
transform 1 0 7912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_94
timestamp 1644511149
transform 1 0 9752 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_102
timestamp 1644511149
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1644511149
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1644511149
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_42
timestamp 1644511149
transform 1 0 4968 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_50
timestamp 1644511149
transform 1 0 5704 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_71
timestamp 1644511149
transform 1 0 7636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_75
timestamp 1644511149
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1644511149
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_92
timestamp 1644511149
transform 1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1644511149
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1644511149
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_73
timestamp 1644511149
transform 1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1644511149
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_10
timestamp 1644511149
transform 1 0 2024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1644511149
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1644511149
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1644511149
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_95
timestamp 1644511149
transform 1 0 9844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_12
timestamp 1644511149
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_26
timestamp 1644511149
transform 1 0 3496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_46
timestamp 1644511149
transform 1 0 5336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1644511149
transform 1 0 7820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1644511149
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_38
timestamp 1644511149
transform 1 0 4600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1644511149
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_78
timestamp 1644511149
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_92
timestamp 1644511149
transform 1 0 9568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1644511149
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_7
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_14
timestamp 1644511149
transform 1 0 2392 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_22
timestamp 1644511149
transform 1 0 3128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_32
timestamp 1644511149
transform 1 0 4048 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1644511149
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_73
timestamp 1644511149
transform 1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_84
timestamp 1644511149
transform 1 0 8832 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1644511149
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_10
timestamp 1644511149
transform 1 0 2024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_17
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1644511149
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 1644511149
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 1644511149
transform 1 0 6716 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_72
timestamp 1644511149
transform 1 0 7728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1644511149
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1644511149
transform 1 0 9200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_95
timestamp 1644511149
transform 1 0 9844 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1644511149
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_20
timestamp 1644511149
transform 1 0 2944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_35
timestamp 1644511149
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_46
timestamp 1644511149
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1644511149
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_64
timestamp 1644511149
transform 1 0 6992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_73
timestamp 1644511149
transform 1 0 7820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_88
timestamp 1644511149
transform 1 0 9200 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_100
timestamp 1644511149
transform 1 0 10304 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_5
timestamp 1644511149
transform 1 0 1564 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_17
timestamp 1644511149
transform 1 0 2668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1644511149
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1644511149
transform 1 0 4048 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_39
timestamp 1644511149
transform 1 0 4692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_48
timestamp 1644511149
transform 1 0 5520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_62
timestamp 1644511149
transform 1 0 6808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_71
timestamp 1644511149
transform 1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_78
timestamp 1644511149
transform 1 0 8280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1644511149
transform 1 0 6256 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__and4_1  _088_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4600 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _089_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4232 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _090_
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _091_
timestamp 1644511149
transform 1 0 4232 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _092_
timestamp 1644511149
transform -1 0 5704 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _093_
timestamp 1644511149
transform -1 0 9660 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _094_
timestamp 1644511149
transform -1 0 8372 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _095_
timestamp 1644511149
transform 1 0 8188 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _096_
timestamp 1644511149
transform -1 0 6808 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _097_
timestamp 1644511149
transform -1 0 6992 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _098_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _099_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _100_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3312 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _101_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7728 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _102_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _103_
timestamp 1644511149
transform 1 0 2576 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _104_
timestamp 1644511149
transform -1 0 4692 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _105_
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _106_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _107_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _108_
timestamp 1644511149
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _109_
timestamp 1644511149
transform -1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _110_
timestamp 1644511149
transform 1 0 4232 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _111_
timestamp 1644511149
transform -1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1644511149
transform -1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _113_
timestamp 1644511149
transform -1 0 2024 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1644511149
transform -1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _115_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1644511149
transform -1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _117_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2208 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _118_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _119_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5060 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1644511149
transform 1 0 9936 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1644511149
transform -1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _122_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _123_
timestamp 1644511149
transform 1 0 2300 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _124_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3496 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1644511149
transform -1 0 2944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _126_
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1644511149
transform -1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1644511149
transform -1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1644511149
transform -1 0 8648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _130_
timestamp 1644511149
transform -1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _131_
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _132_
timestamp 1644511149
transform -1 0 2300 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _133_
timestamp 1644511149
transform 1 0 2208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _134_
timestamp 1644511149
transform -1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _135_
timestamp 1644511149
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _136_
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _137_
timestamp 1644511149
transform 1 0 4508 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _138_
timestamp 1644511149
transform -1 0 3772 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _139_
timestamp 1644511149
transform 1 0 3404 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _141_
timestamp 1644511149
transform -1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _142_
timestamp 1644511149
transform -1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _143_
timestamp 1644511149
transform -1 0 8372 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _144_
timestamp 1644511149
transform -1 0 7544 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _145_
timestamp 1644511149
transform -1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _146_
timestamp 1644511149
transform -1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _147_
timestamp 1644511149
transform -1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _148_
timestamp 1644511149
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _149_
timestamp 1644511149
transform 1 0 8740 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _150_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _151_
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _152_
timestamp 1644511149
transform 1 0 1564 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _154_
timestamp 1644511149
transform -1 0 5796 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _155_
timestamp 1644511149
transform -1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _156_
timestamp 1644511149
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _157_
timestamp 1644511149
transform 1 0 2576 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _158_
timestamp 1644511149
transform -1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _159_
timestamp 1644511149
transform -1 0 3312 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _160_
timestamp 1644511149
transform -1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _161_
timestamp 1644511149
transform -1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _162_
timestamp 1644511149
transform 1 0 7360 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _163_
timestamp 1644511149
transform -1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _164_
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _165_
timestamp 1644511149
transform 1 0 9200 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _166_
timestamp 1644511149
transform -1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _167_
timestamp 1644511149
transform 1 0 7176 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1644511149
transform 1 0 8924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1644511149
transform 1 0 9568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _170_
timestamp 1644511149
transform -1 0 9568 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _171_
timestamp 1644511149
transform 1 0 8188 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _172_
timestamp 1644511149
transform 1 0 6072 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1644511149
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _174_
timestamp 1644511149
transform -1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _175_
timestamp 1644511149
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _176_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 5520 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _177_
timestamp 1644511149
transform 1 0 3956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _178_
timestamp 1644511149
transform 1 0 3864 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _179_
timestamp 1644511149
transform -1 0 7360 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _180_
timestamp 1644511149
transform -1 0 5888 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _181_
timestamp 1644511149
transform -1 0 5888 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _182_
timestamp 1644511149
transform 1 0 4140 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _183_
timestamp 1644511149
transform 1 0 6440 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _184_
timestamp 1644511149
transform 1 0 4232 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _185_
timestamp 1644511149
transform -1 0 4048 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _186_
timestamp 1644511149
transform -1 0 7820 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _187_
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _188_
timestamp 1644511149
transform 1 0 4416 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _189_
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _190_
timestamp 1644511149
transform 1 0 4968 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _191_
timestamp 1644511149
transform 1 0 6348 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _192_
timestamp 1644511149
transform 1 0 1840 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _193_
timestamp 1644511149
transform -1 0 3588 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _194_
timestamp 1644511149
transform 1 0 4416 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _195_
timestamp 1644511149
transform -1 0 7820 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _196_
timestamp 1644511149
transform -1 0 8280 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _197_
timestamp 1644511149
transform 1 0 5244 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _198_
timestamp 1644511149
transform -1 0 9660 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _199_
timestamp 1644511149
transform -1 0 7820 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _200_
timestamp 1644511149
transform 1 0 8280 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _201_
timestamp 1644511149
transform -1 0 9660 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5796 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4968 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 1644511149
transform 1 0 8096 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output2 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9844 0 -1 4352
box -38 -48 406 592
<< labels >>
rlabel metal3 s 11200 6944 12000 7064 6 blink
port 0 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 clk
port 1 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 nrst
port 2 nsew signal input
rlabel metal4 s 2576 2128 2896 11472 6 vccd1
port 3 nsew power input
rlabel metal4 s 5840 2128 6160 11472 6 vccd1
port 3 nsew power input
rlabel metal4 s 9104 2128 9424 11472 6 vccd1
port 3 nsew power input
rlabel metal4 s 4208 2128 4528 11472 6 vssd1
port 4 nsew ground input
rlabel metal4 s 7472 2128 7792 11472 6 vssd1
port 4 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 12000 14000
<< end >>
