VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ExperiarCore
  CLASS BLOCK ;
  FOREIGN ExperiarCore ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 1000.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END addr0[8]
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.880 4.000 655.480 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END addr1[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END clk0
  PIN clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END clk1
  PIN coreIndex[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 996.000 6.350 1000.000 ;
    END
  END coreIndex[0]
  PIN coreIndex[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 996.000 18.770 1000.000 ;
    END
  END coreIndex[1]
  PIN coreIndex[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 996.000 31.650 1000.000 ;
    END
  END coreIndex[2]
  PIN coreIndex[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 996.000 44.530 1000.000 ;
    END
  END coreIndex[3]
  PIN coreIndex[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 996.000 57.410 1000.000 ;
    END
  END coreIndex[4]
  PIN coreIndex[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 996.000 70.290 1000.000 ;
    END
  END coreIndex[5]
  PIN coreIndex[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 996.000 83.170 1000.000 ;
    END
  END coreIndex[6]
  PIN coreIndex[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 996.000 96.050 1000.000 ;
    END
  END coreIndex[7]
  PIN core_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 11.600 500.000 12.200 ;
    END
  END core_wb_ack_i
  PIN core_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 41.520 500.000 42.120 ;
    END
  END core_wb_adr_o[0]
  PIN core_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 209.480 500.000 210.080 ;
    END
  END core_wb_adr_o[10]
  PIN core_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 224.440 500.000 225.040 ;
    END
  END core_wb_adr_o[11]
  PIN core_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 239.400 500.000 240.000 ;
    END
  END core_wb_adr_o[12]
  PIN core_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 254.360 500.000 254.960 ;
    END
  END core_wb_adr_o[13]
  PIN core_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 269.320 500.000 269.920 ;
    END
  END core_wb_adr_o[14]
  PIN core_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 284.280 500.000 284.880 ;
    END
  END core_wb_adr_o[15]
  PIN core_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 298.560 500.000 299.160 ;
    END
  END core_wb_adr_o[16]
  PIN core_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 313.520 500.000 314.120 ;
    END
  END core_wb_adr_o[17]
  PIN core_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 328.480 500.000 329.080 ;
    END
  END core_wb_adr_o[18]
  PIN core_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 343.440 500.000 344.040 ;
    END
  END core_wb_adr_o[19]
  PIN core_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 61.240 500.000 61.840 ;
    END
  END core_wb_adr_o[1]
  PIN core_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 358.400 500.000 359.000 ;
    END
  END core_wb_adr_o[20]
  PIN core_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 373.360 500.000 373.960 ;
    END
  END core_wb_adr_o[21]
  PIN core_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 388.320 500.000 388.920 ;
    END
  END core_wb_adr_o[22]
  PIN core_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 402.600 500.000 403.200 ;
    END
  END core_wb_adr_o[23]
  PIN core_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 417.560 500.000 418.160 ;
    END
  END core_wb_adr_o[24]
  PIN core_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 432.520 500.000 433.120 ;
    END
  END core_wb_adr_o[25]
  PIN core_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 447.480 500.000 448.080 ;
    END
  END core_wb_adr_o[26]
  PIN core_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 462.440 500.000 463.040 ;
    END
  END core_wb_adr_o[27]
  PIN core_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 80.960 500.000 81.560 ;
    END
  END core_wb_adr_o[2]
  PIN core_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 100.680 500.000 101.280 ;
    END
  END core_wb_adr_o[3]
  PIN core_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 120.400 500.000 121.000 ;
    END
  END core_wb_adr_o[4]
  PIN core_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 135.360 500.000 135.960 ;
    END
  END core_wb_adr_o[5]
  PIN core_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 150.320 500.000 150.920 ;
    END
  END core_wb_adr_o[6]
  PIN core_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 165.280 500.000 165.880 ;
    END
  END core_wb_adr_o[7]
  PIN core_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 180.240 500.000 180.840 ;
    END
  END core_wb_adr_o[8]
  PIN core_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 195.200 500.000 195.800 ;
    END
  END core_wb_adr_o[9]
  PIN core_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 16.360 500.000 16.960 ;
    END
  END core_wb_cyc_o
  PIN core_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 46.280 500.000 46.880 ;
    END
  END core_wb_data_i[0]
  PIN core_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 214.920 500.000 215.520 ;
    END
  END core_wb_data_i[10]
  PIN core_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 229.200 500.000 229.800 ;
    END
  END core_wb_data_i[11]
  PIN core_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 244.160 500.000 244.760 ;
    END
  END core_wb_data_i[12]
  PIN core_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 259.120 500.000 259.720 ;
    END
  END core_wb_data_i[13]
  PIN core_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 274.080 500.000 274.680 ;
    END
  END core_wb_data_i[14]
  PIN core_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 289.040 500.000 289.640 ;
    END
  END core_wb_data_i[15]
  PIN core_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 304.000 500.000 304.600 ;
    END
  END core_wb_data_i[16]
  PIN core_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 318.960 500.000 319.560 ;
    END
  END core_wb_data_i[17]
  PIN core_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 333.240 500.000 333.840 ;
    END
  END core_wb_data_i[18]
  PIN core_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 348.200 500.000 348.800 ;
    END
  END core_wb_data_i[19]
  PIN core_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 66.000 500.000 66.600 ;
    END
  END core_wb_data_i[1]
  PIN core_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 363.160 500.000 363.760 ;
    END
  END core_wb_data_i[20]
  PIN core_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 378.120 500.000 378.720 ;
    END
  END core_wb_data_i[21]
  PIN core_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 393.080 500.000 393.680 ;
    END
  END core_wb_data_i[22]
  PIN core_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 408.040 500.000 408.640 ;
    END
  END core_wb_data_i[23]
  PIN core_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 422.320 500.000 422.920 ;
    END
  END core_wb_data_i[24]
  PIN core_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 437.280 500.000 437.880 ;
    END
  END core_wb_data_i[25]
  PIN core_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 452.240 500.000 452.840 ;
    END
  END core_wb_data_i[26]
  PIN core_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 467.200 500.000 467.800 ;
    END
  END core_wb_data_i[27]
  PIN core_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 477.400 500.000 478.000 ;
    END
  END core_wb_data_i[28]
  PIN core_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 486.920 500.000 487.520 ;
    END
  END core_wb_data_i[29]
  PIN core_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 85.720 500.000 86.320 ;
    END
  END core_wb_data_i[2]
  PIN core_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 497.120 500.000 497.720 ;
    END
  END core_wb_data_i[30]
  PIN core_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 506.640 500.000 507.240 ;
    END
  END core_wb_data_i[31]
  PIN core_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 105.440 500.000 106.040 ;
    END
  END core_wb_data_i[3]
  PIN core_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 125.840 500.000 126.440 ;
    END
  END core_wb_data_i[4]
  PIN core_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 140.120 500.000 140.720 ;
    END
  END core_wb_data_i[5]
  PIN core_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 155.080 500.000 155.680 ;
    END
  END core_wb_data_i[6]
  PIN core_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 170.040 500.000 170.640 ;
    END
  END core_wb_data_i[7]
  PIN core_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 185.000 500.000 185.600 ;
    END
  END core_wb_data_i[8]
  PIN core_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 199.960 500.000 200.560 ;
    END
  END core_wb_data_i[9]
  PIN core_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 51.040 500.000 51.640 ;
    END
  END core_wb_data_o[0]
  PIN core_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 219.680 500.000 220.280 ;
    END
  END core_wb_data_o[10]
  PIN core_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 234.640 500.000 235.240 ;
    END
  END core_wb_data_o[11]
  PIN core_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 249.600 500.000 250.200 ;
    END
  END core_wb_data_o[12]
  PIN core_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 263.880 500.000 264.480 ;
    END
  END core_wb_data_o[13]
  PIN core_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 278.840 500.000 279.440 ;
    END
  END core_wb_data_o[14]
  PIN core_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 293.800 500.000 294.400 ;
    END
  END core_wb_data_o[15]
  PIN core_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 308.760 500.000 309.360 ;
    END
  END core_wb_data_o[16]
  PIN core_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 323.720 500.000 324.320 ;
    END
  END core_wb_data_o[17]
  PIN core_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 338.680 500.000 339.280 ;
    END
  END core_wb_data_o[18]
  PIN core_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 353.640 500.000 354.240 ;
    END
  END core_wb_data_o[19]
  PIN core_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 70.760 500.000 71.360 ;
    END
  END core_wb_data_o[1]
  PIN core_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 367.920 500.000 368.520 ;
    END
  END core_wb_data_o[20]
  PIN core_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 382.880 500.000 383.480 ;
    END
  END core_wb_data_o[21]
  PIN core_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 397.840 500.000 398.440 ;
    END
  END core_wb_data_o[22]
  PIN core_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 412.800 500.000 413.400 ;
    END
  END core_wb_data_o[23]
  PIN core_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 427.760 500.000 428.360 ;
    END
  END core_wb_data_o[24]
  PIN core_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 442.720 500.000 443.320 ;
    END
  END core_wb_data_o[25]
  PIN core_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 457.000 500.000 457.600 ;
    END
  END core_wb_data_o[26]
  PIN core_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 471.960 500.000 472.560 ;
    END
  END core_wb_data_o[27]
  PIN core_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 482.160 500.000 482.760 ;
    END
  END core_wb_data_o[28]
  PIN core_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 491.680 500.000 492.280 ;
    END
  END core_wb_data_o[29]
  PIN core_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 91.160 500.000 91.760 ;
    END
  END core_wb_data_o[2]
  PIN core_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 501.880 500.000 502.480 ;
    END
  END core_wb_data_o[30]
  PIN core_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 512.080 500.000 512.680 ;
    END
  END core_wb_data_o[31]
  PIN core_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 110.880 500.000 111.480 ;
    END
  END core_wb_data_o[3]
  PIN core_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 130.600 500.000 131.200 ;
    END
  END core_wb_data_o[4]
  PIN core_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 145.560 500.000 146.160 ;
    END
  END core_wb_data_o[5]
  PIN core_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 160.520 500.000 161.120 ;
    END
  END core_wb_data_o[6]
  PIN core_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 174.800 500.000 175.400 ;
    END
  END core_wb_data_o[7]
  PIN core_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 189.760 500.000 190.360 ;
    END
  END core_wb_data_o[8]
  PIN core_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 204.720 500.000 205.320 ;
    END
  END core_wb_data_o[9]
  PIN core_wb_error_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 21.800 500.000 22.400 ;
    END
  END core_wb_error_i
  PIN core_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 56.480 500.000 57.080 ;
    END
  END core_wb_sel_o[0]
  PIN core_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 76.200 500.000 76.800 ;
    END
  END core_wb_sel_o[1]
  PIN core_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.920 500.000 96.520 ;
    END
  END core_wb_sel_o[2]
  PIN core_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 115.640 500.000 116.240 ;
    END
  END core_wb_sel_o[3]
  PIN core_wb_stall_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 26.560 500.000 27.160 ;
    END
  END core_wb_stall_i
  PIN core_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 31.320 500.000 31.920 ;
    END
  END core_wb_stb_o
  PIN core_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 36.080 500.000 36.680 ;
    END
  END core_wb_we_o
  PIN csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END csb0[0]
  PIN csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END csb0[1]
  PIN csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END csb1[0]
  PIN csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.160 4.000 618.760 ;
    END
  END csb1[1]
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END din0[9]
  PIN dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.560 4.000 401.160 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.400 4.000 427.000 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END dout0[32]
  PIN dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END dout0[33]
  PIN dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END dout0[34]
  PIN dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END dout0[35]
  PIN dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END dout0[36]
  PIN dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END dout0[37]
  PIN dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END dout0[38]
  PIN dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END dout0[39]
  PIN dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END dout0[3]
  PIN dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 483.520 4.000 484.120 ;
    END
  END dout0[40]
  PIN dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END dout0[41]
  PIN dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 494.400 4.000 495.000 ;
    END
  END dout0[42]
  PIN dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END dout0[43]
  PIN dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END dout0[44]
  PIN dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 509.360 4.000 509.960 ;
    END
  END dout0[45]
  PIN dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END dout0[46]
  PIN dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END dout0[47]
  PIN dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END dout0[48]
  PIN dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END dout0[49]
  PIN dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END dout0[4]
  PIN dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END dout0[50]
  PIN dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END dout0[51]
  PIN dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.080 4.000 546.680 ;
    END
  END dout0[52]
  PIN dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END dout0[53]
  PIN dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END dout0[54]
  PIN dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END dout0[55]
  PIN dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 4.000 567.080 ;
    END
  END dout0[56]
  PIN dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END dout0[57]
  PIN dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 577.360 4.000 577.960 ;
    END
  END dout0[58]
  PIN dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END dout0[59]
  PIN dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END dout0[5]
  PIN dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END dout0[60]
  PIN dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END dout0[61]
  PIN dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.760 4.000 598.360 ;
    END
  END dout0[62]
  PIN dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END dout0[63]
  PIN dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END dout0[9]
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 732.400 4.000 733.000 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 742.600 4.000 743.200 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 753.480 4.000 754.080 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.680 4.000 764.280 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.120 4.000 769.720 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.280 4.000 675.880 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.880 4.000 774.480 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.080 4.000 784.680 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 789.520 4.000 790.120 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.960 4.000 795.560 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.160 4.000 805.760 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.920 4.000 810.520 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.800 4.000 821.400 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.000 4.000 831.600 ;
    END
  END dout1[31]
  PIN dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END dout1[32]
  PIN dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 841.200 4.000 841.800 ;
    END
  END dout1[33]
  PIN dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END dout1[34]
  PIN dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 851.400 4.000 852.000 ;
    END
  END dout1[35]
  PIN dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END dout1[36]
  PIN dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END dout1[37]
  PIN dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END dout1[38]
  PIN dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 872.480 4.000 873.080 ;
    END
  END dout1[39]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.160 4.000 686.760 ;
    END
  END dout1[3]
  PIN dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.920 4.000 878.520 ;
    END
  END dout1[40]
  PIN dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 882.680 4.000 883.280 ;
    END
  END dout1[41]
  PIN dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END dout1[42]
  PIN dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.880 4.000 893.480 ;
    END
  END dout1[43]
  PIN dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 898.320 4.000 898.920 ;
    END
  END dout1[44]
  PIN dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.760 4.000 904.360 ;
    END
  END dout1[45]
  PIN dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 908.520 4.000 909.120 ;
    END
  END dout1[46]
  PIN dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 913.960 4.000 914.560 ;
    END
  END dout1[47]
  PIN dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 919.400 4.000 920.000 ;
    END
  END dout1[48]
  PIN dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.160 4.000 924.760 ;
    END
  END dout1[49]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END dout1[4]
  PIN dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 929.600 4.000 930.200 ;
    END
  END dout1[50]
  PIN dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 934.360 4.000 934.960 ;
    END
  END dout1[51]
  PIN dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.800 4.000 940.400 ;
    END
  END dout1[52]
  PIN dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END dout1[53]
  PIN dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.000 4.000 950.600 ;
    END
  END dout1[54]
  PIN dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END dout1[55]
  PIN dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.880 4.000 961.480 ;
    END
  END dout1[56]
  PIN dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END dout1[57]
  PIN dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END dout1[58]
  PIN dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END dout1[59]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END dout1[5]
  PIN dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.280 4.000 981.880 ;
    END
  END dout1[60]
  PIN dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.720 4.000 987.320 ;
    END
  END dout1[61]
  PIN dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 991.480 4.000 992.080 ;
    END
  END dout1[62]
  PIN dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.920 4.000 997.520 ;
    END
  END dout1[63]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.120 4.000 701.720 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 706.560 4.000 707.160 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.000 4.000 712.600 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END dout1[9]
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END irq[0]
  PIN irq[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END irq[10]
  PIN irq[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END irq[11]
  PIN irq[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END irq[12]
  PIN irq[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END irq[13]
  PIN irq[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END irq[14]
  PIN irq[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END irq[15]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END irq[2]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END irq[5]
  PIN irq[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END irq[6]
  PIN irq[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END irq[7]
  PIN irq[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END irq[8]
  PIN irq[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END irq[9]
  PIN jtag_tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END jtag_tms
  PIN localMemory_wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 516.840 500.000 517.440 ;
    END
  END localMemory_wb_ack_o
  PIN localMemory_wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 546.760 500.000 547.360 ;
    END
  END localMemory_wb_adr_i[0]
  PIN localMemory_wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 714.720 500.000 715.320 ;
    END
  END localMemory_wb_adr_i[10]
  PIN localMemory_wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 729.680 500.000 730.280 ;
    END
  END localMemory_wb_adr_i[11]
  PIN localMemory_wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 744.640 500.000 745.240 ;
    END
  END localMemory_wb_adr_i[12]
  PIN localMemory_wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 759.600 500.000 760.200 ;
    END
  END localMemory_wb_adr_i[13]
  PIN localMemory_wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 774.560 500.000 775.160 ;
    END
  END localMemory_wb_adr_i[14]
  PIN localMemory_wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 788.840 500.000 789.440 ;
    END
  END localMemory_wb_adr_i[15]
  PIN localMemory_wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 803.800 500.000 804.400 ;
    END
  END localMemory_wb_adr_i[16]
  PIN localMemory_wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 818.760 500.000 819.360 ;
    END
  END localMemory_wb_adr_i[17]
  PIN localMemory_wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 833.720 500.000 834.320 ;
    END
  END localMemory_wb_adr_i[18]
  PIN localMemory_wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 848.680 500.000 849.280 ;
    END
  END localMemory_wb_adr_i[19]
  PIN localMemory_wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 566.480 500.000 567.080 ;
    END
  END localMemory_wb_adr_i[1]
  PIN localMemory_wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 863.640 500.000 864.240 ;
    END
  END localMemory_wb_adr_i[20]
  PIN localMemory_wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 877.920 500.000 878.520 ;
    END
  END localMemory_wb_adr_i[21]
  PIN localMemory_wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 892.880 500.000 893.480 ;
    END
  END localMemory_wb_adr_i[22]
  PIN localMemory_wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 907.840 500.000 908.440 ;
    END
  END localMemory_wb_adr_i[23]
  PIN localMemory_wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 586.200 500.000 586.800 ;
    END
  END localMemory_wb_adr_i[2]
  PIN localMemory_wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 605.920 500.000 606.520 ;
    END
  END localMemory_wb_adr_i[3]
  PIN localMemory_wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 625.640 500.000 626.240 ;
    END
  END localMemory_wb_adr_i[4]
  PIN localMemory_wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 640.600 500.000 641.200 ;
    END
  END localMemory_wb_adr_i[5]
  PIN localMemory_wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 655.560 500.000 656.160 ;
    END
  END localMemory_wb_adr_i[6]
  PIN localMemory_wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 670.520 500.000 671.120 ;
    END
  END localMemory_wb_adr_i[7]
  PIN localMemory_wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 684.800 500.000 685.400 ;
    END
  END localMemory_wb_adr_i[8]
  PIN localMemory_wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 699.760 500.000 700.360 ;
    END
  END localMemory_wb_adr_i[9]
  PIN localMemory_wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 521.600 500.000 522.200 ;
    END
  END localMemory_wb_cyc_i
  PIN localMemory_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 551.520 500.000 552.120 ;
    END
  END localMemory_wb_data_i[0]
  PIN localMemory_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 719.480 500.000 720.080 ;
    END
  END localMemory_wb_data_i[10]
  PIN localMemory_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 734.440 500.000 735.040 ;
    END
  END localMemory_wb_data_i[11]
  PIN localMemory_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 749.400 500.000 750.000 ;
    END
  END localMemory_wb_data_i[12]
  PIN localMemory_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 764.360 500.000 764.960 ;
    END
  END localMemory_wb_data_i[13]
  PIN localMemory_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 779.320 500.000 779.920 ;
    END
  END localMemory_wb_data_i[14]
  PIN localMemory_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 794.280 500.000 794.880 ;
    END
  END localMemory_wb_data_i[15]
  PIN localMemory_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 808.560 500.000 809.160 ;
    END
  END localMemory_wb_data_i[16]
  PIN localMemory_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 823.520 500.000 824.120 ;
    END
  END localMemory_wb_data_i[17]
  PIN localMemory_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 838.480 500.000 839.080 ;
    END
  END localMemory_wb_data_i[18]
  PIN localMemory_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 853.440 500.000 854.040 ;
    END
  END localMemory_wb_data_i[19]
  PIN localMemory_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 571.240 500.000 571.840 ;
    END
  END localMemory_wb_data_i[1]
  PIN localMemory_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 868.400 500.000 869.000 ;
    END
  END localMemory_wb_data_i[20]
  PIN localMemory_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 883.360 500.000 883.960 ;
    END
  END localMemory_wb_data_i[21]
  PIN localMemory_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 898.320 500.000 898.920 ;
    END
  END localMemory_wb_data_i[22]
  PIN localMemory_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 912.600 500.000 913.200 ;
    END
  END localMemory_wb_data_i[23]
  PIN localMemory_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 922.800 500.000 923.400 ;
    END
  END localMemory_wb_data_i[24]
  PIN localMemory_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 933.000 500.000 933.600 ;
    END
  END localMemory_wb_data_i[25]
  PIN localMemory_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 942.520 500.000 943.120 ;
    END
  END localMemory_wb_data_i[26]
  PIN localMemory_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 952.720 500.000 953.320 ;
    END
  END localMemory_wb_data_i[27]
  PIN localMemory_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 962.240 500.000 962.840 ;
    END
  END localMemory_wb_data_i[28]
  PIN localMemory_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 972.440 500.000 973.040 ;
    END
  END localMemory_wb_data_i[29]
  PIN localMemory_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 590.960 500.000 591.560 ;
    END
  END localMemory_wb_data_i[2]
  PIN localMemory_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 981.960 500.000 982.560 ;
    END
  END localMemory_wb_data_i[30]
  PIN localMemory_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 992.160 500.000 992.760 ;
    END
  END localMemory_wb_data_i[31]
  PIN localMemory_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 610.680 500.000 611.280 ;
    END
  END localMemory_wb_data_i[3]
  PIN localMemory_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 630.400 500.000 631.000 ;
    END
  END localMemory_wb_data_i[4]
  PIN localMemory_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 645.360 500.000 645.960 ;
    END
  END localMemory_wb_data_i[5]
  PIN localMemory_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 660.320 500.000 660.920 ;
    END
  END localMemory_wb_data_i[6]
  PIN localMemory_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 675.280 500.000 675.880 ;
    END
  END localMemory_wb_data_i[7]
  PIN localMemory_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 690.240 500.000 690.840 ;
    END
  END localMemory_wb_data_i[8]
  PIN localMemory_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 705.200 500.000 705.800 ;
    END
  END localMemory_wb_data_i[9]
  PIN localMemory_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 556.280 500.000 556.880 ;
    END
  END localMemory_wb_data_o[0]
  PIN localMemory_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 724.920 500.000 725.520 ;
    END
  END localMemory_wb_data_o[10]
  PIN localMemory_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 739.880 500.000 740.480 ;
    END
  END localMemory_wb_data_o[11]
  PIN localMemory_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 754.160 500.000 754.760 ;
    END
  END localMemory_wb_data_o[12]
  PIN localMemory_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 769.120 500.000 769.720 ;
    END
  END localMemory_wb_data_o[13]
  PIN localMemory_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 784.080 500.000 784.680 ;
    END
  END localMemory_wb_data_o[14]
  PIN localMemory_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 799.040 500.000 799.640 ;
    END
  END localMemory_wb_data_o[15]
  PIN localMemory_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 814.000 500.000 814.600 ;
    END
  END localMemory_wb_data_o[16]
  PIN localMemory_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 828.960 500.000 829.560 ;
    END
  END localMemory_wb_data_o[17]
  PIN localMemory_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 843.240 500.000 843.840 ;
    END
  END localMemory_wb_data_o[18]
  PIN localMemory_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 858.200 500.000 858.800 ;
    END
  END localMemory_wb_data_o[19]
  PIN localMemory_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 576.000 500.000 576.600 ;
    END
  END localMemory_wb_data_o[1]
  PIN localMemory_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 873.160 500.000 873.760 ;
    END
  END localMemory_wb_data_o[20]
  PIN localMemory_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 888.120 500.000 888.720 ;
    END
  END localMemory_wb_data_o[21]
  PIN localMemory_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 903.080 500.000 903.680 ;
    END
  END localMemory_wb_data_o[22]
  PIN localMemory_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 918.040 500.000 918.640 ;
    END
  END localMemory_wb_data_o[23]
  PIN localMemory_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 927.560 500.000 928.160 ;
    END
  END localMemory_wb_data_o[24]
  PIN localMemory_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 937.760 500.000 938.360 ;
    END
  END localMemory_wb_data_o[25]
  PIN localMemory_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 947.280 500.000 947.880 ;
    END
  END localMemory_wb_data_o[26]
  PIN localMemory_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 957.480 500.000 958.080 ;
    END
  END localMemory_wb_data_o[27]
  PIN localMemory_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 967.680 500.000 968.280 ;
    END
  END localMemory_wb_data_o[28]
  PIN localMemory_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 977.200 500.000 977.800 ;
    END
  END localMemory_wb_data_o[29]
  PIN localMemory_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 595.720 500.000 596.320 ;
    END
  END localMemory_wb_data_o[2]
  PIN localMemory_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 987.400 500.000 988.000 ;
    END
  END localMemory_wb_data_o[30]
  PIN localMemory_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 996.920 500.000 997.520 ;
    END
  END localMemory_wb_data_o[31]
  PIN localMemory_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 615.440 500.000 616.040 ;
    END
  END localMemory_wb_data_o[3]
  PIN localMemory_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 635.840 500.000 636.440 ;
    END
  END localMemory_wb_data_o[4]
  PIN localMemory_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 650.120 500.000 650.720 ;
    END
  END localMemory_wb_data_o[5]
  PIN localMemory_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 665.080 500.000 665.680 ;
    END
  END localMemory_wb_data_o[6]
  PIN localMemory_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 680.040 500.000 680.640 ;
    END
  END localMemory_wb_data_o[7]
  PIN localMemory_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 695.000 500.000 695.600 ;
    END
  END localMemory_wb_data_o[8]
  PIN localMemory_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 709.960 500.000 710.560 ;
    END
  END localMemory_wb_data_o[9]
  PIN localMemory_wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 526.360 500.000 526.960 ;
    END
  END localMemory_wb_error_o
  PIN localMemory_wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 561.040 500.000 561.640 ;
    END
  END localMemory_wb_sel_i[0]
  PIN localMemory_wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 581.440 500.000 582.040 ;
    END
  END localMemory_wb_sel_i[1]
  PIN localMemory_wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 601.160 500.000 601.760 ;
    END
  END localMemory_wb_sel_i[2]
  PIN localMemory_wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 620.880 500.000 621.480 ;
    END
  END localMemory_wb_sel_i[3]
  PIN localMemory_wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 531.800 500.000 532.400 ;
    END
  END localMemory_wb_stall_o
  PIN localMemory_wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 536.560 500.000 537.160 ;
    END
  END localMemory_wb_stb_i
  PIN localMemory_wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 541.320 500.000 541.920 ;
    END
  END localMemory_wb_we_i
  PIN manufacturerID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 996.000 108.470 1000.000 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 996.000 236.810 1000.000 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 996.000 121.350 1000.000 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 996.000 134.230 1000.000 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 996.000 147.110 1000.000 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 996.000 159.990 1000.000 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 996.000 172.870 1000.000 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 996.000 185.750 1000.000 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 996.000 198.630 1000.000 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 996.000 211.050 1000.000 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 996.000 223.930 1000.000 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 996.000 249.690 1000.000 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 996.000 378.030 1000.000 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 996.000 390.910 1000.000 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 996.000 403.790 1000.000 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 996.000 416.210 1000.000 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 996.000 429.090 1000.000 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 996.000 441.970 1000.000 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 996.000 262.570 1000.000 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 996.000 275.450 1000.000 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 996.000 288.330 1000.000 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 996.000 301.210 1000.000 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 996.000 313.630 1000.000 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 996.000 326.510 1000.000 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 996.000 339.390 1000.000 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 996.000 352.270 1000.000 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 996.000 365.150 1000.000 ;
    END
  END partID[9]
  PIN probe_env[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END probe_env[0]
  PIN probe_env[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END probe_env[1]
  PIN probe_errorCode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END probe_errorCode[0]
  PIN probe_errorCode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END probe_errorCode[1]
  PIN probe_isBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END probe_isBranch
  PIN probe_isCompressed
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END probe_isCompressed
  PIN probe_isLoad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END probe_isLoad
  PIN probe_isStore
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END probe_isStore
  PIN probe_jtagInstruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END probe_jtagInstruction[0]
  PIN probe_jtagInstruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END probe_jtagInstruction[1]
  PIN probe_jtagInstruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END probe_jtagInstruction[2]
  PIN probe_jtagInstruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END probe_jtagInstruction[3]
  PIN probe_jtagInstruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END probe_jtagInstruction[4]
  PIN probe_opcode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END probe_opcode[0]
  PIN probe_opcode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END probe_opcode[1]
  PIN probe_opcode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END probe_opcode[2]
  PIN probe_opcode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END probe_opcode[3]
  PIN probe_opcode[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END probe_opcode[4]
  PIN probe_opcode[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END probe_opcode[5]
  PIN probe_opcode[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END probe_opcode[6]
  PIN probe_programCounter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END probe_programCounter[0]
  PIN probe_programCounter[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END probe_programCounter[10]
  PIN probe_programCounter[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END probe_programCounter[11]
  PIN probe_programCounter[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END probe_programCounter[12]
  PIN probe_programCounter[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END probe_programCounter[13]
  PIN probe_programCounter[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END probe_programCounter[14]
  PIN probe_programCounter[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END probe_programCounter[15]
  PIN probe_programCounter[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END probe_programCounter[16]
  PIN probe_programCounter[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END probe_programCounter[17]
  PIN probe_programCounter[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END probe_programCounter[18]
  PIN probe_programCounter[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END probe_programCounter[19]
  PIN probe_programCounter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END probe_programCounter[1]
  PIN probe_programCounter[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END probe_programCounter[20]
  PIN probe_programCounter[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END probe_programCounter[21]
  PIN probe_programCounter[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END probe_programCounter[22]
  PIN probe_programCounter[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END probe_programCounter[23]
  PIN probe_programCounter[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END probe_programCounter[24]
  PIN probe_programCounter[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END probe_programCounter[25]
  PIN probe_programCounter[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END probe_programCounter[26]
  PIN probe_programCounter[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END probe_programCounter[27]
  PIN probe_programCounter[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END probe_programCounter[28]
  PIN probe_programCounter[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END probe_programCounter[29]
  PIN probe_programCounter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END probe_programCounter[2]
  PIN probe_programCounter[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END probe_programCounter[30]
  PIN probe_programCounter[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END probe_programCounter[31]
  PIN probe_programCounter[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END probe_programCounter[3]
  PIN probe_programCounter[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END probe_programCounter[4]
  PIN probe_programCounter[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END probe_programCounter[5]
  PIN probe_programCounter[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END probe_programCounter[6]
  PIN probe_programCounter[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END probe_programCounter[7]
  PIN probe_programCounter[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END probe_programCounter[8]
  PIN probe_programCounter[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END probe_programCounter[9]
  PIN probe_state[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END probe_state[0]
  PIN probe_state[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END probe_state[1]
  PIN probe_takeBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END probe_takeBranch
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 987.600 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 996.000 454.850 1000.000 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 996.000 467.730 1000.000 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 996.000 480.610 1000.000 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 996.000 493.490 1000.000 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 987.600 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 2.080 500.000 2.680 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 6.840 500.000 7.440 ;
    END
  END wb_rst_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 987.445 ;
      LAYER met1 ;
        RECT 2.830 6.500 499.950 987.600 ;
      LAYER met2 ;
        RECT 2.860 995.720 5.790 997.405 ;
        RECT 6.630 995.720 18.210 997.405 ;
        RECT 19.050 995.720 31.090 997.405 ;
        RECT 31.930 995.720 43.970 997.405 ;
        RECT 44.810 995.720 56.850 997.405 ;
        RECT 57.690 995.720 69.730 997.405 ;
        RECT 70.570 995.720 82.610 997.405 ;
        RECT 83.450 995.720 95.490 997.405 ;
        RECT 96.330 995.720 107.910 997.405 ;
        RECT 108.750 995.720 120.790 997.405 ;
        RECT 121.630 995.720 133.670 997.405 ;
        RECT 134.510 995.720 146.550 997.405 ;
        RECT 147.390 995.720 159.430 997.405 ;
        RECT 160.270 995.720 172.310 997.405 ;
        RECT 173.150 995.720 185.190 997.405 ;
        RECT 186.030 995.720 198.070 997.405 ;
        RECT 198.910 995.720 210.490 997.405 ;
        RECT 211.330 995.720 223.370 997.405 ;
        RECT 224.210 995.720 236.250 997.405 ;
        RECT 237.090 995.720 249.130 997.405 ;
        RECT 249.970 995.720 262.010 997.405 ;
        RECT 262.850 995.720 274.890 997.405 ;
        RECT 275.730 995.720 287.770 997.405 ;
        RECT 288.610 995.720 300.650 997.405 ;
        RECT 301.490 995.720 313.070 997.405 ;
        RECT 313.910 995.720 325.950 997.405 ;
        RECT 326.790 995.720 338.830 997.405 ;
        RECT 339.670 995.720 351.710 997.405 ;
        RECT 352.550 995.720 364.590 997.405 ;
        RECT 365.430 995.720 377.470 997.405 ;
        RECT 378.310 995.720 390.350 997.405 ;
        RECT 391.190 995.720 403.230 997.405 ;
        RECT 404.070 995.720 415.650 997.405 ;
        RECT 416.490 995.720 428.530 997.405 ;
        RECT 429.370 995.720 441.410 997.405 ;
        RECT 442.250 995.720 454.290 997.405 ;
        RECT 455.130 995.720 467.170 997.405 ;
        RECT 468.010 995.720 480.050 997.405 ;
        RECT 480.890 995.720 492.930 997.405 ;
        RECT 493.770 995.720 499.930 997.405 ;
        RECT 2.860 4.280 499.930 995.720 ;
        RECT 2.860 2.195 3.030 4.280 ;
        RECT 3.870 2.195 9.930 4.280 ;
        RECT 10.770 2.195 16.830 4.280 ;
        RECT 17.670 2.195 23.730 4.280 ;
        RECT 24.570 2.195 31.090 4.280 ;
        RECT 31.930 2.195 37.990 4.280 ;
        RECT 38.830 2.195 44.890 4.280 ;
        RECT 45.730 2.195 52.250 4.280 ;
        RECT 53.090 2.195 59.150 4.280 ;
        RECT 59.990 2.195 66.050 4.280 ;
        RECT 66.890 2.195 73.410 4.280 ;
        RECT 74.250 2.195 80.310 4.280 ;
        RECT 81.150 2.195 87.210 4.280 ;
        RECT 88.050 2.195 94.570 4.280 ;
        RECT 95.410 2.195 101.470 4.280 ;
        RECT 102.310 2.195 108.370 4.280 ;
        RECT 109.210 2.195 115.270 4.280 ;
        RECT 116.110 2.195 122.630 4.280 ;
        RECT 123.470 2.195 129.530 4.280 ;
        RECT 130.370 2.195 136.430 4.280 ;
        RECT 137.270 2.195 143.790 4.280 ;
        RECT 144.630 2.195 150.690 4.280 ;
        RECT 151.530 2.195 157.590 4.280 ;
        RECT 158.430 2.195 164.950 4.280 ;
        RECT 165.790 2.195 171.850 4.280 ;
        RECT 172.690 2.195 178.750 4.280 ;
        RECT 179.590 2.195 186.110 4.280 ;
        RECT 186.950 2.195 193.010 4.280 ;
        RECT 193.850 2.195 199.910 4.280 ;
        RECT 200.750 2.195 206.810 4.280 ;
        RECT 207.650 2.195 214.170 4.280 ;
        RECT 215.010 2.195 221.070 4.280 ;
        RECT 221.910 2.195 227.970 4.280 ;
        RECT 228.810 2.195 235.330 4.280 ;
        RECT 236.170 2.195 242.230 4.280 ;
        RECT 243.070 2.195 249.130 4.280 ;
        RECT 249.970 2.195 256.490 4.280 ;
        RECT 257.330 2.195 263.390 4.280 ;
        RECT 264.230 2.195 270.290 4.280 ;
        RECT 271.130 2.195 277.650 4.280 ;
        RECT 278.490 2.195 284.550 4.280 ;
        RECT 285.390 2.195 291.450 4.280 ;
        RECT 292.290 2.195 298.810 4.280 ;
        RECT 299.650 2.195 305.710 4.280 ;
        RECT 306.550 2.195 312.610 4.280 ;
        RECT 313.450 2.195 319.510 4.280 ;
        RECT 320.350 2.195 326.870 4.280 ;
        RECT 327.710 2.195 333.770 4.280 ;
        RECT 334.610 2.195 340.670 4.280 ;
        RECT 341.510 2.195 348.030 4.280 ;
        RECT 348.870 2.195 354.930 4.280 ;
        RECT 355.770 2.195 361.830 4.280 ;
        RECT 362.670 2.195 369.190 4.280 ;
        RECT 370.030 2.195 376.090 4.280 ;
        RECT 376.930 2.195 382.990 4.280 ;
        RECT 383.830 2.195 390.350 4.280 ;
        RECT 391.190 2.195 397.250 4.280 ;
        RECT 398.090 2.195 404.150 4.280 ;
        RECT 404.990 2.195 411.050 4.280 ;
        RECT 411.890 2.195 418.410 4.280 ;
        RECT 419.250 2.195 425.310 4.280 ;
        RECT 426.150 2.195 432.210 4.280 ;
        RECT 433.050 2.195 439.570 4.280 ;
        RECT 440.410 2.195 446.470 4.280 ;
        RECT 447.310 2.195 453.370 4.280 ;
        RECT 454.210 2.195 460.730 4.280 ;
        RECT 461.570 2.195 467.630 4.280 ;
        RECT 468.470 2.195 474.530 4.280 ;
        RECT 475.370 2.195 481.890 4.280 ;
        RECT 482.730 2.195 488.790 4.280 ;
        RECT 489.630 2.195 495.690 4.280 ;
        RECT 496.530 2.195 499.930 4.280 ;
      LAYER met3 ;
        RECT 4.400 996.520 495.600 997.385 ;
        RECT 3.285 993.160 499.955 996.520 ;
        RECT 3.285 992.480 495.600 993.160 ;
        RECT 4.400 991.760 495.600 992.480 ;
        RECT 4.400 991.080 499.955 991.760 ;
        RECT 3.285 988.400 499.955 991.080 ;
        RECT 3.285 987.720 495.600 988.400 ;
        RECT 4.400 987.000 495.600 987.720 ;
        RECT 4.400 986.320 499.955 987.000 ;
        RECT 3.285 982.960 499.955 986.320 ;
        RECT 3.285 982.280 495.600 982.960 ;
        RECT 4.400 981.560 495.600 982.280 ;
        RECT 4.400 980.880 499.955 981.560 ;
        RECT 3.285 978.200 499.955 980.880 ;
        RECT 3.285 976.840 495.600 978.200 ;
        RECT 4.400 976.800 495.600 976.840 ;
        RECT 4.400 975.440 499.955 976.800 ;
        RECT 3.285 973.440 499.955 975.440 ;
        RECT 3.285 972.080 495.600 973.440 ;
        RECT 4.400 972.040 495.600 972.080 ;
        RECT 4.400 970.680 499.955 972.040 ;
        RECT 3.285 968.680 499.955 970.680 ;
        RECT 3.285 967.280 495.600 968.680 ;
        RECT 3.285 966.640 499.955 967.280 ;
        RECT 4.400 965.240 499.955 966.640 ;
        RECT 3.285 963.240 499.955 965.240 ;
        RECT 3.285 961.880 495.600 963.240 ;
        RECT 4.400 961.840 495.600 961.880 ;
        RECT 4.400 960.480 499.955 961.840 ;
        RECT 3.285 958.480 499.955 960.480 ;
        RECT 3.285 957.080 495.600 958.480 ;
        RECT 3.285 956.440 499.955 957.080 ;
        RECT 4.400 955.040 499.955 956.440 ;
        RECT 3.285 953.720 499.955 955.040 ;
        RECT 3.285 952.320 495.600 953.720 ;
        RECT 3.285 951.000 499.955 952.320 ;
        RECT 4.400 949.600 499.955 951.000 ;
        RECT 3.285 948.280 499.955 949.600 ;
        RECT 3.285 946.880 495.600 948.280 ;
        RECT 3.285 946.240 499.955 946.880 ;
        RECT 4.400 944.840 499.955 946.240 ;
        RECT 3.285 943.520 499.955 944.840 ;
        RECT 3.285 942.120 495.600 943.520 ;
        RECT 3.285 940.800 499.955 942.120 ;
        RECT 4.400 939.400 499.955 940.800 ;
        RECT 3.285 938.760 499.955 939.400 ;
        RECT 3.285 937.360 495.600 938.760 ;
        RECT 3.285 935.360 499.955 937.360 ;
        RECT 4.400 934.000 499.955 935.360 ;
        RECT 4.400 933.960 495.600 934.000 ;
        RECT 3.285 932.600 495.600 933.960 ;
        RECT 3.285 930.600 499.955 932.600 ;
        RECT 4.400 929.200 499.955 930.600 ;
        RECT 3.285 928.560 499.955 929.200 ;
        RECT 3.285 927.160 495.600 928.560 ;
        RECT 3.285 925.160 499.955 927.160 ;
        RECT 4.400 923.800 499.955 925.160 ;
        RECT 4.400 923.760 495.600 923.800 ;
        RECT 3.285 922.400 495.600 923.760 ;
        RECT 3.285 920.400 499.955 922.400 ;
        RECT 4.400 919.040 499.955 920.400 ;
        RECT 4.400 919.000 495.600 919.040 ;
        RECT 3.285 917.640 495.600 919.000 ;
        RECT 3.285 914.960 499.955 917.640 ;
        RECT 4.400 913.600 499.955 914.960 ;
        RECT 4.400 913.560 495.600 913.600 ;
        RECT 3.285 912.200 495.600 913.560 ;
        RECT 3.285 909.520 499.955 912.200 ;
        RECT 4.400 908.840 499.955 909.520 ;
        RECT 4.400 908.120 495.600 908.840 ;
        RECT 3.285 907.440 495.600 908.120 ;
        RECT 3.285 904.760 499.955 907.440 ;
        RECT 4.400 904.080 499.955 904.760 ;
        RECT 4.400 903.360 495.600 904.080 ;
        RECT 3.285 902.680 495.600 903.360 ;
        RECT 3.285 899.320 499.955 902.680 ;
        RECT 4.400 897.920 495.600 899.320 ;
        RECT 3.285 893.880 499.955 897.920 ;
        RECT 4.400 892.480 495.600 893.880 ;
        RECT 3.285 889.120 499.955 892.480 ;
        RECT 4.400 887.720 495.600 889.120 ;
        RECT 3.285 884.360 499.955 887.720 ;
        RECT 3.285 883.680 495.600 884.360 ;
        RECT 4.400 882.960 495.600 883.680 ;
        RECT 4.400 882.280 499.955 882.960 ;
        RECT 3.285 878.920 499.955 882.280 ;
        RECT 4.400 877.520 495.600 878.920 ;
        RECT 3.285 874.160 499.955 877.520 ;
        RECT 3.285 873.480 495.600 874.160 ;
        RECT 4.400 872.760 495.600 873.480 ;
        RECT 4.400 872.080 499.955 872.760 ;
        RECT 3.285 869.400 499.955 872.080 ;
        RECT 3.285 868.040 495.600 869.400 ;
        RECT 4.400 868.000 495.600 868.040 ;
        RECT 4.400 866.640 499.955 868.000 ;
        RECT 3.285 864.640 499.955 866.640 ;
        RECT 3.285 863.280 495.600 864.640 ;
        RECT 4.400 863.240 495.600 863.280 ;
        RECT 4.400 861.880 499.955 863.240 ;
        RECT 3.285 859.200 499.955 861.880 ;
        RECT 3.285 857.840 495.600 859.200 ;
        RECT 4.400 857.800 495.600 857.840 ;
        RECT 4.400 856.440 499.955 857.800 ;
        RECT 3.285 854.440 499.955 856.440 ;
        RECT 3.285 853.040 495.600 854.440 ;
        RECT 3.285 852.400 499.955 853.040 ;
        RECT 4.400 851.000 499.955 852.400 ;
        RECT 3.285 849.680 499.955 851.000 ;
        RECT 3.285 848.280 495.600 849.680 ;
        RECT 3.285 847.640 499.955 848.280 ;
        RECT 4.400 846.240 499.955 847.640 ;
        RECT 3.285 844.240 499.955 846.240 ;
        RECT 3.285 842.840 495.600 844.240 ;
        RECT 3.285 842.200 499.955 842.840 ;
        RECT 4.400 840.800 499.955 842.200 ;
        RECT 3.285 839.480 499.955 840.800 ;
        RECT 3.285 838.080 495.600 839.480 ;
        RECT 3.285 837.440 499.955 838.080 ;
        RECT 4.400 836.040 499.955 837.440 ;
        RECT 3.285 834.720 499.955 836.040 ;
        RECT 3.285 833.320 495.600 834.720 ;
        RECT 3.285 832.000 499.955 833.320 ;
        RECT 4.400 830.600 499.955 832.000 ;
        RECT 3.285 829.960 499.955 830.600 ;
        RECT 3.285 828.560 495.600 829.960 ;
        RECT 3.285 826.560 499.955 828.560 ;
        RECT 4.400 825.160 499.955 826.560 ;
        RECT 3.285 824.520 499.955 825.160 ;
        RECT 3.285 823.120 495.600 824.520 ;
        RECT 3.285 821.800 499.955 823.120 ;
        RECT 4.400 820.400 499.955 821.800 ;
        RECT 3.285 819.760 499.955 820.400 ;
        RECT 3.285 818.360 495.600 819.760 ;
        RECT 3.285 816.360 499.955 818.360 ;
        RECT 4.400 815.000 499.955 816.360 ;
        RECT 4.400 814.960 495.600 815.000 ;
        RECT 3.285 813.600 495.600 814.960 ;
        RECT 3.285 810.920 499.955 813.600 ;
        RECT 4.400 809.560 499.955 810.920 ;
        RECT 4.400 809.520 495.600 809.560 ;
        RECT 3.285 808.160 495.600 809.520 ;
        RECT 3.285 806.160 499.955 808.160 ;
        RECT 4.400 804.800 499.955 806.160 ;
        RECT 4.400 804.760 495.600 804.800 ;
        RECT 3.285 803.400 495.600 804.760 ;
        RECT 3.285 800.720 499.955 803.400 ;
        RECT 4.400 800.040 499.955 800.720 ;
        RECT 4.400 799.320 495.600 800.040 ;
        RECT 3.285 798.640 495.600 799.320 ;
        RECT 3.285 795.960 499.955 798.640 ;
        RECT 4.400 795.280 499.955 795.960 ;
        RECT 4.400 794.560 495.600 795.280 ;
        RECT 3.285 793.880 495.600 794.560 ;
        RECT 3.285 790.520 499.955 793.880 ;
        RECT 4.400 789.840 499.955 790.520 ;
        RECT 4.400 789.120 495.600 789.840 ;
        RECT 3.285 788.440 495.600 789.120 ;
        RECT 3.285 785.080 499.955 788.440 ;
        RECT 4.400 783.680 495.600 785.080 ;
        RECT 3.285 780.320 499.955 783.680 ;
        RECT 4.400 778.920 495.600 780.320 ;
        RECT 3.285 775.560 499.955 778.920 ;
        RECT 3.285 774.880 495.600 775.560 ;
        RECT 4.400 774.160 495.600 774.880 ;
        RECT 4.400 773.480 499.955 774.160 ;
        RECT 3.285 770.120 499.955 773.480 ;
        RECT 4.400 768.720 495.600 770.120 ;
        RECT 3.285 765.360 499.955 768.720 ;
        RECT 3.285 764.680 495.600 765.360 ;
        RECT 4.400 763.960 495.600 764.680 ;
        RECT 4.400 763.280 499.955 763.960 ;
        RECT 3.285 760.600 499.955 763.280 ;
        RECT 3.285 759.240 495.600 760.600 ;
        RECT 4.400 759.200 495.600 759.240 ;
        RECT 4.400 757.840 499.955 759.200 ;
        RECT 3.285 755.160 499.955 757.840 ;
        RECT 3.285 754.480 495.600 755.160 ;
        RECT 4.400 753.760 495.600 754.480 ;
        RECT 4.400 753.080 499.955 753.760 ;
        RECT 3.285 750.400 499.955 753.080 ;
        RECT 3.285 749.040 495.600 750.400 ;
        RECT 4.400 749.000 495.600 749.040 ;
        RECT 4.400 747.640 499.955 749.000 ;
        RECT 3.285 745.640 499.955 747.640 ;
        RECT 3.285 744.240 495.600 745.640 ;
        RECT 3.285 743.600 499.955 744.240 ;
        RECT 4.400 742.200 499.955 743.600 ;
        RECT 3.285 740.880 499.955 742.200 ;
        RECT 3.285 739.480 495.600 740.880 ;
        RECT 3.285 738.840 499.955 739.480 ;
        RECT 4.400 737.440 499.955 738.840 ;
        RECT 3.285 735.440 499.955 737.440 ;
        RECT 3.285 734.040 495.600 735.440 ;
        RECT 3.285 733.400 499.955 734.040 ;
        RECT 4.400 732.000 499.955 733.400 ;
        RECT 3.285 730.680 499.955 732.000 ;
        RECT 3.285 729.280 495.600 730.680 ;
        RECT 3.285 728.640 499.955 729.280 ;
        RECT 4.400 727.240 499.955 728.640 ;
        RECT 3.285 725.920 499.955 727.240 ;
        RECT 3.285 724.520 495.600 725.920 ;
        RECT 3.285 723.200 499.955 724.520 ;
        RECT 4.400 721.800 499.955 723.200 ;
        RECT 3.285 720.480 499.955 721.800 ;
        RECT 3.285 719.080 495.600 720.480 ;
        RECT 3.285 717.760 499.955 719.080 ;
        RECT 4.400 716.360 499.955 717.760 ;
        RECT 3.285 715.720 499.955 716.360 ;
        RECT 3.285 714.320 495.600 715.720 ;
        RECT 3.285 713.000 499.955 714.320 ;
        RECT 4.400 711.600 499.955 713.000 ;
        RECT 3.285 710.960 499.955 711.600 ;
        RECT 3.285 709.560 495.600 710.960 ;
        RECT 3.285 707.560 499.955 709.560 ;
        RECT 4.400 706.200 499.955 707.560 ;
        RECT 4.400 706.160 495.600 706.200 ;
        RECT 3.285 704.800 495.600 706.160 ;
        RECT 3.285 702.120 499.955 704.800 ;
        RECT 4.400 700.760 499.955 702.120 ;
        RECT 4.400 700.720 495.600 700.760 ;
        RECT 3.285 699.360 495.600 700.720 ;
        RECT 3.285 697.360 499.955 699.360 ;
        RECT 4.400 696.000 499.955 697.360 ;
        RECT 4.400 695.960 495.600 696.000 ;
        RECT 3.285 694.600 495.600 695.960 ;
        RECT 3.285 691.920 499.955 694.600 ;
        RECT 4.400 691.240 499.955 691.920 ;
        RECT 4.400 690.520 495.600 691.240 ;
        RECT 3.285 689.840 495.600 690.520 ;
        RECT 3.285 687.160 499.955 689.840 ;
        RECT 4.400 685.800 499.955 687.160 ;
        RECT 4.400 685.760 495.600 685.800 ;
        RECT 3.285 684.400 495.600 685.760 ;
        RECT 3.285 681.720 499.955 684.400 ;
        RECT 4.400 681.040 499.955 681.720 ;
        RECT 4.400 680.320 495.600 681.040 ;
        RECT 3.285 679.640 495.600 680.320 ;
        RECT 3.285 676.280 499.955 679.640 ;
        RECT 4.400 674.880 495.600 676.280 ;
        RECT 3.285 671.520 499.955 674.880 ;
        RECT 4.400 670.120 495.600 671.520 ;
        RECT 3.285 666.080 499.955 670.120 ;
        RECT 4.400 664.680 495.600 666.080 ;
        RECT 3.285 661.320 499.955 664.680 ;
        RECT 3.285 660.640 495.600 661.320 ;
        RECT 4.400 659.920 495.600 660.640 ;
        RECT 4.400 659.240 499.955 659.920 ;
        RECT 3.285 656.560 499.955 659.240 ;
        RECT 3.285 655.880 495.600 656.560 ;
        RECT 4.400 655.160 495.600 655.880 ;
        RECT 4.400 654.480 499.955 655.160 ;
        RECT 3.285 651.120 499.955 654.480 ;
        RECT 3.285 650.440 495.600 651.120 ;
        RECT 4.400 649.720 495.600 650.440 ;
        RECT 4.400 649.040 499.955 649.720 ;
        RECT 3.285 646.360 499.955 649.040 ;
        RECT 3.285 645.680 495.600 646.360 ;
        RECT 4.400 644.960 495.600 645.680 ;
        RECT 4.400 644.280 499.955 644.960 ;
        RECT 3.285 641.600 499.955 644.280 ;
        RECT 3.285 640.240 495.600 641.600 ;
        RECT 4.400 640.200 495.600 640.240 ;
        RECT 4.400 638.840 499.955 640.200 ;
        RECT 3.285 636.840 499.955 638.840 ;
        RECT 3.285 635.440 495.600 636.840 ;
        RECT 3.285 634.800 499.955 635.440 ;
        RECT 4.400 633.400 499.955 634.800 ;
        RECT 3.285 631.400 499.955 633.400 ;
        RECT 3.285 630.040 495.600 631.400 ;
        RECT 4.400 630.000 495.600 630.040 ;
        RECT 4.400 628.640 499.955 630.000 ;
        RECT 3.285 626.640 499.955 628.640 ;
        RECT 3.285 625.240 495.600 626.640 ;
        RECT 3.285 624.600 499.955 625.240 ;
        RECT 4.400 623.200 499.955 624.600 ;
        RECT 3.285 621.880 499.955 623.200 ;
        RECT 3.285 620.480 495.600 621.880 ;
        RECT 3.285 619.160 499.955 620.480 ;
        RECT 4.400 617.760 499.955 619.160 ;
        RECT 3.285 616.440 499.955 617.760 ;
        RECT 3.285 615.040 495.600 616.440 ;
        RECT 3.285 614.400 499.955 615.040 ;
        RECT 4.400 613.000 499.955 614.400 ;
        RECT 3.285 611.680 499.955 613.000 ;
        RECT 3.285 610.280 495.600 611.680 ;
        RECT 3.285 608.960 499.955 610.280 ;
        RECT 4.400 607.560 499.955 608.960 ;
        RECT 3.285 606.920 499.955 607.560 ;
        RECT 3.285 605.520 495.600 606.920 ;
        RECT 3.285 604.200 499.955 605.520 ;
        RECT 4.400 602.800 499.955 604.200 ;
        RECT 3.285 602.160 499.955 602.800 ;
        RECT 3.285 600.760 495.600 602.160 ;
        RECT 3.285 598.760 499.955 600.760 ;
        RECT 4.400 597.360 499.955 598.760 ;
        RECT 3.285 596.720 499.955 597.360 ;
        RECT 3.285 595.320 495.600 596.720 ;
        RECT 3.285 593.320 499.955 595.320 ;
        RECT 4.400 591.960 499.955 593.320 ;
        RECT 4.400 591.920 495.600 591.960 ;
        RECT 3.285 590.560 495.600 591.920 ;
        RECT 3.285 588.560 499.955 590.560 ;
        RECT 4.400 587.200 499.955 588.560 ;
        RECT 4.400 587.160 495.600 587.200 ;
        RECT 3.285 585.800 495.600 587.160 ;
        RECT 3.285 583.120 499.955 585.800 ;
        RECT 4.400 582.440 499.955 583.120 ;
        RECT 4.400 581.720 495.600 582.440 ;
        RECT 3.285 581.040 495.600 581.720 ;
        RECT 3.285 578.360 499.955 581.040 ;
        RECT 4.400 577.000 499.955 578.360 ;
        RECT 4.400 576.960 495.600 577.000 ;
        RECT 3.285 575.600 495.600 576.960 ;
        RECT 3.285 572.920 499.955 575.600 ;
        RECT 4.400 572.240 499.955 572.920 ;
        RECT 4.400 571.520 495.600 572.240 ;
        RECT 3.285 570.840 495.600 571.520 ;
        RECT 3.285 567.480 499.955 570.840 ;
        RECT 4.400 566.080 495.600 567.480 ;
        RECT 3.285 562.720 499.955 566.080 ;
        RECT 4.400 562.040 499.955 562.720 ;
        RECT 4.400 561.320 495.600 562.040 ;
        RECT 3.285 560.640 495.600 561.320 ;
        RECT 3.285 557.280 499.955 560.640 ;
        RECT 4.400 555.880 495.600 557.280 ;
        RECT 3.285 552.520 499.955 555.880 ;
        RECT 3.285 551.840 495.600 552.520 ;
        RECT 4.400 551.120 495.600 551.840 ;
        RECT 4.400 550.440 499.955 551.120 ;
        RECT 3.285 547.760 499.955 550.440 ;
        RECT 3.285 547.080 495.600 547.760 ;
        RECT 4.400 546.360 495.600 547.080 ;
        RECT 4.400 545.680 499.955 546.360 ;
        RECT 3.285 542.320 499.955 545.680 ;
        RECT 3.285 541.640 495.600 542.320 ;
        RECT 4.400 540.920 495.600 541.640 ;
        RECT 4.400 540.240 499.955 540.920 ;
        RECT 3.285 537.560 499.955 540.240 ;
        RECT 3.285 536.880 495.600 537.560 ;
        RECT 4.400 536.160 495.600 536.880 ;
        RECT 4.400 535.480 499.955 536.160 ;
        RECT 3.285 532.800 499.955 535.480 ;
        RECT 3.285 531.440 495.600 532.800 ;
        RECT 4.400 531.400 495.600 531.440 ;
        RECT 4.400 530.040 499.955 531.400 ;
        RECT 3.285 527.360 499.955 530.040 ;
        RECT 3.285 526.000 495.600 527.360 ;
        RECT 4.400 525.960 495.600 526.000 ;
        RECT 4.400 524.600 499.955 525.960 ;
        RECT 3.285 522.600 499.955 524.600 ;
        RECT 3.285 521.240 495.600 522.600 ;
        RECT 4.400 521.200 495.600 521.240 ;
        RECT 4.400 519.840 499.955 521.200 ;
        RECT 3.285 517.840 499.955 519.840 ;
        RECT 3.285 516.440 495.600 517.840 ;
        RECT 3.285 515.800 499.955 516.440 ;
        RECT 4.400 514.400 499.955 515.800 ;
        RECT 3.285 513.080 499.955 514.400 ;
        RECT 3.285 511.680 495.600 513.080 ;
        RECT 3.285 510.360 499.955 511.680 ;
        RECT 4.400 508.960 499.955 510.360 ;
        RECT 3.285 507.640 499.955 508.960 ;
        RECT 3.285 506.240 495.600 507.640 ;
        RECT 3.285 505.600 499.955 506.240 ;
        RECT 4.400 504.200 499.955 505.600 ;
        RECT 3.285 502.880 499.955 504.200 ;
        RECT 3.285 501.480 495.600 502.880 ;
        RECT 3.285 500.160 499.955 501.480 ;
        RECT 4.400 498.760 499.955 500.160 ;
        RECT 3.285 498.120 499.955 498.760 ;
        RECT 3.285 496.720 495.600 498.120 ;
        RECT 3.285 495.400 499.955 496.720 ;
        RECT 4.400 494.000 499.955 495.400 ;
        RECT 3.285 492.680 499.955 494.000 ;
        RECT 3.285 491.280 495.600 492.680 ;
        RECT 3.285 489.960 499.955 491.280 ;
        RECT 4.400 488.560 499.955 489.960 ;
        RECT 3.285 487.920 499.955 488.560 ;
        RECT 3.285 486.520 495.600 487.920 ;
        RECT 3.285 484.520 499.955 486.520 ;
        RECT 4.400 483.160 499.955 484.520 ;
        RECT 4.400 483.120 495.600 483.160 ;
        RECT 3.285 481.760 495.600 483.120 ;
        RECT 3.285 479.760 499.955 481.760 ;
        RECT 4.400 478.400 499.955 479.760 ;
        RECT 4.400 478.360 495.600 478.400 ;
        RECT 3.285 477.000 495.600 478.360 ;
        RECT 3.285 474.320 499.955 477.000 ;
        RECT 4.400 472.960 499.955 474.320 ;
        RECT 4.400 472.920 495.600 472.960 ;
        RECT 3.285 471.560 495.600 472.920 ;
        RECT 3.285 468.880 499.955 471.560 ;
        RECT 4.400 468.200 499.955 468.880 ;
        RECT 4.400 467.480 495.600 468.200 ;
        RECT 3.285 466.800 495.600 467.480 ;
        RECT 3.285 464.120 499.955 466.800 ;
        RECT 4.400 463.440 499.955 464.120 ;
        RECT 4.400 462.720 495.600 463.440 ;
        RECT 3.285 462.040 495.600 462.720 ;
        RECT 3.285 458.680 499.955 462.040 ;
        RECT 4.400 458.000 499.955 458.680 ;
        RECT 4.400 457.280 495.600 458.000 ;
        RECT 3.285 456.600 495.600 457.280 ;
        RECT 3.285 453.920 499.955 456.600 ;
        RECT 4.400 453.240 499.955 453.920 ;
        RECT 4.400 452.520 495.600 453.240 ;
        RECT 3.285 451.840 495.600 452.520 ;
        RECT 3.285 448.480 499.955 451.840 ;
        RECT 4.400 447.080 495.600 448.480 ;
        RECT 3.285 443.720 499.955 447.080 ;
        RECT 3.285 443.040 495.600 443.720 ;
        RECT 4.400 442.320 495.600 443.040 ;
        RECT 4.400 441.640 499.955 442.320 ;
        RECT 3.285 438.280 499.955 441.640 ;
        RECT 4.400 436.880 495.600 438.280 ;
        RECT 3.285 433.520 499.955 436.880 ;
        RECT 3.285 432.840 495.600 433.520 ;
        RECT 4.400 432.120 495.600 432.840 ;
        RECT 4.400 431.440 499.955 432.120 ;
        RECT 3.285 428.760 499.955 431.440 ;
        RECT 3.285 427.400 495.600 428.760 ;
        RECT 4.400 427.360 495.600 427.400 ;
        RECT 4.400 426.000 499.955 427.360 ;
        RECT 3.285 423.320 499.955 426.000 ;
        RECT 3.285 422.640 495.600 423.320 ;
        RECT 4.400 421.920 495.600 422.640 ;
        RECT 4.400 421.240 499.955 421.920 ;
        RECT 3.285 418.560 499.955 421.240 ;
        RECT 3.285 417.200 495.600 418.560 ;
        RECT 4.400 417.160 495.600 417.200 ;
        RECT 4.400 415.800 499.955 417.160 ;
        RECT 3.285 413.800 499.955 415.800 ;
        RECT 3.285 412.440 495.600 413.800 ;
        RECT 4.400 412.400 495.600 412.440 ;
        RECT 4.400 411.040 499.955 412.400 ;
        RECT 3.285 409.040 499.955 411.040 ;
        RECT 3.285 407.640 495.600 409.040 ;
        RECT 3.285 407.000 499.955 407.640 ;
        RECT 4.400 405.600 499.955 407.000 ;
        RECT 3.285 403.600 499.955 405.600 ;
        RECT 3.285 402.200 495.600 403.600 ;
        RECT 3.285 401.560 499.955 402.200 ;
        RECT 4.400 400.160 499.955 401.560 ;
        RECT 3.285 398.840 499.955 400.160 ;
        RECT 3.285 397.440 495.600 398.840 ;
        RECT 3.285 396.800 499.955 397.440 ;
        RECT 4.400 395.400 499.955 396.800 ;
        RECT 3.285 394.080 499.955 395.400 ;
        RECT 3.285 392.680 495.600 394.080 ;
        RECT 3.285 391.360 499.955 392.680 ;
        RECT 4.400 389.960 499.955 391.360 ;
        RECT 3.285 389.320 499.955 389.960 ;
        RECT 3.285 387.920 495.600 389.320 ;
        RECT 3.285 386.600 499.955 387.920 ;
        RECT 4.400 385.200 499.955 386.600 ;
        RECT 3.285 383.880 499.955 385.200 ;
        RECT 3.285 382.480 495.600 383.880 ;
        RECT 3.285 381.160 499.955 382.480 ;
        RECT 4.400 379.760 499.955 381.160 ;
        RECT 3.285 379.120 499.955 379.760 ;
        RECT 3.285 377.720 495.600 379.120 ;
        RECT 3.285 375.720 499.955 377.720 ;
        RECT 4.400 374.360 499.955 375.720 ;
        RECT 4.400 374.320 495.600 374.360 ;
        RECT 3.285 372.960 495.600 374.320 ;
        RECT 3.285 370.960 499.955 372.960 ;
        RECT 4.400 369.560 499.955 370.960 ;
        RECT 3.285 368.920 499.955 369.560 ;
        RECT 3.285 367.520 495.600 368.920 ;
        RECT 3.285 365.520 499.955 367.520 ;
        RECT 4.400 364.160 499.955 365.520 ;
        RECT 4.400 364.120 495.600 364.160 ;
        RECT 3.285 362.760 495.600 364.120 ;
        RECT 3.285 360.080 499.955 362.760 ;
        RECT 4.400 359.400 499.955 360.080 ;
        RECT 4.400 358.680 495.600 359.400 ;
        RECT 3.285 358.000 495.600 358.680 ;
        RECT 3.285 355.320 499.955 358.000 ;
        RECT 4.400 354.640 499.955 355.320 ;
        RECT 4.400 353.920 495.600 354.640 ;
        RECT 3.285 353.240 495.600 353.920 ;
        RECT 3.285 349.880 499.955 353.240 ;
        RECT 4.400 349.200 499.955 349.880 ;
        RECT 4.400 348.480 495.600 349.200 ;
        RECT 3.285 347.800 495.600 348.480 ;
        RECT 3.285 345.120 499.955 347.800 ;
        RECT 4.400 344.440 499.955 345.120 ;
        RECT 4.400 343.720 495.600 344.440 ;
        RECT 3.285 343.040 495.600 343.720 ;
        RECT 3.285 339.680 499.955 343.040 ;
        RECT 4.400 338.280 495.600 339.680 ;
        RECT 3.285 334.240 499.955 338.280 ;
        RECT 4.400 332.840 495.600 334.240 ;
        RECT 3.285 329.480 499.955 332.840 ;
        RECT 4.400 328.080 495.600 329.480 ;
        RECT 3.285 324.720 499.955 328.080 ;
        RECT 3.285 324.040 495.600 324.720 ;
        RECT 4.400 323.320 495.600 324.040 ;
        RECT 4.400 322.640 499.955 323.320 ;
        RECT 3.285 319.960 499.955 322.640 ;
        RECT 3.285 318.600 495.600 319.960 ;
        RECT 4.400 318.560 495.600 318.600 ;
        RECT 4.400 317.200 499.955 318.560 ;
        RECT 3.285 314.520 499.955 317.200 ;
        RECT 3.285 313.840 495.600 314.520 ;
        RECT 4.400 313.120 495.600 313.840 ;
        RECT 4.400 312.440 499.955 313.120 ;
        RECT 3.285 309.760 499.955 312.440 ;
        RECT 3.285 308.400 495.600 309.760 ;
        RECT 4.400 308.360 495.600 308.400 ;
        RECT 4.400 307.000 499.955 308.360 ;
        RECT 3.285 305.000 499.955 307.000 ;
        RECT 3.285 303.640 495.600 305.000 ;
        RECT 4.400 303.600 495.600 303.640 ;
        RECT 4.400 302.240 499.955 303.600 ;
        RECT 3.285 299.560 499.955 302.240 ;
        RECT 3.285 298.200 495.600 299.560 ;
        RECT 4.400 298.160 495.600 298.200 ;
        RECT 4.400 296.800 499.955 298.160 ;
        RECT 3.285 294.800 499.955 296.800 ;
        RECT 3.285 293.400 495.600 294.800 ;
        RECT 3.285 292.760 499.955 293.400 ;
        RECT 4.400 291.360 499.955 292.760 ;
        RECT 3.285 290.040 499.955 291.360 ;
        RECT 3.285 288.640 495.600 290.040 ;
        RECT 3.285 288.000 499.955 288.640 ;
        RECT 4.400 286.600 499.955 288.000 ;
        RECT 3.285 285.280 499.955 286.600 ;
        RECT 3.285 283.880 495.600 285.280 ;
        RECT 3.285 282.560 499.955 283.880 ;
        RECT 4.400 281.160 499.955 282.560 ;
        RECT 3.285 279.840 499.955 281.160 ;
        RECT 3.285 278.440 495.600 279.840 ;
        RECT 3.285 277.120 499.955 278.440 ;
        RECT 4.400 275.720 499.955 277.120 ;
        RECT 3.285 275.080 499.955 275.720 ;
        RECT 3.285 273.680 495.600 275.080 ;
        RECT 3.285 272.360 499.955 273.680 ;
        RECT 4.400 270.960 499.955 272.360 ;
        RECT 3.285 270.320 499.955 270.960 ;
        RECT 3.285 268.920 495.600 270.320 ;
        RECT 3.285 266.920 499.955 268.920 ;
        RECT 4.400 265.520 499.955 266.920 ;
        RECT 3.285 264.880 499.955 265.520 ;
        RECT 3.285 263.480 495.600 264.880 ;
        RECT 3.285 262.160 499.955 263.480 ;
        RECT 4.400 260.760 499.955 262.160 ;
        RECT 3.285 260.120 499.955 260.760 ;
        RECT 3.285 258.720 495.600 260.120 ;
        RECT 3.285 256.720 499.955 258.720 ;
        RECT 4.400 255.360 499.955 256.720 ;
        RECT 4.400 255.320 495.600 255.360 ;
        RECT 3.285 253.960 495.600 255.320 ;
        RECT 3.285 251.280 499.955 253.960 ;
        RECT 4.400 250.600 499.955 251.280 ;
        RECT 4.400 249.880 495.600 250.600 ;
        RECT 3.285 249.200 495.600 249.880 ;
        RECT 3.285 246.520 499.955 249.200 ;
        RECT 4.400 245.160 499.955 246.520 ;
        RECT 4.400 245.120 495.600 245.160 ;
        RECT 3.285 243.760 495.600 245.120 ;
        RECT 3.285 241.080 499.955 243.760 ;
        RECT 4.400 240.400 499.955 241.080 ;
        RECT 4.400 239.680 495.600 240.400 ;
        RECT 3.285 239.000 495.600 239.680 ;
        RECT 3.285 235.640 499.955 239.000 ;
        RECT 4.400 234.240 495.600 235.640 ;
        RECT 3.285 230.880 499.955 234.240 ;
        RECT 4.400 230.200 499.955 230.880 ;
        RECT 4.400 229.480 495.600 230.200 ;
        RECT 3.285 228.800 495.600 229.480 ;
        RECT 3.285 225.440 499.955 228.800 ;
        RECT 4.400 224.040 495.600 225.440 ;
        RECT 3.285 220.680 499.955 224.040 ;
        RECT 4.400 219.280 495.600 220.680 ;
        RECT 3.285 215.920 499.955 219.280 ;
        RECT 3.285 215.240 495.600 215.920 ;
        RECT 4.400 214.520 495.600 215.240 ;
        RECT 4.400 213.840 499.955 214.520 ;
        RECT 3.285 210.480 499.955 213.840 ;
        RECT 3.285 209.800 495.600 210.480 ;
        RECT 4.400 209.080 495.600 209.800 ;
        RECT 4.400 208.400 499.955 209.080 ;
        RECT 3.285 205.720 499.955 208.400 ;
        RECT 3.285 205.040 495.600 205.720 ;
        RECT 4.400 204.320 495.600 205.040 ;
        RECT 4.400 203.640 499.955 204.320 ;
        RECT 3.285 200.960 499.955 203.640 ;
        RECT 3.285 199.600 495.600 200.960 ;
        RECT 4.400 199.560 495.600 199.600 ;
        RECT 4.400 198.200 499.955 199.560 ;
        RECT 3.285 196.200 499.955 198.200 ;
        RECT 3.285 194.840 495.600 196.200 ;
        RECT 4.400 194.800 495.600 194.840 ;
        RECT 4.400 193.440 499.955 194.800 ;
        RECT 3.285 190.760 499.955 193.440 ;
        RECT 3.285 189.400 495.600 190.760 ;
        RECT 4.400 189.360 495.600 189.400 ;
        RECT 4.400 188.000 499.955 189.360 ;
        RECT 3.285 186.000 499.955 188.000 ;
        RECT 3.285 184.600 495.600 186.000 ;
        RECT 3.285 183.960 499.955 184.600 ;
        RECT 4.400 182.560 499.955 183.960 ;
        RECT 3.285 181.240 499.955 182.560 ;
        RECT 3.285 179.840 495.600 181.240 ;
        RECT 3.285 179.200 499.955 179.840 ;
        RECT 4.400 177.800 499.955 179.200 ;
        RECT 3.285 175.800 499.955 177.800 ;
        RECT 3.285 174.400 495.600 175.800 ;
        RECT 3.285 173.760 499.955 174.400 ;
        RECT 4.400 172.360 499.955 173.760 ;
        RECT 3.285 171.040 499.955 172.360 ;
        RECT 3.285 169.640 495.600 171.040 ;
        RECT 3.285 168.320 499.955 169.640 ;
        RECT 4.400 166.920 499.955 168.320 ;
        RECT 3.285 166.280 499.955 166.920 ;
        RECT 3.285 164.880 495.600 166.280 ;
        RECT 3.285 163.560 499.955 164.880 ;
        RECT 4.400 162.160 499.955 163.560 ;
        RECT 3.285 161.520 499.955 162.160 ;
        RECT 3.285 160.120 495.600 161.520 ;
        RECT 3.285 158.120 499.955 160.120 ;
        RECT 4.400 156.720 499.955 158.120 ;
        RECT 3.285 156.080 499.955 156.720 ;
        RECT 3.285 154.680 495.600 156.080 ;
        RECT 3.285 153.360 499.955 154.680 ;
        RECT 4.400 151.960 499.955 153.360 ;
        RECT 3.285 151.320 499.955 151.960 ;
        RECT 3.285 149.920 495.600 151.320 ;
        RECT 3.285 147.920 499.955 149.920 ;
        RECT 4.400 146.560 499.955 147.920 ;
        RECT 4.400 146.520 495.600 146.560 ;
        RECT 3.285 145.160 495.600 146.520 ;
        RECT 3.285 142.480 499.955 145.160 ;
        RECT 4.400 141.120 499.955 142.480 ;
        RECT 4.400 141.080 495.600 141.120 ;
        RECT 3.285 139.720 495.600 141.080 ;
        RECT 3.285 137.720 499.955 139.720 ;
        RECT 4.400 136.360 499.955 137.720 ;
        RECT 4.400 136.320 495.600 136.360 ;
        RECT 3.285 134.960 495.600 136.320 ;
        RECT 3.285 132.280 499.955 134.960 ;
        RECT 4.400 131.600 499.955 132.280 ;
        RECT 4.400 130.880 495.600 131.600 ;
        RECT 3.285 130.200 495.600 130.880 ;
        RECT 3.285 126.840 499.955 130.200 ;
        RECT 4.400 125.440 495.600 126.840 ;
        RECT 3.285 122.080 499.955 125.440 ;
        RECT 4.400 121.400 499.955 122.080 ;
        RECT 4.400 120.680 495.600 121.400 ;
        RECT 3.285 120.000 495.600 120.680 ;
        RECT 3.285 116.640 499.955 120.000 ;
        RECT 4.400 115.240 495.600 116.640 ;
        RECT 3.285 111.880 499.955 115.240 ;
        RECT 4.400 110.480 495.600 111.880 ;
        RECT 3.285 106.440 499.955 110.480 ;
        RECT 4.400 105.040 495.600 106.440 ;
        RECT 3.285 101.680 499.955 105.040 ;
        RECT 3.285 101.000 495.600 101.680 ;
        RECT 4.400 100.280 495.600 101.000 ;
        RECT 4.400 99.600 499.955 100.280 ;
        RECT 3.285 96.920 499.955 99.600 ;
        RECT 3.285 96.240 495.600 96.920 ;
        RECT 4.400 95.520 495.600 96.240 ;
        RECT 4.400 94.840 499.955 95.520 ;
        RECT 3.285 92.160 499.955 94.840 ;
        RECT 3.285 90.800 495.600 92.160 ;
        RECT 4.400 90.760 495.600 90.800 ;
        RECT 4.400 89.400 499.955 90.760 ;
        RECT 3.285 86.720 499.955 89.400 ;
        RECT 3.285 85.360 495.600 86.720 ;
        RECT 4.400 85.320 495.600 85.360 ;
        RECT 4.400 83.960 499.955 85.320 ;
        RECT 3.285 81.960 499.955 83.960 ;
        RECT 3.285 80.600 495.600 81.960 ;
        RECT 4.400 80.560 495.600 80.600 ;
        RECT 4.400 79.200 499.955 80.560 ;
        RECT 3.285 77.200 499.955 79.200 ;
        RECT 3.285 75.800 495.600 77.200 ;
        RECT 3.285 75.160 499.955 75.800 ;
        RECT 4.400 73.760 499.955 75.160 ;
        RECT 3.285 71.760 499.955 73.760 ;
        RECT 3.285 70.400 495.600 71.760 ;
        RECT 4.400 70.360 495.600 70.400 ;
        RECT 4.400 69.000 499.955 70.360 ;
        RECT 3.285 67.000 499.955 69.000 ;
        RECT 3.285 65.600 495.600 67.000 ;
        RECT 3.285 64.960 499.955 65.600 ;
        RECT 4.400 63.560 499.955 64.960 ;
        RECT 3.285 62.240 499.955 63.560 ;
        RECT 3.285 60.840 495.600 62.240 ;
        RECT 3.285 59.520 499.955 60.840 ;
        RECT 4.400 58.120 499.955 59.520 ;
        RECT 3.285 57.480 499.955 58.120 ;
        RECT 3.285 56.080 495.600 57.480 ;
        RECT 3.285 54.760 499.955 56.080 ;
        RECT 4.400 53.360 499.955 54.760 ;
        RECT 3.285 52.040 499.955 53.360 ;
        RECT 3.285 50.640 495.600 52.040 ;
        RECT 3.285 49.320 499.955 50.640 ;
        RECT 4.400 47.920 499.955 49.320 ;
        RECT 3.285 47.280 499.955 47.920 ;
        RECT 3.285 45.880 495.600 47.280 ;
        RECT 3.285 43.880 499.955 45.880 ;
        RECT 4.400 42.520 499.955 43.880 ;
        RECT 4.400 42.480 495.600 42.520 ;
        RECT 3.285 41.120 495.600 42.480 ;
        RECT 3.285 39.120 499.955 41.120 ;
        RECT 4.400 37.720 499.955 39.120 ;
        RECT 3.285 37.080 499.955 37.720 ;
        RECT 3.285 35.680 495.600 37.080 ;
        RECT 3.285 33.680 499.955 35.680 ;
        RECT 4.400 32.320 499.955 33.680 ;
        RECT 4.400 32.280 495.600 32.320 ;
        RECT 3.285 30.920 495.600 32.280 ;
        RECT 3.285 28.920 499.955 30.920 ;
        RECT 4.400 27.560 499.955 28.920 ;
        RECT 4.400 27.520 495.600 27.560 ;
        RECT 3.285 26.160 495.600 27.520 ;
        RECT 3.285 23.480 499.955 26.160 ;
        RECT 4.400 22.800 499.955 23.480 ;
        RECT 4.400 22.080 495.600 22.800 ;
        RECT 3.285 21.400 495.600 22.080 ;
        RECT 3.285 18.040 499.955 21.400 ;
        RECT 4.400 17.360 499.955 18.040 ;
        RECT 4.400 16.640 495.600 17.360 ;
        RECT 3.285 15.960 495.600 16.640 ;
        RECT 3.285 13.280 499.955 15.960 ;
        RECT 4.400 12.600 499.955 13.280 ;
        RECT 4.400 11.880 495.600 12.600 ;
        RECT 3.285 11.200 495.600 11.880 ;
        RECT 3.285 7.840 499.955 11.200 ;
        RECT 4.400 6.440 495.600 7.840 ;
        RECT 3.285 3.080 499.955 6.440 ;
        RECT 4.400 2.215 495.600 3.080 ;
      LAYER met4 ;
        RECT 7.655 34.175 20.640 925.305 ;
        RECT 23.040 34.175 97.440 925.305 ;
        RECT 99.840 34.175 174.240 925.305 ;
        RECT 176.640 34.175 251.040 925.305 ;
        RECT 253.440 34.175 327.840 925.305 ;
        RECT 330.240 34.175 404.640 925.305 ;
        RECT 407.040 34.175 481.440 925.305 ;
        RECT 483.840 34.175 499.265 925.305 ;
  END
END ExperiarCore
END LIBRARY

