magic
tech sky130A
magscale 1 2
timestamp 1653402246
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 290 1708 69630 67584
<< metal2 >>
rect 294 69200 350 70000
rect 938 69200 994 70000
rect 1582 69200 1638 70000
rect 2318 69200 2374 70000
rect 2962 69200 3018 70000
rect 3698 69200 3754 70000
rect 4342 69200 4398 70000
rect 5078 69200 5134 70000
rect 5722 69200 5778 70000
rect 6458 69200 6514 70000
rect 7102 69200 7158 70000
rect 7838 69200 7894 70000
rect 8482 69200 8538 70000
rect 9126 69200 9182 70000
rect 9862 69200 9918 70000
rect 10506 69200 10562 70000
rect 11242 69200 11298 70000
rect 11886 69200 11942 70000
rect 12622 69200 12678 70000
rect 13266 69200 13322 70000
rect 14002 69200 14058 70000
rect 14646 69200 14702 70000
rect 15382 69200 15438 70000
rect 16026 69200 16082 70000
rect 16762 69200 16818 70000
rect 17406 69200 17462 70000
rect 18050 69200 18106 70000
rect 18786 69200 18842 70000
rect 19430 69200 19486 70000
rect 20166 69200 20222 70000
rect 20810 69200 20866 70000
rect 21546 69200 21602 70000
rect 22190 69200 22246 70000
rect 22926 69200 22982 70000
rect 23570 69200 23626 70000
rect 24306 69200 24362 70000
rect 24950 69200 25006 70000
rect 25686 69200 25742 70000
rect 26330 69200 26386 70000
rect 26974 69200 27030 70000
rect 27710 69200 27766 70000
rect 28354 69200 28410 70000
rect 29090 69200 29146 70000
rect 29734 69200 29790 70000
rect 30470 69200 30526 70000
rect 31114 69200 31170 70000
rect 31850 69200 31906 70000
rect 32494 69200 32550 70000
rect 33230 69200 33286 70000
rect 33874 69200 33930 70000
rect 34610 69200 34666 70000
rect 35254 69200 35310 70000
rect 35898 69200 35954 70000
rect 36634 69200 36690 70000
rect 37278 69200 37334 70000
rect 38014 69200 38070 70000
rect 38658 69200 38714 70000
rect 39394 69200 39450 70000
rect 40038 69200 40094 70000
rect 40774 69200 40830 70000
rect 41418 69200 41474 70000
rect 42154 69200 42210 70000
rect 42798 69200 42854 70000
rect 43534 69200 43590 70000
rect 44178 69200 44234 70000
rect 44822 69200 44878 70000
rect 45558 69200 45614 70000
rect 46202 69200 46258 70000
rect 46938 69200 46994 70000
rect 47582 69200 47638 70000
rect 48318 69200 48374 70000
rect 48962 69200 49018 70000
rect 49698 69200 49754 70000
rect 50342 69200 50398 70000
rect 51078 69200 51134 70000
rect 51722 69200 51778 70000
rect 52458 69200 52514 70000
rect 53102 69200 53158 70000
rect 53746 69200 53802 70000
rect 54482 69200 54538 70000
rect 55126 69200 55182 70000
rect 55862 69200 55918 70000
rect 56506 69200 56562 70000
rect 57242 69200 57298 70000
rect 57886 69200 57942 70000
rect 58622 69200 58678 70000
rect 59266 69200 59322 70000
rect 60002 69200 60058 70000
rect 60646 69200 60702 70000
rect 61382 69200 61438 70000
rect 62026 69200 62082 70000
rect 62670 69200 62726 70000
rect 63406 69200 63462 70000
rect 64050 69200 64106 70000
rect 64786 69200 64842 70000
rect 65430 69200 65486 70000
rect 66166 69200 66222 70000
rect 66810 69200 66866 70000
rect 67546 69200 67602 70000
rect 68190 69200 68246 70000
rect 68926 69200 68982 70000
rect 69570 69200 69626 70000
rect 294 0 350 800
rect 938 0 994 800
rect 1582 0 1638 800
rect 2226 0 2282 800
rect 2870 0 2926 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 4894 0 4950 800
rect 5538 0 5594 800
rect 6182 0 6238 800
rect 6826 0 6882 800
rect 7470 0 7526 800
rect 8206 0 8262 800
rect 8850 0 8906 800
rect 9494 0 9550 800
rect 10138 0 10194 800
rect 10782 0 10838 800
rect 11518 0 11574 800
rect 12162 0 12218 800
rect 12806 0 12862 800
rect 13450 0 13506 800
rect 14094 0 14150 800
rect 14738 0 14794 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18786 0 18842 800
rect 19430 0 19486 800
rect 20074 0 20130 800
rect 20718 0 20774 800
rect 21362 0 21418 800
rect 22006 0 22062 800
rect 22742 0 22798 800
rect 23386 0 23442 800
rect 24030 0 24086 800
rect 24674 0 24730 800
rect 25318 0 25374 800
rect 25962 0 26018 800
rect 26698 0 26754 800
rect 27342 0 27398 800
rect 27986 0 28042 800
rect 28630 0 28686 800
rect 29274 0 29330 800
rect 30010 0 30066 800
rect 30654 0 30710 800
rect 31298 0 31354 800
rect 31942 0 31998 800
rect 32586 0 32642 800
rect 33230 0 33286 800
rect 33966 0 34022 800
rect 34610 0 34666 800
rect 35254 0 35310 800
rect 35898 0 35954 800
rect 36542 0 36598 800
rect 37278 0 37334 800
rect 37922 0 37978 800
rect 38566 0 38622 800
rect 39210 0 39266 800
rect 39854 0 39910 800
rect 40498 0 40554 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44546 0 44602 800
rect 45190 0 45246 800
rect 45834 0 45890 800
rect 46478 0 46534 800
rect 47122 0 47178 800
rect 47766 0 47822 800
rect 48502 0 48558 800
rect 49146 0 49202 800
rect 49790 0 49846 800
rect 50434 0 50490 800
rect 51078 0 51134 800
rect 51722 0 51778 800
rect 52458 0 52514 800
rect 53102 0 53158 800
rect 53746 0 53802 800
rect 54390 0 54446 800
rect 55034 0 55090 800
rect 55770 0 55826 800
rect 56414 0 56470 800
rect 57058 0 57114 800
rect 57702 0 57758 800
rect 58346 0 58402 800
rect 58990 0 59046 800
rect 59726 0 59782 800
rect 60370 0 60426 800
rect 61014 0 61070 800
rect 61658 0 61714 800
rect 62302 0 62358 800
rect 63038 0 63094 800
rect 63682 0 63738 800
rect 64326 0 64382 800
rect 64970 0 65026 800
rect 65614 0 65670 800
rect 66258 0 66314 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
<< obsm2 >>
rect 18 69144 238 69306
rect 406 69144 882 69306
rect 1050 69144 1526 69306
rect 1694 69144 2262 69306
rect 2430 69144 2906 69306
rect 3074 69144 3642 69306
rect 3810 69144 4286 69306
rect 4454 69144 5022 69306
rect 5190 69144 5666 69306
rect 5834 69144 6402 69306
rect 6570 69144 7046 69306
rect 7214 69144 7782 69306
rect 7950 69144 8426 69306
rect 8594 69144 9070 69306
rect 9238 69144 9806 69306
rect 9974 69144 10450 69306
rect 10618 69144 11186 69306
rect 11354 69144 11830 69306
rect 11998 69144 12566 69306
rect 12734 69144 13210 69306
rect 13378 69144 13946 69306
rect 14114 69144 14590 69306
rect 14758 69144 15326 69306
rect 15494 69144 15970 69306
rect 16138 69144 16706 69306
rect 16874 69144 17350 69306
rect 17518 69144 17994 69306
rect 18162 69144 18730 69306
rect 18898 69144 19374 69306
rect 19542 69144 20110 69306
rect 20278 69144 20754 69306
rect 20922 69144 21490 69306
rect 21658 69144 22134 69306
rect 22302 69144 22870 69306
rect 23038 69144 23514 69306
rect 23682 69144 24250 69306
rect 24418 69144 24894 69306
rect 25062 69144 25630 69306
rect 25798 69144 26274 69306
rect 26442 69144 26918 69306
rect 27086 69144 27654 69306
rect 27822 69144 28298 69306
rect 28466 69144 29034 69306
rect 29202 69144 29678 69306
rect 29846 69144 30414 69306
rect 30582 69144 31058 69306
rect 31226 69144 31794 69306
rect 31962 69144 32438 69306
rect 32606 69144 33174 69306
rect 33342 69144 33818 69306
rect 33986 69144 34554 69306
rect 34722 69144 35198 69306
rect 35366 69144 35842 69306
rect 36010 69144 36578 69306
rect 36746 69144 37222 69306
rect 37390 69144 37958 69306
rect 38126 69144 38602 69306
rect 38770 69144 39338 69306
rect 39506 69144 39982 69306
rect 40150 69144 40718 69306
rect 40886 69144 41362 69306
rect 41530 69144 42098 69306
rect 42266 69144 42742 69306
rect 42910 69144 43478 69306
rect 43646 69144 44122 69306
rect 44290 69144 44766 69306
rect 44934 69144 45502 69306
rect 45670 69144 46146 69306
rect 46314 69144 46882 69306
rect 47050 69144 47526 69306
rect 47694 69144 48262 69306
rect 48430 69144 48906 69306
rect 49074 69144 49642 69306
rect 49810 69144 50286 69306
rect 50454 69144 51022 69306
rect 51190 69144 51666 69306
rect 51834 69144 52402 69306
rect 52570 69144 53046 69306
rect 53214 69144 53690 69306
rect 53858 69144 54426 69306
rect 54594 69144 55070 69306
rect 55238 69144 55806 69306
rect 55974 69144 56450 69306
rect 56618 69144 57186 69306
rect 57354 69144 57830 69306
rect 57998 69144 58566 69306
rect 58734 69144 59210 69306
rect 59378 69144 59946 69306
rect 60114 69144 60590 69306
rect 60758 69144 61326 69306
rect 61494 69144 61970 69306
rect 62138 69144 62614 69306
rect 62782 69144 63350 69306
rect 63518 69144 63994 69306
rect 64162 69144 64730 69306
rect 64898 69144 65374 69306
rect 65542 69144 66110 69306
rect 66278 69144 66754 69306
rect 66922 69144 67490 69306
rect 67658 69144 68134 69306
rect 68302 69144 68870 69306
rect 69038 69144 69514 69306
rect 18 856 69624 69144
rect 18 734 238 856
rect 406 734 882 856
rect 1050 734 1526 856
rect 1694 734 2170 856
rect 2338 734 2814 856
rect 2982 734 3458 856
rect 3626 734 4194 856
rect 4362 734 4838 856
rect 5006 734 5482 856
rect 5650 734 6126 856
rect 6294 734 6770 856
rect 6938 734 7414 856
rect 7582 734 8150 856
rect 8318 734 8794 856
rect 8962 734 9438 856
rect 9606 734 10082 856
rect 10250 734 10726 856
rect 10894 734 11462 856
rect 11630 734 12106 856
rect 12274 734 12750 856
rect 12918 734 13394 856
rect 13562 734 14038 856
rect 14206 734 14682 856
rect 14850 734 15418 856
rect 15586 734 16062 856
rect 16230 734 16706 856
rect 16874 734 17350 856
rect 17518 734 17994 856
rect 18162 734 18730 856
rect 18898 734 19374 856
rect 19542 734 20018 856
rect 20186 734 20662 856
rect 20830 734 21306 856
rect 21474 734 21950 856
rect 22118 734 22686 856
rect 22854 734 23330 856
rect 23498 734 23974 856
rect 24142 734 24618 856
rect 24786 734 25262 856
rect 25430 734 25906 856
rect 26074 734 26642 856
rect 26810 734 27286 856
rect 27454 734 27930 856
rect 28098 734 28574 856
rect 28742 734 29218 856
rect 29386 734 29954 856
rect 30122 734 30598 856
rect 30766 734 31242 856
rect 31410 734 31886 856
rect 32054 734 32530 856
rect 32698 734 33174 856
rect 33342 734 33910 856
rect 34078 734 34554 856
rect 34722 734 35198 856
rect 35366 734 35842 856
rect 36010 734 36486 856
rect 36654 734 37222 856
rect 37390 734 37866 856
rect 38034 734 38510 856
rect 38678 734 39154 856
rect 39322 734 39798 856
rect 39966 734 40442 856
rect 40610 734 41178 856
rect 41346 734 41822 856
rect 41990 734 42466 856
rect 42634 734 43110 856
rect 43278 734 43754 856
rect 43922 734 44490 856
rect 44658 734 45134 856
rect 45302 734 45778 856
rect 45946 734 46422 856
rect 46590 734 47066 856
rect 47234 734 47710 856
rect 47878 734 48446 856
rect 48614 734 49090 856
rect 49258 734 49734 856
rect 49902 734 50378 856
rect 50546 734 51022 856
rect 51190 734 51666 856
rect 51834 734 52402 856
rect 52570 734 53046 856
rect 53214 734 53690 856
rect 53858 734 54334 856
rect 54502 734 54978 856
rect 55146 734 55714 856
rect 55882 734 56358 856
rect 56526 734 57002 856
rect 57170 734 57646 856
rect 57814 734 58290 856
rect 58458 734 58934 856
rect 59102 734 59670 856
rect 59838 734 60314 856
rect 60482 734 60958 856
rect 61126 734 61602 856
rect 61770 734 62246 856
rect 62414 734 62982 856
rect 63150 734 63626 856
rect 63794 734 64270 856
rect 64438 734 64914 856
rect 65082 734 65558 856
rect 65726 734 66202 856
rect 66370 734 66938 856
rect 67106 734 67582 856
rect 67750 734 68226 856
rect 68394 734 68870 856
rect 69038 734 69514 856
<< metal3 >>
rect 0 69232 800 69352
rect 0 67736 800 67856
rect 0 66240 800 66360
rect 0 64744 800 64864
rect 0 63248 800 63368
rect 0 61752 800 61872
rect 0 60256 800 60376
rect 0 58760 800 58880
rect 0 57264 800 57384
rect 0 55768 800 55888
rect 0 54272 800 54392
rect 0 52776 800 52896
rect 69200 52368 70000 52488
rect 0 51280 800 51400
rect 0 49784 800 49904
rect 0 48288 800 48408
rect 0 46792 800 46912
rect 0 45296 800 45416
rect 0 43800 800 43920
rect 0 42304 800 42424
rect 0 40808 800 40928
rect 0 39312 800 39432
rect 0 37816 800 37936
rect 0 36320 800 36440
rect 0 34960 800 35080
rect 0 33464 800 33584
rect 0 31968 800 32088
rect 0 30472 800 30592
rect 0 28976 800 29096
rect 0 27480 800 27600
rect 0 25984 800 26104
rect 0 24488 800 24608
rect 0 22992 800 23112
rect 0 21496 800 21616
rect 0 20000 800 20120
rect 0 18504 800 18624
rect 69200 17416 70000 17536
rect 0 17008 800 17128
rect 0 15512 800 15632
rect 0 14016 800 14136
rect 0 12520 800 12640
rect 0 11024 800 11144
rect 0 9528 800 9648
rect 0 8032 800 8152
rect 0 6536 800 6656
rect 0 5040 800 5160
rect 0 3544 800 3664
rect 0 2048 800 2168
rect 0 688 800 808
<< obsm3 >>
rect 880 69152 69200 69322
rect 13 67936 69200 69152
rect 880 67656 69200 67936
rect 13 66440 69200 67656
rect 880 66160 69200 66440
rect 13 64944 69200 66160
rect 880 64664 69200 64944
rect 13 63448 69200 64664
rect 880 63168 69200 63448
rect 13 61952 69200 63168
rect 880 61672 69200 61952
rect 13 60456 69200 61672
rect 880 60176 69200 60456
rect 13 58960 69200 60176
rect 880 58680 69200 58960
rect 13 57464 69200 58680
rect 880 57184 69200 57464
rect 13 55968 69200 57184
rect 880 55688 69200 55968
rect 13 54472 69200 55688
rect 880 54192 69200 54472
rect 13 52976 69200 54192
rect 880 52696 69200 52976
rect 13 52568 69200 52696
rect 13 52288 69120 52568
rect 13 51480 69200 52288
rect 880 51200 69200 51480
rect 13 49984 69200 51200
rect 880 49704 69200 49984
rect 13 48488 69200 49704
rect 880 48208 69200 48488
rect 13 46992 69200 48208
rect 880 46712 69200 46992
rect 13 45496 69200 46712
rect 880 45216 69200 45496
rect 13 44000 69200 45216
rect 880 43720 69200 44000
rect 13 42504 69200 43720
rect 880 42224 69200 42504
rect 13 41008 69200 42224
rect 880 40728 69200 41008
rect 13 39512 69200 40728
rect 880 39232 69200 39512
rect 13 38016 69200 39232
rect 880 37736 69200 38016
rect 13 36520 69200 37736
rect 880 36240 69200 36520
rect 13 35160 69200 36240
rect 880 34880 69200 35160
rect 13 33664 69200 34880
rect 880 33384 69200 33664
rect 13 32168 69200 33384
rect 880 31888 69200 32168
rect 13 30672 69200 31888
rect 880 30392 69200 30672
rect 13 29176 69200 30392
rect 880 28896 69200 29176
rect 13 27680 69200 28896
rect 880 27400 69200 27680
rect 13 26184 69200 27400
rect 880 25904 69200 26184
rect 13 24688 69200 25904
rect 880 24408 69200 24688
rect 13 23192 69200 24408
rect 880 22912 69200 23192
rect 13 21696 69200 22912
rect 880 21416 69200 21696
rect 13 20200 69200 21416
rect 880 19920 69200 20200
rect 13 18704 69200 19920
rect 880 18424 69200 18704
rect 13 17616 69200 18424
rect 13 17336 69120 17616
rect 13 17208 69200 17336
rect 880 16928 69200 17208
rect 13 15712 69200 16928
rect 880 15432 69200 15712
rect 13 14216 69200 15432
rect 880 13936 69200 14216
rect 13 12720 69200 13936
rect 880 12440 69200 12720
rect 13 11224 69200 12440
rect 880 10944 69200 11224
rect 13 9728 69200 10944
rect 880 9448 69200 9728
rect 13 8232 69200 9448
rect 880 7952 69200 8232
rect 13 6736 69200 7952
rect 880 6456 69200 6736
rect 13 5240 69200 6456
rect 880 4960 69200 5240
rect 13 3744 69200 4960
rect 880 3464 69200 3744
rect 13 2248 69200 3464
rect 880 1968 69200 2248
rect 13 888 69200 1968
rect 880 718 69200 888
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< obsm4 >>
rect 6315 2483 19488 66605
rect 19968 2483 34848 66605
rect 35328 2483 50208 66605
rect 50688 2483 64157 66605
<< labels >>
rlabel metal3 s 69200 17416 70000 17536 6 caravel_uart_rx
port 1 nsew signal input
rlabel metal3 s 69200 52368 70000 52488 6 caravel_uart_tx
port 2 nsew signal output
rlabel metal2 s 294 69200 350 70000 6 caravel_wb_ack_i
port 3 nsew signal input
rlabel metal2 s 4342 69200 4398 70000 6 caravel_wb_adr_o[0]
port 4 nsew signal output
rlabel metal2 s 27710 69200 27766 70000 6 caravel_wb_adr_o[10]
port 5 nsew signal output
rlabel metal2 s 29734 69200 29790 70000 6 caravel_wb_adr_o[11]
port 6 nsew signal output
rlabel metal2 s 31850 69200 31906 70000 6 caravel_wb_adr_o[12]
port 7 nsew signal output
rlabel metal2 s 33874 69200 33930 70000 6 caravel_wb_adr_o[13]
port 8 nsew signal output
rlabel metal2 s 35898 69200 35954 70000 6 caravel_wb_adr_o[14]
port 9 nsew signal output
rlabel metal2 s 38014 69200 38070 70000 6 caravel_wb_adr_o[15]
port 10 nsew signal output
rlabel metal2 s 40038 69200 40094 70000 6 caravel_wb_adr_o[16]
port 11 nsew signal output
rlabel metal2 s 42154 69200 42210 70000 6 caravel_wb_adr_o[17]
port 12 nsew signal output
rlabel metal2 s 44178 69200 44234 70000 6 caravel_wb_adr_o[18]
port 13 nsew signal output
rlabel metal2 s 46202 69200 46258 70000 6 caravel_wb_adr_o[19]
port 14 nsew signal output
rlabel metal2 s 7102 69200 7158 70000 6 caravel_wb_adr_o[1]
port 15 nsew signal output
rlabel metal2 s 48318 69200 48374 70000 6 caravel_wb_adr_o[20]
port 16 nsew signal output
rlabel metal2 s 50342 69200 50398 70000 6 caravel_wb_adr_o[21]
port 17 nsew signal output
rlabel metal2 s 52458 69200 52514 70000 6 caravel_wb_adr_o[22]
port 18 nsew signal output
rlabel metal2 s 54482 69200 54538 70000 6 caravel_wb_adr_o[23]
port 19 nsew signal output
rlabel metal2 s 56506 69200 56562 70000 6 caravel_wb_adr_o[24]
port 20 nsew signal output
rlabel metal2 s 58622 69200 58678 70000 6 caravel_wb_adr_o[25]
port 21 nsew signal output
rlabel metal2 s 60646 69200 60702 70000 6 caravel_wb_adr_o[26]
port 22 nsew signal output
rlabel metal2 s 62670 69200 62726 70000 6 caravel_wb_adr_o[27]
port 23 nsew signal output
rlabel metal2 s 9862 69200 9918 70000 6 caravel_wb_adr_o[2]
port 24 nsew signal output
rlabel metal2 s 12622 69200 12678 70000 6 caravel_wb_adr_o[3]
port 25 nsew signal output
rlabel metal2 s 15382 69200 15438 70000 6 caravel_wb_adr_o[4]
port 26 nsew signal output
rlabel metal2 s 17406 69200 17462 70000 6 caravel_wb_adr_o[5]
port 27 nsew signal output
rlabel metal2 s 19430 69200 19486 70000 6 caravel_wb_adr_o[6]
port 28 nsew signal output
rlabel metal2 s 21546 69200 21602 70000 6 caravel_wb_adr_o[7]
port 29 nsew signal output
rlabel metal2 s 23570 69200 23626 70000 6 caravel_wb_adr_o[8]
port 30 nsew signal output
rlabel metal2 s 25686 69200 25742 70000 6 caravel_wb_adr_o[9]
port 31 nsew signal output
rlabel metal2 s 938 69200 994 70000 6 caravel_wb_cyc_o
port 32 nsew signal output
rlabel metal2 s 5078 69200 5134 70000 6 caravel_wb_data_i[0]
port 33 nsew signal input
rlabel metal2 s 28354 69200 28410 70000 6 caravel_wb_data_i[10]
port 34 nsew signal input
rlabel metal2 s 30470 69200 30526 70000 6 caravel_wb_data_i[11]
port 35 nsew signal input
rlabel metal2 s 32494 69200 32550 70000 6 caravel_wb_data_i[12]
port 36 nsew signal input
rlabel metal2 s 34610 69200 34666 70000 6 caravel_wb_data_i[13]
port 37 nsew signal input
rlabel metal2 s 36634 69200 36690 70000 6 caravel_wb_data_i[14]
port 38 nsew signal input
rlabel metal2 s 38658 69200 38714 70000 6 caravel_wb_data_i[15]
port 39 nsew signal input
rlabel metal2 s 40774 69200 40830 70000 6 caravel_wb_data_i[16]
port 40 nsew signal input
rlabel metal2 s 42798 69200 42854 70000 6 caravel_wb_data_i[17]
port 41 nsew signal input
rlabel metal2 s 44822 69200 44878 70000 6 caravel_wb_data_i[18]
port 42 nsew signal input
rlabel metal2 s 46938 69200 46994 70000 6 caravel_wb_data_i[19]
port 43 nsew signal input
rlabel metal2 s 7838 69200 7894 70000 6 caravel_wb_data_i[1]
port 44 nsew signal input
rlabel metal2 s 48962 69200 49018 70000 6 caravel_wb_data_i[20]
port 45 nsew signal input
rlabel metal2 s 51078 69200 51134 70000 6 caravel_wb_data_i[21]
port 46 nsew signal input
rlabel metal2 s 53102 69200 53158 70000 6 caravel_wb_data_i[22]
port 47 nsew signal input
rlabel metal2 s 55126 69200 55182 70000 6 caravel_wb_data_i[23]
port 48 nsew signal input
rlabel metal2 s 57242 69200 57298 70000 6 caravel_wb_data_i[24]
port 49 nsew signal input
rlabel metal2 s 59266 69200 59322 70000 6 caravel_wb_data_i[25]
port 50 nsew signal input
rlabel metal2 s 61382 69200 61438 70000 6 caravel_wb_data_i[26]
port 51 nsew signal input
rlabel metal2 s 63406 69200 63462 70000 6 caravel_wb_data_i[27]
port 52 nsew signal input
rlabel metal2 s 64786 69200 64842 70000 6 caravel_wb_data_i[28]
port 53 nsew signal input
rlabel metal2 s 66166 69200 66222 70000 6 caravel_wb_data_i[29]
port 54 nsew signal input
rlabel metal2 s 10506 69200 10562 70000 6 caravel_wb_data_i[2]
port 55 nsew signal input
rlabel metal2 s 67546 69200 67602 70000 6 caravel_wb_data_i[30]
port 56 nsew signal input
rlabel metal2 s 68926 69200 68982 70000 6 caravel_wb_data_i[31]
port 57 nsew signal input
rlabel metal2 s 13266 69200 13322 70000 6 caravel_wb_data_i[3]
port 58 nsew signal input
rlabel metal2 s 16026 69200 16082 70000 6 caravel_wb_data_i[4]
port 59 nsew signal input
rlabel metal2 s 18050 69200 18106 70000 6 caravel_wb_data_i[5]
port 60 nsew signal input
rlabel metal2 s 20166 69200 20222 70000 6 caravel_wb_data_i[6]
port 61 nsew signal input
rlabel metal2 s 22190 69200 22246 70000 6 caravel_wb_data_i[7]
port 62 nsew signal input
rlabel metal2 s 24306 69200 24362 70000 6 caravel_wb_data_i[8]
port 63 nsew signal input
rlabel metal2 s 26330 69200 26386 70000 6 caravel_wb_data_i[9]
port 64 nsew signal input
rlabel metal2 s 5722 69200 5778 70000 6 caravel_wb_data_o[0]
port 65 nsew signal output
rlabel metal2 s 29090 69200 29146 70000 6 caravel_wb_data_o[10]
port 66 nsew signal output
rlabel metal2 s 31114 69200 31170 70000 6 caravel_wb_data_o[11]
port 67 nsew signal output
rlabel metal2 s 33230 69200 33286 70000 6 caravel_wb_data_o[12]
port 68 nsew signal output
rlabel metal2 s 35254 69200 35310 70000 6 caravel_wb_data_o[13]
port 69 nsew signal output
rlabel metal2 s 37278 69200 37334 70000 6 caravel_wb_data_o[14]
port 70 nsew signal output
rlabel metal2 s 39394 69200 39450 70000 6 caravel_wb_data_o[15]
port 71 nsew signal output
rlabel metal2 s 41418 69200 41474 70000 6 caravel_wb_data_o[16]
port 72 nsew signal output
rlabel metal2 s 43534 69200 43590 70000 6 caravel_wb_data_o[17]
port 73 nsew signal output
rlabel metal2 s 45558 69200 45614 70000 6 caravel_wb_data_o[18]
port 74 nsew signal output
rlabel metal2 s 47582 69200 47638 70000 6 caravel_wb_data_o[19]
port 75 nsew signal output
rlabel metal2 s 8482 69200 8538 70000 6 caravel_wb_data_o[1]
port 76 nsew signal output
rlabel metal2 s 49698 69200 49754 70000 6 caravel_wb_data_o[20]
port 77 nsew signal output
rlabel metal2 s 51722 69200 51778 70000 6 caravel_wb_data_o[21]
port 78 nsew signal output
rlabel metal2 s 53746 69200 53802 70000 6 caravel_wb_data_o[22]
port 79 nsew signal output
rlabel metal2 s 55862 69200 55918 70000 6 caravel_wb_data_o[23]
port 80 nsew signal output
rlabel metal2 s 57886 69200 57942 70000 6 caravel_wb_data_o[24]
port 81 nsew signal output
rlabel metal2 s 60002 69200 60058 70000 6 caravel_wb_data_o[25]
port 82 nsew signal output
rlabel metal2 s 62026 69200 62082 70000 6 caravel_wb_data_o[26]
port 83 nsew signal output
rlabel metal2 s 64050 69200 64106 70000 6 caravel_wb_data_o[27]
port 84 nsew signal output
rlabel metal2 s 65430 69200 65486 70000 6 caravel_wb_data_o[28]
port 85 nsew signal output
rlabel metal2 s 66810 69200 66866 70000 6 caravel_wb_data_o[29]
port 86 nsew signal output
rlabel metal2 s 11242 69200 11298 70000 6 caravel_wb_data_o[2]
port 87 nsew signal output
rlabel metal2 s 68190 69200 68246 70000 6 caravel_wb_data_o[30]
port 88 nsew signal output
rlabel metal2 s 69570 69200 69626 70000 6 caravel_wb_data_o[31]
port 89 nsew signal output
rlabel metal2 s 14002 69200 14058 70000 6 caravel_wb_data_o[3]
port 90 nsew signal output
rlabel metal2 s 16762 69200 16818 70000 6 caravel_wb_data_o[4]
port 91 nsew signal output
rlabel metal2 s 18786 69200 18842 70000 6 caravel_wb_data_o[5]
port 92 nsew signal output
rlabel metal2 s 20810 69200 20866 70000 6 caravel_wb_data_o[6]
port 93 nsew signal output
rlabel metal2 s 22926 69200 22982 70000 6 caravel_wb_data_o[7]
port 94 nsew signal output
rlabel metal2 s 24950 69200 25006 70000 6 caravel_wb_data_o[8]
port 95 nsew signal output
rlabel metal2 s 26974 69200 27030 70000 6 caravel_wb_data_o[9]
port 96 nsew signal output
rlabel metal2 s 1582 69200 1638 70000 6 caravel_wb_error_i
port 97 nsew signal input
rlabel metal2 s 6458 69200 6514 70000 6 caravel_wb_sel_o[0]
port 98 nsew signal output
rlabel metal2 s 9126 69200 9182 70000 6 caravel_wb_sel_o[1]
port 99 nsew signal output
rlabel metal2 s 11886 69200 11942 70000 6 caravel_wb_sel_o[2]
port 100 nsew signal output
rlabel metal2 s 14646 69200 14702 70000 6 caravel_wb_sel_o[3]
port 101 nsew signal output
rlabel metal2 s 2318 69200 2374 70000 6 caravel_wb_stall_i
port 102 nsew signal input
rlabel metal2 s 2962 69200 3018 70000 6 caravel_wb_stb_o
port 103 nsew signal output
rlabel metal2 s 3698 69200 3754 70000 6 caravel_wb_we_o
port 104 nsew signal output
rlabel metal3 s 0 688 800 808 6 core0Index[0]
port 105 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 core0Index[1]
port 106 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 core0Index[2]
port 107 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 core0Index[3]
port 108 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 core0Index[4]
port 109 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 core0Index[5]
port 110 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 core0Index[6]
port 111 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 core0Index[7]
port 112 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 core1Index[0]
port 113 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 core1Index[1]
port 114 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 core1Index[2]
port 115 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 core1Index[3]
port 116 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 core1Index[4]
port 117 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 core1Index[5]
port 118 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 core1Index[6]
port 119 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 core1Index[7]
port 120 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 manufacturerID[0]
port 121 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 manufacturerID[10]
port 122 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 manufacturerID[1]
port 123 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 manufacturerID[2]
port 124 nsew signal output
rlabel metal3 s 0 28976 800 29096 6 manufacturerID[3]
port 125 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 manufacturerID[4]
port 126 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 manufacturerID[5]
port 127 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 manufacturerID[6]
port 128 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 manufacturerID[7]
port 129 nsew signal output
rlabel metal3 s 0 36320 800 36440 6 manufacturerID[8]
port 130 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 manufacturerID[9]
port 131 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 partID[0]
port 132 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 partID[10]
port 133 nsew signal output
rlabel metal3 s 0 57264 800 57384 6 partID[11]
port 134 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 partID[12]
port 135 nsew signal output
rlabel metal3 s 0 60256 800 60376 6 partID[13]
port 136 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 partID[14]
port 137 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 partID[15]
port 138 nsew signal output
rlabel metal3 s 0 42304 800 42424 6 partID[1]
port 139 nsew signal output
rlabel metal3 s 0 43800 800 43920 6 partID[2]
port 140 nsew signal output
rlabel metal3 s 0 45296 800 45416 6 partID[3]
port 141 nsew signal output
rlabel metal3 s 0 46792 800 46912 6 partID[4]
port 142 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 partID[5]
port 143 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 partID[6]
port 144 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 partID[7]
port 145 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 partID[8]
port 146 nsew signal output
rlabel metal3 s 0 54272 800 54392 6 partID[9]
port 147 nsew signal output
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 148 nsew power input
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 148 nsew power input
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 148 nsew power input
rlabel metal3 s 0 64744 800 64864 6 versionID[0]
port 149 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 versionID[1]
port 150 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 versionID[2]
port 151 nsew signal output
rlabel metal3 s 0 69232 800 69352 6 versionID[3]
port 152 nsew signal output
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 153 nsew ground input
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 153 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 154 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_rst_i
port 155 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_ack_o
port 156 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[0]
port 157 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[10]
port 158 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[11]
port 159 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[12]
port 160 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_adr_i[13]
port 161 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[14]
port 162 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_adr_i[15]
port 163 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_adr_i[16]
port 164 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_adr_i[17]
port 165 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[18]
port 166 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_adr_i[19]
port 167 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[1]
port 168 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[20]
port 169 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 wbs_adr_i[21]
port 170 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[22]
port 171 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_adr_i[23]
port 172 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_adr_i[24]
port 173 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 wbs_adr_i[25]
port 174 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 wbs_adr_i[26]
port 175 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 wbs_adr_i[27]
port 176 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 wbs_adr_i[28]
port 177 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 wbs_adr_i[29]
port 178 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_adr_i[2]
port 179 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 wbs_adr_i[30]
port 180 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 wbs_adr_i[31]
port 181 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_adr_i[3]
port 182 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[4]
port 183 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[5]
port 184 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[6]
port 185 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_adr_i[7]
port 186 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[8]
port 187 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[9]
port 188 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_cyc_i
port 189 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_data_i[0]
port 190 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_data_i[10]
port 191 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_data_i[11]
port 192 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_data_i[12]
port 193 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_data_i[13]
port 194 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_data_i[14]
port 195 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_data_i[15]
port 196 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 wbs_data_i[16]
port 197 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 wbs_data_i[17]
port 198 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_data_i[18]
port 199 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 wbs_data_i[19]
port 200 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_data_i[1]
port 201 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_data_i[20]
port 202 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_data_i[21]
port 203 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_data_i[22]
port 204 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_data_i[23]
port 205 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_data_i[24]
port 206 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 wbs_data_i[25]
port 207 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wbs_data_i[26]
port 208 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 wbs_data_i[27]
port 209 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_data_i[28]
port 210 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 wbs_data_i[29]
port 211 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_data_i[2]
port 212 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 wbs_data_i[30]
port 213 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 wbs_data_i[31]
port 214 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_data_i[3]
port 215 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_data_i[4]
port 216 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_data_i[5]
port 217 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_data_i[6]
port 218 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_data_i[7]
port 219 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_data_i[8]
port 220 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_data_i[9]
port 221 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_data_o[0]
port 222 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_data_o[10]
port 223 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 wbs_data_o[11]
port 224 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_data_o[12]
port 225 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 wbs_data_o[13]
port 226 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 wbs_data_o[14]
port 227 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_data_o[15]
port 228 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 wbs_data_o[16]
port 229 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 wbs_data_o[17]
port 230 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 wbs_data_o[18]
port 231 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 wbs_data_o[19]
port 232 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 wbs_data_o[1]
port 233 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 wbs_data_o[20]
port 234 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 wbs_data_o[21]
port 235 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_data_o[22]
port 236 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 wbs_data_o[23]
port 237 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 wbs_data_o[24]
port 238 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 wbs_data_o[25]
port 239 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 wbs_data_o[26]
port 240 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 wbs_data_o[27]
port 241 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 wbs_data_o[28]
port 242 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 wbs_data_o[29]
port 243 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_data_o[2]
port 244 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 wbs_data_o[30]
port 245 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 wbs_data_o[31]
port 246 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_data_o[3]
port 247 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_data_o[4]
port 248 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wbs_data_o[5]
port 249 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_data_o[6]
port 250 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_data_o[7]
port 251 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_data_o[8]
port 252 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 wbs_data_o[9]
port 253 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_sel_i[0]
port 254 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_sel_i[1]
port 255 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_sel_i[2]
port 256 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_sel_i[3]
port 257 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_stb_i
port 258 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_we_i
port 259 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12327164
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/CaravelHost/runs/CaravelHost/results/finishing/CaravelHost.magic.gds
string GDS_START 841728
<< end >>

