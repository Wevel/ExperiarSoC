VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SPI
  CLASS BLOCK ;
  FOREIGN SPI ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 196.000 50.050 200.000 ;
    END
  END clk
  PIN peripheralBus_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END peripheralBus_address[0]
  PIN peripheralBus_address[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END peripheralBus_address[10]
  PIN peripheralBus_address[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END peripheralBus_address[11]
  PIN peripheralBus_address[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END peripheralBus_address[12]
  PIN peripheralBus_address[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END peripheralBus_address[13]
  PIN peripheralBus_address[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END peripheralBus_address[14]
  PIN peripheralBus_address[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END peripheralBus_address[15]
  PIN peripheralBus_address[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END peripheralBus_address[16]
  PIN peripheralBus_address[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END peripheralBus_address[17]
  PIN peripheralBus_address[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END peripheralBus_address[18]
  PIN peripheralBus_address[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END peripheralBus_address[19]
  PIN peripheralBus_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END peripheralBus_address[1]
  PIN peripheralBus_address[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END peripheralBus_address[20]
  PIN peripheralBus_address[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END peripheralBus_address[21]
  PIN peripheralBus_address[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END peripheralBus_address[22]
  PIN peripheralBus_address[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END peripheralBus_address[23]
  PIN peripheralBus_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END peripheralBus_address[2]
  PIN peripheralBus_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END peripheralBus_address[3]
  PIN peripheralBus_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END peripheralBus_address[4]
  PIN peripheralBus_address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END peripheralBus_address[5]
  PIN peripheralBus_address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END peripheralBus_address[6]
  PIN peripheralBus_address[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END peripheralBus_address[7]
  PIN peripheralBus_address[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END peripheralBus_address[8]
  PIN peripheralBus_address[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END peripheralBus_address[9]
  PIN peripheralBus_busy
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END peripheralBus_busy
  PIN peripheralBus_data[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END peripheralBus_data[0]
  PIN peripheralBus_data[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END peripheralBus_data[10]
  PIN peripheralBus_data[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END peripheralBus_data[11]
  PIN peripheralBus_data[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END peripheralBus_data[12]
  PIN peripheralBus_data[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END peripheralBus_data[13]
  PIN peripheralBus_data[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END peripheralBus_data[14]
  PIN peripheralBus_data[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END peripheralBus_data[15]
  PIN peripheralBus_data[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END peripheralBus_data[16]
  PIN peripheralBus_data[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END peripheralBus_data[17]
  PIN peripheralBus_data[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END peripheralBus_data[18]
  PIN peripheralBus_data[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END peripheralBus_data[19]
  PIN peripheralBus_data[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END peripheralBus_data[1]
  PIN peripheralBus_data[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END peripheralBus_data[20]
  PIN peripheralBus_data[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END peripheralBus_data[21]
  PIN peripheralBus_data[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END peripheralBus_data[22]
  PIN peripheralBus_data[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END peripheralBus_data[23]
  PIN peripheralBus_data[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END peripheralBus_data[24]
  PIN peripheralBus_data[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END peripheralBus_data[25]
  PIN peripheralBus_data[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END peripheralBus_data[26]
  PIN peripheralBus_data[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END peripheralBus_data[27]
  PIN peripheralBus_data[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END peripheralBus_data[28]
  PIN peripheralBus_data[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END peripheralBus_data[29]
  PIN peripheralBus_data[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END peripheralBus_data[2]
  PIN peripheralBus_data[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END peripheralBus_data[30]
  PIN peripheralBus_data[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END peripheralBus_data[31]
  PIN peripheralBus_data[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END peripheralBus_data[3]
  PIN peripheralBus_data[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END peripheralBus_data[4]
  PIN peripheralBus_data[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END peripheralBus_data[5]
  PIN peripheralBus_data[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END peripheralBus_data[6]
  PIN peripheralBus_data[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END peripheralBus_data[7]
  PIN peripheralBus_data[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END peripheralBus_data[8]
  PIN peripheralBus_data[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END peripheralBus_data[9]
  PIN peripheralBus_oe
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END peripheralBus_oe
  PIN peripheralBus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END peripheralBus_we
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 196.000 149.870 200.000 ;
    END
  END rst
  PIN spi_clk[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 9.560 200.000 10.160 ;
    END
  END spi_clk[0]
  PIN spi_clk[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 109.520 200.000 110.120 ;
    END
  END spi_clk[1]
  PIN spi_cs[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 29.280 200.000 29.880 ;
    END
  END spi_cs[0]
  PIN spi_cs[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 129.240 200.000 129.840 ;
    END
  END spi_cs[1]
  PIN spi_en[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 49.000 200.000 49.600 ;
    END
  END spi_en[0]
  PIN spi_en[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 148.960 200.000 149.560 ;
    END
  END spi_en[1]
  PIN spi_miso[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 69.400 200.000 70.000 ;
    END
  END spi_miso[0]
  PIN spi_miso[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 169.360 200.000 169.960 ;
    END
  END spi_miso[1]
  PIN spi_mosi[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 89.120 200.000 89.720 ;
    END
  END spi_mosi[0]
  PIN spi_mosi[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 189.080 200.000 189.680 ;
    END
  END spi_mosi[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 5.520 10.640 194.120 187.920 ;
      LAYER met2 ;
        RECT 6.990 195.720 49.490 198.405 ;
        RECT 50.330 195.720 149.310 198.405 ;
        RECT 150.150 195.720 190.810 198.405 ;
        RECT 6.990 1.515 190.810 195.720 ;
      LAYER met3 ;
        RECT 4.400 197.520 196.000 198.385 ;
        RECT 4.000 195.520 196.000 197.520 ;
        RECT 4.400 194.120 196.000 195.520 ;
        RECT 4.000 192.120 196.000 194.120 ;
        RECT 4.400 190.720 196.000 192.120 ;
        RECT 4.000 190.080 196.000 190.720 ;
        RECT 4.000 188.720 195.600 190.080 ;
        RECT 4.400 188.680 195.600 188.720 ;
        RECT 4.400 187.320 196.000 188.680 ;
        RECT 4.000 185.320 196.000 187.320 ;
        RECT 4.400 183.920 196.000 185.320 ;
        RECT 4.000 181.920 196.000 183.920 ;
        RECT 4.400 180.520 196.000 181.920 ;
        RECT 4.000 178.520 196.000 180.520 ;
        RECT 4.400 177.120 196.000 178.520 ;
        RECT 4.000 175.120 196.000 177.120 ;
        RECT 4.400 173.720 196.000 175.120 ;
        RECT 4.000 171.720 196.000 173.720 ;
        RECT 4.400 170.360 196.000 171.720 ;
        RECT 4.400 170.320 195.600 170.360 ;
        RECT 4.000 168.960 195.600 170.320 ;
        RECT 4.000 168.320 196.000 168.960 ;
        RECT 4.400 166.920 196.000 168.320 ;
        RECT 4.000 164.920 196.000 166.920 ;
        RECT 4.400 163.520 196.000 164.920 ;
        RECT 4.000 161.520 196.000 163.520 ;
        RECT 4.400 160.120 196.000 161.520 ;
        RECT 4.000 158.120 196.000 160.120 ;
        RECT 4.400 156.720 196.000 158.120 ;
        RECT 4.000 154.720 196.000 156.720 ;
        RECT 4.400 153.320 196.000 154.720 ;
        RECT 4.000 151.320 196.000 153.320 ;
        RECT 4.400 149.960 196.000 151.320 ;
        RECT 4.400 149.920 195.600 149.960 ;
        RECT 4.000 148.560 195.600 149.920 ;
        RECT 4.000 147.920 196.000 148.560 ;
        RECT 4.400 146.520 196.000 147.920 ;
        RECT 4.000 144.520 196.000 146.520 ;
        RECT 4.400 143.120 196.000 144.520 ;
        RECT 4.000 141.120 196.000 143.120 ;
        RECT 4.400 139.720 196.000 141.120 ;
        RECT 4.000 137.720 196.000 139.720 ;
        RECT 4.400 136.320 196.000 137.720 ;
        RECT 4.000 134.320 196.000 136.320 ;
        RECT 4.400 132.920 196.000 134.320 ;
        RECT 4.000 130.920 196.000 132.920 ;
        RECT 4.400 130.240 196.000 130.920 ;
        RECT 4.400 129.520 195.600 130.240 ;
        RECT 4.000 128.840 195.600 129.520 ;
        RECT 4.000 127.520 196.000 128.840 ;
        RECT 4.400 126.120 196.000 127.520 ;
        RECT 4.000 124.120 196.000 126.120 ;
        RECT 4.400 122.720 196.000 124.120 ;
        RECT 4.000 120.720 196.000 122.720 ;
        RECT 4.400 119.320 196.000 120.720 ;
        RECT 4.000 117.320 196.000 119.320 ;
        RECT 4.400 115.920 196.000 117.320 ;
        RECT 4.000 113.920 196.000 115.920 ;
        RECT 4.400 112.520 196.000 113.920 ;
        RECT 4.000 110.520 196.000 112.520 ;
        RECT 4.400 109.120 195.600 110.520 ;
        RECT 4.000 107.120 196.000 109.120 ;
        RECT 4.400 105.720 196.000 107.120 ;
        RECT 4.000 103.720 196.000 105.720 ;
        RECT 4.400 102.320 196.000 103.720 ;
        RECT 4.000 100.320 196.000 102.320 ;
        RECT 4.400 98.920 196.000 100.320 ;
        RECT 4.000 96.920 196.000 98.920 ;
        RECT 4.400 95.520 196.000 96.920 ;
        RECT 4.000 93.520 196.000 95.520 ;
        RECT 4.400 92.120 196.000 93.520 ;
        RECT 4.000 90.120 196.000 92.120 ;
        RECT 4.400 88.720 195.600 90.120 ;
        RECT 4.000 86.720 196.000 88.720 ;
        RECT 4.400 85.320 196.000 86.720 ;
        RECT 4.000 83.320 196.000 85.320 ;
        RECT 4.400 81.920 196.000 83.320 ;
        RECT 4.000 79.920 196.000 81.920 ;
        RECT 4.400 78.520 196.000 79.920 ;
        RECT 4.000 76.520 196.000 78.520 ;
        RECT 4.400 75.120 196.000 76.520 ;
        RECT 4.000 73.120 196.000 75.120 ;
        RECT 4.400 71.720 196.000 73.120 ;
        RECT 4.000 70.400 196.000 71.720 ;
        RECT 4.000 69.720 195.600 70.400 ;
        RECT 4.400 69.000 195.600 69.720 ;
        RECT 4.400 68.320 196.000 69.000 ;
        RECT 4.000 66.320 196.000 68.320 ;
        RECT 4.400 64.920 196.000 66.320 ;
        RECT 4.000 62.920 196.000 64.920 ;
        RECT 4.400 61.520 196.000 62.920 ;
        RECT 4.000 59.520 196.000 61.520 ;
        RECT 4.400 58.120 196.000 59.520 ;
        RECT 4.000 56.120 196.000 58.120 ;
        RECT 4.400 54.720 196.000 56.120 ;
        RECT 4.000 52.720 196.000 54.720 ;
        RECT 4.400 51.320 196.000 52.720 ;
        RECT 4.000 50.000 196.000 51.320 ;
        RECT 4.000 49.320 195.600 50.000 ;
        RECT 4.400 48.600 195.600 49.320 ;
        RECT 4.400 47.920 196.000 48.600 ;
        RECT 4.000 45.920 196.000 47.920 ;
        RECT 4.400 44.520 196.000 45.920 ;
        RECT 4.000 42.520 196.000 44.520 ;
        RECT 4.400 41.120 196.000 42.520 ;
        RECT 4.000 39.120 196.000 41.120 ;
        RECT 4.400 37.720 196.000 39.120 ;
        RECT 4.000 35.720 196.000 37.720 ;
        RECT 4.400 34.320 196.000 35.720 ;
        RECT 4.000 32.320 196.000 34.320 ;
        RECT 4.400 30.920 196.000 32.320 ;
        RECT 4.000 30.280 196.000 30.920 ;
        RECT 4.000 28.920 195.600 30.280 ;
        RECT 4.400 28.880 195.600 28.920 ;
        RECT 4.400 27.520 196.000 28.880 ;
        RECT 4.000 25.520 196.000 27.520 ;
        RECT 4.400 24.120 196.000 25.520 ;
        RECT 4.000 22.120 196.000 24.120 ;
        RECT 4.400 20.720 196.000 22.120 ;
        RECT 4.000 18.720 196.000 20.720 ;
        RECT 4.400 17.320 196.000 18.720 ;
        RECT 4.000 15.320 196.000 17.320 ;
        RECT 4.400 13.920 196.000 15.320 ;
        RECT 4.000 11.920 196.000 13.920 ;
        RECT 4.400 10.560 196.000 11.920 ;
        RECT 4.400 10.520 195.600 10.560 ;
        RECT 4.000 9.160 195.600 10.520 ;
        RECT 4.000 8.520 196.000 9.160 ;
        RECT 4.400 7.120 196.000 8.520 ;
        RECT 4.000 5.120 196.000 7.120 ;
        RECT 4.400 3.720 196.000 5.120 ;
        RECT 4.000 2.400 196.000 3.720 ;
        RECT 4.400 1.535 196.000 2.400 ;
  END
END SPI
END LIBRARY

