magic
tech sky130A
magscale 1 2
timestamp 1651278043
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 290 212 39638 37584
<< metal2 >>
rect 19982 39200 20038 40000
rect 294 0 350 800
rect 938 0 994 800
rect 1582 0 1638 800
rect 2318 0 2374 800
rect 2962 0 3018 800
rect 3606 0 3662 800
rect 4342 0 4398 800
rect 4986 0 5042 800
rect 5630 0 5686 800
rect 6366 0 6422 800
rect 7010 0 7066 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9770 0 9826 800
rect 10414 0 10470 800
rect 11058 0 11114 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 13174 0 13230 800
rect 13818 0 13874 800
rect 14462 0 14518 800
rect 15198 0 15254 800
rect 15842 0 15898 800
rect 16486 0 16542 800
rect 17222 0 17278 800
rect 17866 0 17922 800
rect 18602 0 18658 800
rect 19246 0 19302 800
rect 19890 0 19946 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22650 0 22706 800
rect 23294 0 23350 800
rect 24030 0 24086 800
rect 24674 0 24730 800
rect 25318 0 25374 800
rect 26054 0 26110 800
rect 26698 0 26754 800
rect 27342 0 27398 800
rect 28078 0 28134 800
rect 28722 0 28778 800
rect 29458 0 29514 800
rect 30102 0 30158 800
rect 30746 0 30802 800
rect 31482 0 31538 800
rect 32126 0 32182 800
rect 32770 0 32826 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34886 0 34942 800
rect 35530 0 35586 800
rect 36174 0 36230 800
rect 36910 0 36966 800
rect 37554 0 37610 800
rect 38198 0 38254 800
rect 38934 0 38990 800
rect 39578 0 39634 800
<< obsm2 >>
rect 296 39144 19926 39681
rect 20094 39144 39632 39681
rect 296 856 39632 39144
rect 406 167 882 856
rect 1050 167 1526 856
rect 1694 167 2262 856
rect 2430 167 2906 856
rect 3074 167 3550 856
rect 3718 167 4286 856
rect 4454 167 4930 856
rect 5098 167 5574 856
rect 5742 167 6310 856
rect 6478 167 6954 856
rect 7122 167 7690 856
rect 7858 167 8334 856
rect 8502 167 8978 856
rect 9146 167 9714 856
rect 9882 167 10358 856
rect 10526 167 11002 856
rect 11170 167 11738 856
rect 11906 167 12382 856
rect 12550 167 13118 856
rect 13286 167 13762 856
rect 13930 167 14406 856
rect 14574 167 15142 856
rect 15310 167 15786 856
rect 15954 167 16430 856
rect 16598 167 17166 856
rect 17334 167 17810 856
rect 17978 167 18546 856
rect 18714 167 19190 856
rect 19358 167 19834 856
rect 20002 167 20570 856
rect 20738 167 21214 856
rect 21382 167 21858 856
rect 22026 167 22594 856
rect 22762 167 23238 856
rect 23406 167 23974 856
rect 24142 167 24618 856
rect 24786 167 25262 856
rect 25430 167 25998 856
rect 26166 167 26642 856
rect 26810 167 27286 856
rect 27454 167 28022 856
rect 28190 167 28666 856
rect 28834 167 29402 856
rect 29570 167 30046 856
rect 30214 167 30690 856
rect 30858 167 31426 856
rect 31594 167 32070 856
rect 32238 167 32714 856
rect 32882 167 33450 856
rect 33618 167 34094 856
rect 34262 167 34830 856
rect 34998 167 35474 856
rect 35642 167 36118 856
rect 36286 167 36854 856
rect 37022 167 37498 856
rect 37666 167 38142 856
rect 38310 167 38878 856
rect 39046 167 39522 856
<< metal3 >>
rect 0 39584 800 39704
rect 39200 39448 40000 39568
rect 0 39176 800 39296
rect 0 38768 800 38888
rect 39200 38768 40000 38888
rect 0 38360 800 38480
rect 39200 38088 40000 38208
rect 0 37816 800 37936
rect 0 37408 800 37528
rect 39200 37408 40000 37528
rect 0 37000 800 37120
rect 0 36592 800 36712
rect 39200 36728 40000 36848
rect 0 36048 800 36168
rect 39200 36048 40000 36168
rect 0 35640 800 35760
rect 0 35232 800 35352
rect 39200 35232 40000 35352
rect 0 34824 800 34944
rect 0 34416 800 34536
rect 39200 34552 40000 34672
rect 0 33872 800 33992
rect 39200 33872 40000 33992
rect 0 33464 800 33584
rect 0 33056 800 33176
rect 39200 33192 40000 33312
rect 0 32648 800 32768
rect 39200 32512 40000 32632
rect 0 32104 800 32224
rect 0 31696 800 31816
rect 39200 31832 40000 31952
rect 0 31288 800 31408
rect 0 30880 800 31000
rect 39200 31016 40000 31136
rect 0 30336 800 30456
rect 39200 30336 40000 30456
rect 0 29928 800 30048
rect 0 29520 800 29640
rect 39200 29656 40000 29776
rect 0 29112 800 29232
rect 39200 28976 40000 29096
rect 0 28704 800 28824
rect 0 28160 800 28280
rect 39200 28296 40000 28416
rect 0 27752 800 27872
rect 39200 27616 40000 27736
rect 0 27344 800 27464
rect 0 26936 800 27056
rect 39200 26936 40000 27056
rect 0 26392 800 26512
rect 0 25984 800 26104
rect 39200 26120 40000 26240
rect 0 25576 800 25696
rect 39200 25440 40000 25560
rect 0 25168 800 25288
rect 0 24624 800 24744
rect 39200 24760 40000 24880
rect 0 24216 800 24336
rect 39200 24080 40000 24200
rect 0 23808 800 23928
rect 0 23400 800 23520
rect 39200 23400 40000 23520
rect 0 22992 800 23112
rect 39200 22720 40000 22840
rect 0 22448 800 22568
rect 0 22040 800 22160
rect 39200 21904 40000 22024
rect 0 21632 800 21752
rect 0 21224 800 21344
rect 39200 21224 40000 21344
rect 0 20680 800 20800
rect 39200 20544 40000 20664
rect 0 20272 800 20392
rect 0 19864 800 19984
rect 39200 19864 40000 19984
rect 0 19456 800 19576
rect 39200 19184 40000 19304
rect 0 18912 800 19032
rect 0 18504 800 18624
rect 39200 18504 40000 18624
rect 0 18096 800 18216
rect 0 17688 800 17808
rect 39200 17688 40000 17808
rect 0 17280 800 17400
rect 39200 17008 40000 17128
rect 0 16736 800 16856
rect 0 16328 800 16448
rect 39200 16328 40000 16448
rect 0 15920 800 16040
rect 0 15512 800 15632
rect 39200 15648 40000 15768
rect 0 14968 800 15088
rect 39200 14968 40000 15088
rect 0 14560 800 14680
rect 0 14152 800 14272
rect 39200 14288 40000 14408
rect 0 13744 800 13864
rect 39200 13608 40000 13728
rect 0 13200 800 13320
rect 0 12792 800 12912
rect 39200 12792 40000 12912
rect 0 12384 800 12504
rect 0 11976 800 12096
rect 39200 12112 40000 12232
rect 0 11568 800 11688
rect 39200 11432 40000 11552
rect 0 11024 800 11144
rect 0 10616 800 10736
rect 39200 10752 40000 10872
rect 0 10208 800 10328
rect 39200 10072 40000 10192
rect 0 9800 800 9920
rect 0 9256 800 9376
rect 39200 9392 40000 9512
rect 0 8848 800 8968
rect 0 8440 800 8560
rect 39200 8576 40000 8696
rect 0 8032 800 8152
rect 39200 7896 40000 8016
rect 0 7488 800 7608
rect 0 7080 800 7200
rect 39200 7216 40000 7336
rect 0 6672 800 6792
rect 39200 6536 40000 6656
rect 0 6264 800 6384
rect 0 5856 800 5976
rect 39200 5856 40000 5976
rect 0 5312 800 5432
rect 39200 5176 40000 5296
rect 0 4904 800 5024
rect 0 4496 800 4616
rect 39200 4360 40000 4480
rect 0 4088 800 4208
rect 0 3544 800 3664
rect 39200 3680 40000 3800
rect 0 3136 800 3256
rect 39200 3000 40000 3120
rect 0 2728 800 2848
rect 0 2320 800 2440
rect 39200 2320 40000 2440
rect 0 1776 800 1896
rect 39200 1640 40000 1760
rect 0 1368 800 1488
rect 0 960 800 1080
rect 39200 960 40000 1080
rect 0 552 800 672
rect 0 144 800 264
rect 39200 280 40000 400
<< obsm3 >>
rect 880 39648 39200 39677
rect 880 39504 39120 39648
rect 800 39376 39120 39504
rect 880 39368 39120 39376
rect 880 39096 39200 39368
rect 800 38968 39200 39096
rect 880 38688 39120 38968
rect 800 38560 39200 38688
rect 880 38288 39200 38560
rect 880 38280 39120 38288
rect 800 38016 39120 38280
rect 880 38008 39120 38016
rect 880 37736 39200 38008
rect 800 37608 39200 37736
rect 880 37328 39120 37608
rect 800 37200 39200 37328
rect 880 36928 39200 37200
rect 880 36920 39120 36928
rect 800 36792 39120 36920
rect 880 36648 39120 36792
rect 880 36512 39200 36648
rect 800 36248 39200 36512
rect 880 35968 39120 36248
rect 800 35840 39200 35968
rect 880 35560 39200 35840
rect 800 35432 39200 35560
rect 880 35152 39120 35432
rect 800 35024 39200 35152
rect 880 34752 39200 35024
rect 880 34744 39120 34752
rect 800 34616 39120 34744
rect 880 34472 39120 34616
rect 880 34336 39200 34472
rect 800 34072 39200 34336
rect 880 33792 39120 34072
rect 800 33664 39200 33792
rect 880 33392 39200 33664
rect 880 33384 39120 33392
rect 800 33256 39120 33384
rect 880 33112 39120 33256
rect 880 32976 39200 33112
rect 800 32848 39200 32976
rect 880 32712 39200 32848
rect 880 32568 39120 32712
rect 800 32432 39120 32568
rect 800 32304 39200 32432
rect 880 32032 39200 32304
rect 880 32024 39120 32032
rect 800 31896 39120 32024
rect 880 31752 39120 31896
rect 880 31616 39200 31752
rect 800 31488 39200 31616
rect 880 31216 39200 31488
rect 880 31208 39120 31216
rect 800 31080 39120 31208
rect 880 30936 39120 31080
rect 880 30800 39200 30936
rect 800 30536 39200 30800
rect 880 30256 39120 30536
rect 800 30128 39200 30256
rect 880 29856 39200 30128
rect 880 29848 39120 29856
rect 800 29720 39120 29848
rect 880 29576 39120 29720
rect 880 29440 39200 29576
rect 800 29312 39200 29440
rect 880 29176 39200 29312
rect 880 29032 39120 29176
rect 800 28904 39120 29032
rect 880 28896 39120 28904
rect 880 28624 39200 28896
rect 800 28496 39200 28624
rect 800 28360 39120 28496
rect 880 28216 39120 28360
rect 880 28080 39200 28216
rect 800 27952 39200 28080
rect 880 27816 39200 27952
rect 880 27672 39120 27816
rect 800 27544 39120 27672
rect 880 27536 39120 27544
rect 880 27264 39200 27536
rect 800 27136 39200 27264
rect 880 26856 39120 27136
rect 800 26592 39200 26856
rect 880 26320 39200 26592
rect 880 26312 39120 26320
rect 800 26184 39120 26312
rect 880 26040 39120 26184
rect 880 25904 39200 26040
rect 800 25776 39200 25904
rect 880 25640 39200 25776
rect 880 25496 39120 25640
rect 800 25368 39120 25496
rect 880 25360 39120 25368
rect 880 25088 39200 25360
rect 800 24960 39200 25088
rect 800 24824 39120 24960
rect 880 24680 39120 24824
rect 880 24544 39200 24680
rect 800 24416 39200 24544
rect 880 24280 39200 24416
rect 880 24136 39120 24280
rect 800 24008 39120 24136
rect 880 24000 39120 24008
rect 880 23728 39200 24000
rect 800 23600 39200 23728
rect 880 23320 39120 23600
rect 800 23192 39200 23320
rect 880 22920 39200 23192
rect 880 22912 39120 22920
rect 800 22648 39120 22912
rect 880 22640 39120 22648
rect 880 22368 39200 22640
rect 800 22240 39200 22368
rect 880 22104 39200 22240
rect 880 21960 39120 22104
rect 800 21832 39120 21960
rect 880 21824 39120 21832
rect 880 21552 39200 21824
rect 800 21424 39200 21552
rect 880 21144 39120 21424
rect 800 20880 39200 21144
rect 880 20744 39200 20880
rect 880 20600 39120 20744
rect 800 20472 39120 20600
rect 880 20464 39120 20472
rect 880 20192 39200 20464
rect 800 20064 39200 20192
rect 880 19784 39120 20064
rect 800 19656 39200 19784
rect 880 19384 39200 19656
rect 880 19376 39120 19384
rect 800 19112 39120 19376
rect 880 19104 39120 19112
rect 880 18832 39200 19104
rect 800 18704 39200 18832
rect 880 18424 39120 18704
rect 800 18296 39200 18424
rect 880 18016 39200 18296
rect 800 17888 39200 18016
rect 880 17608 39120 17888
rect 800 17480 39200 17608
rect 880 17208 39200 17480
rect 880 17200 39120 17208
rect 800 16936 39120 17200
rect 880 16928 39120 16936
rect 880 16656 39200 16928
rect 800 16528 39200 16656
rect 880 16248 39120 16528
rect 800 16120 39200 16248
rect 880 15848 39200 16120
rect 880 15840 39120 15848
rect 800 15712 39120 15840
rect 880 15568 39120 15712
rect 880 15432 39200 15568
rect 800 15168 39200 15432
rect 880 14888 39120 15168
rect 800 14760 39200 14888
rect 880 14488 39200 14760
rect 880 14480 39120 14488
rect 800 14352 39120 14480
rect 880 14208 39120 14352
rect 880 14072 39200 14208
rect 800 13944 39200 14072
rect 880 13808 39200 13944
rect 880 13664 39120 13808
rect 800 13528 39120 13664
rect 800 13400 39200 13528
rect 880 13120 39200 13400
rect 800 12992 39200 13120
rect 880 12712 39120 12992
rect 800 12584 39200 12712
rect 880 12312 39200 12584
rect 880 12304 39120 12312
rect 800 12176 39120 12304
rect 880 12032 39120 12176
rect 880 11896 39200 12032
rect 800 11768 39200 11896
rect 880 11632 39200 11768
rect 880 11488 39120 11632
rect 800 11352 39120 11488
rect 800 11224 39200 11352
rect 880 10952 39200 11224
rect 880 10944 39120 10952
rect 800 10816 39120 10944
rect 880 10672 39120 10816
rect 880 10536 39200 10672
rect 800 10408 39200 10536
rect 880 10272 39200 10408
rect 880 10128 39120 10272
rect 800 10000 39120 10128
rect 880 9992 39120 10000
rect 880 9720 39200 9992
rect 800 9592 39200 9720
rect 800 9456 39120 9592
rect 880 9312 39120 9456
rect 880 9176 39200 9312
rect 800 9048 39200 9176
rect 880 8776 39200 9048
rect 880 8768 39120 8776
rect 800 8640 39120 8768
rect 880 8496 39120 8640
rect 880 8360 39200 8496
rect 800 8232 39200 8360
rect 880 8096 39200 8232
rect 880 7952 39120 8096
rect 800 7816 39120 7952
rect 800 7688 39200 7816
rect 880 7416 39200 7688
rect 880 7408 39120 7416
rect 800 7280 39120 7408
rect 880 7136 39120 7280
rect 880 7000 39200 7136
rect 800 6872 39200 7000
rect 880 6736 39200 6872
rect 880 6592 39120 6736
rect 800 6464 39120 6592
rect 880 6456 39120 6464
rect 880 6184 39200 6456
rect 800 6056 39200 6184
rect 880 5776 39120 6056
rect 800 5512 39200 5776
rect 880 5376 39200 5512
rect 880 5232 39120 5376
rect 800 5104 39120 5232
rect 880 5096 39120 5104
rect 880 4824 39200 5096
rect 800 4696 39200 4824
rect 880 4560 39200 4696
rect 880 4416 39120 4560
rect 800 4288 39120 4416
rect 880 4280 39120 4288
rect 880 4008 39200 4280
rect 800 3880 39200 4008
rect 800 3744 39120 3880
rect 880 3600 39120 3744
rect 880 3464 39200 3600
rect 800 3336 39200 3464
rect 880 3200 39200 3336
rect 880 3056 39120 3200
rect 800 2928 39120 3056
rect 880 2920 39120 2928
rect 880 2648 39200 2920
rect 800 2520 39200 2648
rect 880 2240 39120 2520
rect 800 1976 39200 2240
rect 880 1840 39200 1976
rect 880 1696 39120 1840
rect 800 1568 39120 1696
rect 880 1560 39120 1568
rect 880 1288 39200 1560
rect 800 1160 39200 1288
rect 880 880 39120 1160
rect 800 752 39200 880
rect 880 480 39200 752
rect 880 472 39120 480
rect 800 344 39120 472
rect 880 200 39120 344
rect 880 171 39200 200
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal2 s 38934 0 38990 800 6 clk
port 1 nsew signal input
rlabel metal3 s 39200 280 40000 400 6 gpio0_input[0]
port 2 nsew signal input
rlabel metal3 s 39200 21224 40000 21344 6 gpio0_input[10]
port 3 nsew signal input
rlabel metal3 s 39200 23400 40000 23520 6 gpio0_input[11]
port 4 nsew signal input
rlabel metal3 s 39200 25440 40000 25560 6 gpio0_input[12]
port 5 nsew signal input
rlabel metal3 s 39200 27616 40000 27736 6 gpio0_input[13]
port 6 nsew signal input
rlabel metal3 s 39200 29656 40000 29776 6 gpio0_input[14]
port 7 nsew signal input
rlabel metal3 s 39200 31832 40000 31952 6 gpio0_input[15]
port 8 nsew signal input
rlabel metal3 s 39200 33872 40000 33992 6 gpio0_input[16]
port 9 nsew signal input
rlabel metal3 s 39200 36048 40000 36168 6 gpio0_input[17]
port 10 nsew signal input
rlabel metal3 s 39200 38088 40000 38208 6 gpio0_input[18]
port 11 nsew signal input
rlabel metal3 s 39200 2320 40000 2440 6 gpio0_input[1]
port 12 nsew signal input
rlabel metal3 s 39200 4360 40000 4480 6 gpio0_input[2]
port 13 nsew signal input
rlabel metal3 s 39200 6536 40000 6656 6 gpio0_input[3]
port 14 nsew signal input
rlabel metal3 s 39200 8576 40000 8696 6 gpio0_input[4]
port 15 nsew signal input
rlabel metal3 s 39200 10752 40000 10872 6 gpio0_input[5]
port 16 nsew signal input
rlabel metal3 s 39200 12792 40000 12912 6 gpio0_input[6]
port 17 nsew signal input
rlabel metal3 s 39200 14968 40000 15088 6 gpio0_input[7]
port 18 nsew signal input
rlabel metal3 s 39200 17008 40000 17128 6 gpio0_input[8]
port 19 nsew signal input
rlabel metal3 s 39200 19184 40000 19304 6 gpio0_input[9]
port 20 nsew signal input
rlabel metal3 s 39200 960 40000 1080 6 gpio0_oe[0]
port 21 nsew signal output
rlabel metal3 s 39200 21904 40000 22024 6 gpio0_oe[10]
port 22 nsew signal output
rlabel metal3 s 39200 24080 40000 24200 6 gpio0_oe[11]
port 23 nsew signal output
rlabel metal3 s 39200 26120 40000 26240 6 gpio0_oe[12]
port 24 nsew signal output
rlabel metal3 s 39200 28296 40000 28416 6 gpio0_oe[13]
port 25 nsew signal output
rlabel metal3 s 39200 30336 40000 30456 6 gpio0_oe[14]
port 26 nsew signal output
rlabel metal3 s 39200 32512 40000 32632 6 gpio0_oe[15]
port 27 nsew signal output
rlabel metal3 s 39200 34552 40000 34672 6 gpio0_oe[16]
port 28 nsew signal output
rlabel metal3 s 39200 36728 40000 36848 6 gpio0_oe[17]
port 29 nsew signal output
rlabel metal3 s 39200 38768 40000 38888 6 gpio0_oe[18]
port 30 nsew signal output
rlabel metal3 s 39200 3000 40000 3120 6 gpio0_oe[1]
port 31 nsew signal output
rlabel metal3 s 39200 5176 40000 5296 6 gpio0_oe[2]
port 32 nsew signal output
rlabel metal3 s 39200 7216 40000 7336 6 gpio0_oe[3]
port 33 nsew signal output
rlabel metal3 s 39200 9392 40000 9512 6 gpio0_oe[4]
port 34 nsew signal output
rlabel metal3 s 39200 11432 40000 11552 6 gpio0_oe[5]
port 35 nsew signal output
rlabel metal3 s 39200 13608 40000 13728 6 gpio0_oe[6]
port 36 nsew signal output
rlabel metal3 s 39200 15648 40000 15768 6 gpio0_oe[7]
port 37 nsew signal output
rlabel metal3 s 39200 17688 40000 17808 6 gpio0_oe[8]
port 38 nsew signal output
rlabel metal3 s 39200 19864 40000 19984 6 gpio0_oe[9]
port 39 nsew signal output
rlabel metal3 s 39200 1640 40000 1760 6 gpio0_output[0]
port 40 nsew signal output
rlabel metal3 s 39200 22720 40000 22840 6 gpio0_output[10]
port 41 nsew signal output
rlabel metal3 s 39200 24760 40000 24880 6 gpio0_output[11]
port 42 nsew signal output
rlabel metal3 s 39200 26936 40000 27056 6 gpio0_output[12]
port 43 nsew signal output
rlabel metal3 s 39200 28976 40000 29096 6 gpio0_output[13]
port 44 nsew signal output
rlabel metal3 s 39200 31016 40000 31136 6 gpio0_output[14]
port 45 nsew signal output
rlabel metal3 s 39200 33192 40000 33312 6 gpio0_output[15]
port 46 nsew signal output
rlabel metal3 s 39200 35232 40000 35352 6 gpio0_output[16]
port 47 nsew signal output
rlabel metal3 s 39200 37408 40000 37528 6 gpio0_output[17]
port 48 nsew signal output
rlabel metal3 s 39200 39448 40000 39568 6 gpio0_output[18]
port 49 nsew signal output
rlabel metal3 s 39200 3680 40000 3800 6 gpio0_output[1]
port 50 nsew signal output
rlabel metal3 s 39200 5856 40000 5976 6 gpio0_output[2]
port 51 nsew signal output
rlabel metal3 s 39200 7896 40000 8016 6 gpio0_output[3]
port 52 nsew signal output
rlabel metal3 s 39200 10072 40000 10192 6 gpio0_output[4]
port 53 nsew signal output
rlabel metal3 s 39200 12112 40000 12232 6 gpio0_output[5]
port 54 nsew signal output
rlabel metal3 s 39200 14288 40000 14408 6 gpio0_output[6]
port 55 nsew signal output
rlabel metal3 s 39200 16328 40000 16448 6 gpio0_output[7]
port 56 nsew signal output
rlabel metal3 s 39200 18504 40000 18624 6 gpio0_output[8]
port 57 nsew signal output
rlabel metal3 s 39200 20544 40000 20664 6 gpio0_output[9]
port 58 nsew signal output
rlabel metal2 s 294 0 350 800 6 gpio1_input[0]
port 59 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 gpio1_input[10]
port 60 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 gpio1_input[11]
port 61 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 gpio1_input[12]
port 62 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 gpio1_input[13]
port 63 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 gpio1_input[14]
port 64 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 gpio1_input[15]
port 65 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 gpio1_input[16]
port 66 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 gpio1_input[17]
port 67 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 gpio1_input[18]
port 68 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 gpio1_input[1]
port 69 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 gpio1_input[2]
port 70 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 gpio1_input[3]
port 71 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 gpio1_input[4]
port 72 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 gpio1_input[5]
port 73 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 gpio1_input[6]
port 74 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 gpio1_input[7]
port 75 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 gpio1_input[8]
port 76 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 gpio1_input[9]
port 77 nsew signal input
rlabel metal2 s 938 0 994 800 6 gpio1_oe[0]
port 78 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 gpio1_oe[10]
port 79 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 gpio1_oe[11]
port 80 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 gpio1_oe[12]
port 81 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 gpio1_oe[13]
port 82 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 gpio1_oe[14]
port 83 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 gpio1_oe[15]
port 84 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 gpio1_oe[16]
port 85 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 gpio1_oe[17]
port 86 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 gpio1_oe[18]
port 87 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 gpio1_oe[1]
port 88 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 gpio1_oe[2]
port 89 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 gpio1_oe[3]
port 90 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 gpio1_oe[4]
port 91 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 gpio1_oe[5]
port 92 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 gpio1_oe[6]
port 93 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 gpio1_oe[7]
port 94 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 gpio1_oe[8]
port 95 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 gpio1_oe[9]
port 96 nsew signal output
rlabel metal2 s 1582 0 1638 800 6 gpio1_output[0]
port 97 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 gpio1_output[10]
port 98 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 gpio1_output[11]
port 99 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 gpio1_output[12]
port 100 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 gpio1_output[13]
port 101 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 gpio1_output[14]
port 102 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 gpio1_output[15]
port 103 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 gpio1_output[16]
port 104 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 gpio1_output[17]
port 105 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 gpio1_output[18]
port 106 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 gpio1_output[1]
port 107 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 gpio1_output[2]
port 108 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 gpio1_output[3]
port 109 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 gpio1_output[4]
port 110 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 gpio1_output[5]
port 111 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 gpio1_output[6]
port 112 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 gpio1_output[7]
port 113 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 gpio1_output[8]
port 114 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 gpio1_output[9]
port 115 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 peripheralBus_address[0]
port 116 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 peripheralBus_address[10]
port 117 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 peripheralBus_address[11]
port 118 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 peripheralBus_address[12]
port 119 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 peripheralBus_address[13]
port 120 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 peripheralBus_address[14]
port 121 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 peripheralBus_address[15]
port 122 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 peripheralBus_address[16]
port 123 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 peripheralBus_address[17]
port 124 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 peripheralBus_address[18]
port 125 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 peripheralBus_address[19]
port 126 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 peripheralBus_address[1]
port 127 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 peripheralBus_address[20]
port 128 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 peripheralBus_address[21]
port 129 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 peripheralBus_address[22]
port 130 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 peripheralBus_address[23]
port 131 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 peripheralBus_address[2]
port 132 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 peripheralBus_address[3]
port 133 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 peripheralBus_address[4]
port 134 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 peripheralBus_address[5]
port 135 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 peripheralBus_address[6]
port 136 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 peripheralBus_address[7]
port 137 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 peripheralBus_address[8]
port 138 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 peripheralBus_address[9]
port 139 nsew signal input
rlabel metal3 s 0 144 800 264 6 peripheralBus_busy
port 140 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 peripheralBus_dataIn[0]
port 141 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 peripheralBus_dataIn[10]
port 142 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 peripheralBus_dataIn[11]
port 143 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 peripheralBus_dataIn[12]
port 144 nsew signal input
rlabel metal3 s 0 18912 800 19032 6 peripheralBus_dataIn[13]
port 145 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 peripheralBus_dataIn[14]
port 146 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 peripheralBus_dataIn[15]
port 147 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 peripheralBus_dataIn[16]
port 148 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 peripheralBus_dataIn[17]
port 149 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 peripheralBus_dataIn[18]
port 150 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 peripheralBus_dataIn[19]
port 151 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 peripheralBus_dataIn[1]
port 152 nsew signal input
rlabel metal3 s 0 28160 800 28280 6 peripheralBus_dataIn[20]
port 153 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 peripheralBus_dataIn[21]
port 154 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 peripheralBus_dataIn[22]
port 155 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 peripheralBus_dataIn[23]
port 156 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 peripheralBus_dataIn[24]
port 157 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 peripheralBus_dataIn[25]
port 158 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 peripheralBus_dataIn[26]
port 159 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 peripheralBus_dataIn[27]
port 160 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 peripheralBus_dataIn[28]
port 161 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 peripheralBus_dataIn[29]
port 162 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 peripheralBus_dataIn[2]
port 163 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 peripheralBus_dataIn[30]
port 164 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 peripheralBus_dataIn[31]
port 165 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 peripheralBus_dataIn[3]
port 166 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 peripheralBus_dataIn[4]
port 167 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 peripheralBus_dataIn[5]
port 168 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 peripheralBus_dataIn[6]
port 169 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 peripheralBus_dataIn[7]
port 170 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 peripheralBus_dataIn[8]
port 171 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 peripheralBus_dataIn[9]
port 172 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 peripheralBus_dataOut[0]
port 173 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 peripheralBus_dataOut[10]
port 174 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 peripheralBus_dataOut[11]
port 175 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 peripheralBus_dataOut[12]
port 176 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 peripheralBus_dataOut[13]
port 177 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 peripheralBus_dataOut[14]
port 178 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 peripheralBus_dataOut[15]
port 179 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 peripheralBus_dataOut[16]
port 180 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 peripheralBus_dataOut[17]
port 181 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 peripheralBus_dataOut[18]
port 182 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 peripheralBus_dataOut[19]
port 183 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 peripheralBus_dataOut[1]
port 184 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 peripheralBus_dataOut[20]
port 185 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 peripheralBus_dataOut[21]
port 186 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 peripheralBus_dataOut[22]
port 187 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 peripheralBus_dataOut[23]
port 188 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 peripheralBus_dataOut[24]
port 189 nsew signal output
rlabel metal3 s 0 34416 800 34536 6 peripheralBus_dataOut[25]
port 190 nsew signal output
rlabel metal3 s 0 35232 800 35352 6 peripheralBus_dataOut[26]
port 191 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 peripheralBus_dataOut[27]
port 192 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 peripheralBus_dataOut[28]
port 193 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 peripheralBus_dataOut[29]
port 194 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 peripheralBus_dataOut[2]
port 195 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 peripheralBus_dataOut[30]
port 196 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 peripheralBus_dataOut[31]
port 197 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 peripheralBus_dataOut[3]
port 198 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 peripheralBus_dataOut[4]
port 199 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 peripheralBus_dataOut[5]
port 200 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 peripheralBus_dataOut[6]
port 201 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 peripheralBus_dataOut[7]
port 202 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 peripheralBus_dataOut[8]
port 203 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 peripheralBus_dataOut[9]
port 204 nsew signal output
rlabel metal3 s 0 552 800 672 6 peripheralBus_oe
port 205 nsew signal input
rlabel metal3 s 0 960 800 1080 6 peripheralBus_we
port 206 nsew signal input
rlabel metal2 s 19982 39200 20038 40000 6 requestOutput
port 207 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 rst
port 208 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 209 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 209 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 210 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2552386
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripheral_GPIO/runs/Peripheral_GPIO/results/finishing/GPIO.magic.gds
string GDS_START 286020
<< end >>

