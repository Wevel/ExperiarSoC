magic
tech sky130A
magscale 1 2
timestamp 1652654706
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 474 1368 99990 97424
<< metal2 >>
rect 478 0 534 800
rect 1398 0 1454 800
rect 2410 0 2466 800
rect 3422 0 3478 800
rect 4434 0 4490 800
rect 5446 0 5502 800
rect 6458 0 6514 800
rect 7470 0 7526 800
rect 8390 0 8446 800
rect 9402 0 9458 800
rect 10414 0 10470 800
rect 11426 0 11482 800
rect 12438 0 12494 800
rect 13450 0 13506 800
rect 14462 0 14518 800
rect 15474 0 15530 800
rect 16394 0 16450 800
rect 17406 0 17462 800
rect 18418 0 18474 800
rect 19430 0 19486 800
rect 20442 0 20498 800
rect 21454 0 21510 800
rect 22466 0 22522 800
rect 23478 0 23534 800
rect 24398 0 24454 800
rect 25410 0 25466 800
rect 26422 0 26478 800
rect 27434 0 27490 800
rect 28446 0 28502 800
rect 29458 0 29514 800
rect 30470 0 30526 800
rect 31390 0 31446 800
rect 32402 0 32458 800
rect 33414 0 33470 800
rect 34426 0 34482 800
rect 35438 0 35494 800
rect 36450 0 36506 800
rect 37462 0 37518 800
rect 38474 0 38530 800
rect 39394 0 39450 800
rect 40406 0 40462 800
rect 41418 0 41474 800
rect 42430 0 42486 800
rect 43442 0 43498 800
rect 44454 0 44510 800
rect 45466 0 45522 800
rect 46478 0 46534 800
rect 47398 0 47454 800
rect 48410 0 48466 800
rect 49422 0 49478 800
rect 50434 0 50490 800
rect 51446 0 51502 800
rect 52458 0 52514 800
rect 53470 0 53526 800
rect 54390 0 54446 800
rect 55402 0 55458 800
rect 56414 0 56470 800
rect 57426 0 57482 800
rect 58438 0 58494 800
rect 59450 0 59506 800
rect 60462 0 60518 800
rect 61474 0 61530 800
rect 62394 0 62450 800
rect 63406 0 63462 800
rect 64418 0 64474 800
rect 65430 0 65486 800
rect 66442 0 66498 800
rect 67454 0 67510 800
rect 68466 0 68522 800
rect 69478 0 69534 800
rect 70398 0 70454 800
rect 71410 0 71466 800
rect 72422 0 72478 800
rect 73434 0 73490 800
rect 74446 0 74502 800
rect 75458 0 75514 800
rect 76470 0 76526 800
rect 77390 0 77446 800
rect 78402 0 78458 800
rect 79414 0 79470 800
rect 80426 0 80482 800
rect 81438 0 81494 800
rect 82450 0 82506 800
rect 83462 0 83518 800
rect 84474 0 84530 800
rect 85394 0 85450 800
rect 86406 0 86462 800
rect 87418 0 87474 800
rect 88430 0 88486 800
rect 89442 0 89498 800
rect 90454 0 90510 800
rect 91466 0 91522 800
rect 92478 0 92534 800
rect 93398 0 93454 800
rect 94410 0 94466 800
rect 95422 0 95478 800
rect 96434 0 96490 800
rect 97446 0 97502 800
rect 98458 0 98514 800
rect 99470 0 99526 800
<< obsm2 >>
rect 480 856 99986 99657
rect 590 167 1342 856
rect 1510 167 2354 856
rect 2522 167 3366 856
rect 3534 167 4378 856
rect 4546 167 5390 856
rect 5558 167 6402 856
rect 6570 167 7414 856
rect 7582 167 8334 856
rect 8502 167 9346 856
rect 9514 167 10358 856
rect 10526 167 11370 856
rect 11538 167 12382 856
rect 12550 167 13394 856
rect 13562 167 14406 856
rect 14574 167 15418 856
rect 15586 167 16338 856
rect 16506 167 17350 856
rect 17518 167 18362 856
rect 18530 167 19374 856
rect 19542 167 20386 856
rect 20554 167 21398 856
rect 21566 167 22410 856
rect 22578 167 23422 856
rect 23590 167 24342 856
rect 24510 167 25354 856
rect 25522 167 26366 856
rect 26534 167 27378 856
rect 27546 167 28390 856
rect 28558 167 29402 856
rect 29570 167 30414 856
rect 30582 167 31334 856
rect 31502 167 32346 856
rect 32514 167 33358 856
rect 33526 167 34370 856
rect 34538 167 35382 856
rect 35550 167 36394 856
rect 36562 167 37406 856
rect 37574 167 38418 856
rect 38586 167 39338 856
rect 39506 167 40350 856
rect 40518 167 41362 856
rect 41530 167 42374 856
rect 42542 167 43386 856
rect 43554 167 44398 856
rect 44566 167 45410 856
rect 45578 167 46422 856
rect 46590 167 47342 856
rect 47510 167 48354 856
rect 48522 167 49366 856
rect 49534 167 50378 856
rect 50546 167 51390 856
rect 51558 167 52402 856
rect 52570 167 53414 856
rect 53582 167 54334 856
rect 54502 167 55346 856
rect 55514 167 56358 856
rect 56526 167 57370 856
rect 57538 167 58382 856
rect 58550 167 59394 856
rect 59562 167 60406 856
rect 60574 167 61418 856
rect 61586 167 62338 856
rect 62506 167 63350 856
rect 63518 167 64362 856
rect 64530 167 65374 856
rect 65542 167 66386 856
rect 66554 167 67398 856
rect 67566 167 68410 856
rect 68578 167 69422 856
rect 69590 167 70342 856
rect 70510 167 71354 856
rect 71522 167 72366 856
rect 72534 167 73378 856
rect 73546 167 74390 856
rect 74558 167 75402 856
rect 75570 167 76414 856
rect 76582 167 77334 856
rect 77502 167 78346 856
rect 78514 167 79358 856
rect 79526 167 80370 856
rect 80538 167 81382 856
rect 81550 167 82394 856
rect 82562 167 83406 856
rect 83574 167 84418 856
rect 84586 167 85338 856
rect 85506 167 86350 856
rect 86518 167 87362 856
rect 87530 167 88374 856
rect 88542 167 89386 856
rect 89554 167 90398 856
rect 90566 167 91410 856
rect 91578 167 92422 856
rect 92590 167 93342 856
rect 93510 167 94354 856
rect 94522 167 95366 856
rect 95534 167 96378 856
rect 96546 167 97390 856
rect 97558 167 98402 856
rect 98570 167 99414 856
rect 99582 167 99986 856
<< metal3 >>
rect 99200 99560 100000 99680
rect 99200 99016 100000 99136
rect 99200 98472 100000 98592
rect 99200 98064 100000 98184
rect 99200 97520 100000 97640
rect 99200 96976 100000 97096
rect 99200 96432 100000 96552
rect 99200 96024 100000 96144
rect 99200 95480 100000 95600
rect 99200 94936 100000 95056
rect 99200 94392 100000 94512
rect 99200 93984 100000 94104
rect 99200 93440 100000 93560
rect 99200 92896 100000 93016
rect 99200 92488 100000 92608
rect 99200 91944 100000 92064
rect 99200 91400 100000 91520
rect 99200 90856 100000 90976
rect 99200 90448 100000 90568
rect 99200 89904 100000 90024
rect 99200 89360 100000 89480
rect 99200 88816 100000 88936
rect 99200 88408 100000 88528
rect 99200 87864 100000 87984
rect 99200 87320 100000 87440
rect 99200 86776 100000 86896
rect 99200 86368 100000 86488
rect 99200 85824 100000 85944
rect 99200 85280 100000 85400
rect 99200 84872 100000 84992
rect 99200 84328 100000 84448
rect 99200 83784 100000 83904
rect 99200 83240 100000 83360
rect 99200 82832 100000 82952
rect 99200 82288 100000 82408
rect 99200 81744 100000 81864
rect 99200 81200 100000 81320
rect 99200 80792 100000 80912
rect 99200 80248 100000 80368
rect 99200 79704 100000 79824
rect 99200 79296 100000 79416
rect 99200 78752 100000 78872
rect 99200 78208 100000 78328
rect 99200 77664 100000 77784
rect 99200 77256 100000 77376
rect 99200 76712 100000 76832
rect 99200 76168 100000 76288
rect 99200 75624 100000 75744
rect 99200 75216 100000 75336
rect 99200 74672 100000 74792
rect 99200 74128 100000 74248
rect 99200 73584 100000 73704
rect 99200 73176 100000 73296
rect 99200 72632 100000 72752
rect 99200 72088 100000 72208
rect 99200 71680 100000 71800
rect 99200 71136 100000 71256
rect 99200 70592 100000 70712
rect 99200 70048 100000 70168
rect 99200 69640 100000 69760
rect 99200 69096 100000 69216
rect 99200 68552 100000 68672
rect 99200 68008 100000 68128
rect 99200 67600 100000 67720
rect 99200 67056 100000 67176
rect 99200 66512 100000 66632
rect 99200 66104 100000 66224
rect 99200 65560 100000 65680
rect 99200 65016 100000 65136
rect 99200 64472 100000 64592
rect 99200 64064 100000 64184
rect 99200 63520 100000 63640
rect 99200 62976 100000 63096
rect 99200 62432 100000 62552
rect 99200 62024 100000 62144
rect 99200 61480 100000 61600
rect 99200 60936 100000 61056
rect 99200 60392 100000 60512
rect 99200 59984 100000 60104
rect 99200 59440 100000 59560
rect 99200 58896 100000 59016
rect 99200 58488 100000 58608
rect 99200 57944 100000 58064
rect 99200 57400 100000 57520
rect 99200 56856 100000 56976
rect 99200 56448 100000 56568
rect 99200 55904 100000 56024
rect 99200 55360 100000 55480
rect 99200 54816 100000 54936
rect 99200 54408 100000 54528
rect 99200 53864 100000 53984
rect 99200 53320 100000 53440
rect 99200 52912 100000 53032
rect 99200 52368 100000 52488
rect 99200 51824 100000 51944
rect 99200 51280 100000 51400
rect 99200 50872 100000 50992
rect 99200 50328 100000 50448
rect 99200 49784 100000 49904
rect 99200 49240 100000 49360
rect 99200 48832 100000 48952
rect 99200 48288 100000 48408
rect 99200 47744 100000 47864
rect 99200 47200 100000 47320
rect 99200 46792 100000 46912
rect 99200 46248 100000 46368
rect 99200 45704 100000 45824
rect 99200 45296 100000 45416
rect 99200 44752 100000 44872
rect 99200 44208 100000 44328
rect 99200 43664 100000 43784
rect 99200 43256 100000 43376
rect 99200 42712 100000 42832
rect 99200 42168 100000 42288
rect 99200 41624 100000 41744
rect 99200 41216 100000 41336
rect 99200 40672 100000 40792
rect 99200 40128 100000 40248
rect 99200 39720 100000 39840
rect 99200 39176 100000 39296
rect 99200 38632 100000 38752
rect 99200 38088 100000 38208
rect 99200 37680 100000 37800
rect 99200 37136 100000 37256
rect 99200 36592 100000 36712
rect 99200 36048 100000 36168
rect 99200 35640 100000 35760
rect 99200 35096 100000 35216
rect 99200 34552 100000 34672
rect 99200 34008 100000 34128
rect 99200 33600 100000 33720
rect 99200 33056 100000 33176
rect 99200 32512 100000 32632
rect 99200 32104 100000 32224
rect 99200 31560 100000 31680
rect 99200 31016 100000 31136
rect 99200 30472 100000 30592
rect 99200 30064 100000 30184
rect 99200 29520 100000 29640
rect 99200 28976 100000 29096
rect 99200 28432 100000 28552
rect 99200 28024 100000 28144
rect 99200 27480 100000 27600
rect 99200 26936 100000 27056
rect 99200 26528 100000 26648
rect 99200 25984 100000 26104
rect 99200 25440 100000 25560
rect 99200 24896 100000 25016
rect 99200 24488 100000 24608
rect 99200 23944 100000 24064
rect 99200 23400 100000 23520
rect 99200 22856 100000 22976
rect 99200 22448 100000 22568
rect 99200 21904 100000 22024
rect 99200 21360 100000 21480
rect 99200 20816 100000 20936
rect 99200 20408 100000 20528
rect 99200 19864 100000 19984
rect 99200 19320 100000 19440
rect 99200 18912 100000 19032
rect 99200 18368 100000 18488
rect 99200 17824 100000 17944
rect 99200 17280 100000 17400
rect 99200 16872 100000 16992
rect 99200 16328 100000 16448
rect 99200 15784 100000 15904
rect 99200 15240 100000 15360
rect 99200 14832 100000 14952
rect 99200 14288 100000 14408
rect 99200 13744 100000 13864
rect 99200 13336 100000 13456
rect 99200 12792 100000 12912
rect 99200 12248 100000 12368
rect 99200 11704 100000 11824
rect 99200 11296 100000 11416
rect 99200 10752 100000 10872
rect 99200 10208 100000 10328
rect 99200 9664 100000 9784
rect 99200 9256 100000 9376
rect 99200 8712 100000 8832
rect 99200 8168 100000 8288
rect 99200 7624 100000 7744
rect 99200 7216 100000 7336
rect 99200 6672 100000 6792
rect 99200 6128 100000 6248
rect 99200 5720 100000 5840
rect 99200 5176 100000 5296
rect 99200 4632 100000 4752
rect 99200 4088 100000 4208
rect 99200 3680 100000 3800
rect 99200 3136 100000 3256
rect 99200 2592 100000 2712
rect 99200 2048 100000 2168
rect 99200 1640 100000 1760
rect 99200 1096 100000 1216
rect 99200 552 100000 672
rect 99200 144 100000 264
<< obsm3 >>
rect 1853 99480 99120 99653
rect 1853 99216 99991 99480
rect 1853 98936 99120 99216
rect 1853 98672 99991 98936
rect 1853 98392 99120 98672
rect 1853 98264 99991 98392
rect 1853 97984 99120 98264
rect 1853 97720 99991 97984
rect 1853 97440 99120 97720
rect 1853 97176 99991 97440
rect 1853 96896 99120 97176
rect 1853 96632 99991 96896
rect 1853 96352 99120 96632
rect 1853 96224 99991 96352
rect 1853 95944 99120 96224
rect 1853 95680 99991 95944
rect 1853 95400 99120 95680
rect 1853 95136 99991 95400
rect 1853 94856 99120 95136
rect 1853 94592 99991 94856
rect 1853 94312 99120 94592
rect 1853 94184 99991 94312
rect 1853 93904 99120 94184
rect 1853 93640 99991 93904
rect 1853 93360 99120 93640
rect 1853 93096 99991 93360
rect 1853 92816 99120 93096
rect 1853 92688 99991 92816
rect 1853 92408 99120 92688
rect 1853 92144 99991 92408
rect 1853 91864 99120 92144
rect 1853 91600 99991 91864
rect 1853 91320 99120 91600
rect 1853 91056 99991 91320
rect 1853 90776 99120 91056
rect 1853 90648 99991 90776
rect 1853 90368 99120 90648
rect 1853 90104 99991 90368
rect 1853 89824 99120 90104
rect 1853 89560 99991 89824
rect 1853 89280 99120 89560
rect 1853 89016 99991 89280
rect 1853 88736 99120 89016
rect 1853 88608 99991 88736
rect 1853 88328 99120 88608
rect 1853 88064 99991 88328
rect 1853 87784 99120 88064
rect 1853 87520 99991 87784
rect 1853 87240 99120 87520
rect 1853 86976 99991 87240
rect 1853 86696 99120 86976
rect 1853 86568 99991 86696
rect 1853 86288 99120 86568
rect 1853 86024 99991 86288
rect 1853 85744 99120 86024
rect 1853 85480 99991 85744
rect 1853 85200 99120 85480
rect 1853 85072 99991 85200
rect 1853 84792 99120 85072
rect 1853 84528 99991 84792
rect 1853 84248 99120 84528
rect 1853 83984 99991 84248
rect 1853 83704 99120 83984
rect 1853 83440 99991 83704
rect 1853 83160 99120 83440
rect 1853 83032 99991 83160
rect 1853 82752 99120 83032
rect 1853 82488 99991 82752
rect 1853 82208 99120 82488
rect 1853 81944 99991 82208
rect 1853 81664 99120 81944
rect 1853 81400 99991 81664
rect 1853 81120 99120 81400
rect 1853 80992 99991 81120
rect 1853 80712 99120 80992
rect 1853 80448 99991 80712
rect 1853 80168 99120 80448
rect 1853 79904 99991 80168
rect 1853 79624 99120 79904
rect 1853 79496 99991 79624
rect 1853 79216 99120 79496
rect 1853 78952 99991 79216
rect 1853 78672 99120 78952
rect 1853 78408 99991 78672
rect 1853 78128 99120 78408
rect 1853 77864 99991 78128
rect 1853 77584 99120 77864
rect 1853 77456 99991 77584
rect 1853 77176 99120 77456
rect 1853 76912 99991 77176
rect 1853 76632 99120 76912
rect 1853 76368 99991 76632
rect 1853 76088 99120 76368
rect 1853 75824 99991 76088
rect 1853 75544 99120 75824
rect 1853 75416 99991 75544
rect 1853 75136 99120 75416
rect 1853 74872 99991 75136
rect 1853 74592 99120 74872
rect 1853 74328 99991 74592
rect 1853 74048 99120 74328
rect 1853 73784 99991 74048
rect 1853 73504 99120 73784
rect 1853 73376 99991 73504
rect 1853 73096 99120 73376
rect 1853 72832 99991 73096
rect 1853 72552 99120 72832
rect 1853 72288 99991 72552
rect 1853 72008 99120 72288
rect 1853 71880 99991 72008
rect 1853 71600 99120 71880
rect 1853 71336 99991 71600
rect 1853 71056 99120 71336
rect 1853 70792 99991 71056
rect 1853 70512 99120 70792
rect 1853 70248 99991 70512
rect 1853 69968 99120 70248
rect 1853 69840 99991 69968
rect 1853 69560 99120 69840
rect 1853 69296 99991 69560
rect 1853 69016 99120 69296
rect 1853 68752 99991 69016
rect 1853 68472 99120 68752
rect 1853 68208 99991 68472
rect 1853 67928 99120 68208
rect 1853 67800 99991 67928
rect 1853 67520 99120 67800
rect 1853 67256 99991 67520
rect 1853 66976 99120 67256
rect 1853 66712 99991 66976
rect 1853 66432 99120 66712
rect 1853 66304 99991 66432
rect 1853 66024 99120 66304
rect 1853 65760 99991 66024
rect 1853 65480 99120 65760
rect 1853 65216 99991 65480
rect 1853 64936 99120 65216
rect 1853 64672 99991 64936
rect 1853 64392 99120 64672
rect 1853 64264 99991 64392
rect 1853 63984 99120 64264
rect 1853 63720 99991 63984
rect 1853 63440 99120 63720
rect 1853 63176 99991 63440
rect 1853 62896 99120 63176
rect 1853 62632 99991 62896
rect 1853 62352 99120 62632
rect 1853 62224 99991 62352
rect 1853 61944 99120 62224
rect 1853 61680 99991 61944
rect 1853 61400 99120 61680
rect 1853 61136 99991 61400
rect 1853 60856 99120 61136
rect 1853 60592 99991 60856
rect 1853 60312 99120 60592
rect 1853 60184 99991 60312
rect 1853 59904 99120 60184
rect 1853 59640 99991 59904
rect 1853 59360 99120 59640
rect 1853 59096 99991 59360
rect 1853 58816 99120 59096
rect 1853 58688 99991 58816
rect 1853 58408 99120 58688
rect 1853 58144 99991 58408
rect 1853 57864 99120 58144
rect 1853 57600 99991 57864
rect 1853 57320 99120 57600
rect 1853 57056 99991 57320
rect 1853 56776 99120 57056
rect 1853 56648 99991 56776
rect 1853 56368 99120 56648
rect 1853 56104 99991 56368
rect 1853 55824 99120 56104
rect 1853 55560 99991 55824
rect 1853 55280 99120 55560
rect 1853 55016 99991 55280
rect 1853 54736 99120 55016
rect 1853 54608 99991 54736
rect 1853 54328 99120 54608
rect 1853 54064 99991 54328
rect 1853 53784 99120 54064
rect 1853 53520 99991 53784
rect 1853 53240 99120 53520
rect 1853 53112 99991 53240
rect 1853 52832 99120 53112
rect 1853 52568 99991 52832
rect 1853 52288 99120 52568
rect 1853 52024 99991 52288
rect 1853 51744 99120 52024
rect 1853 51480 99991 51744
rect 1853 51200 99120 51480
rect 1853 51072 99991 51200
rect 1853 50792 99120 51072
rect 1853 50528 99991 50792
rect 1853 50248 99120 50528
rect 1853 49984 99991 50248
rect 1853 49704 99120 49984
rect 1853 49440 99991 49704
rect 1853 49160 99120 49440
rect 1853 49032 99991 49160
rect 1853 48752 99120 49032
rect 1853 48488 99991 48752
rect 1853 48208 99120 48488
rect 1853 47944 99991 48208
rect 1853 47664 99120 47944
rect 1853 47400 99991 47664
rect 1853 47120 99120 47400
rect 1853 46992 99991 47120
rect 1853 46712 99120 46992
rect 1853 46448 99991 46712
rect 1853 46168 99120 46448
rect 1853 45904 99991 46168
rect 1853 45624 99120 45904
rect 1853 45496 99991 45624
rect 1853 45216 99120 45496
rect 1853 44952 99991 45216
rect 1853 44672 99120 44952
rect 1853 44408 99991 44672
rect 1853 44128 99120 44408
rect 1853 43864 99991 44128
rect 1853 43584 99120 43864
rect 1853 43456 99991 43584
rect 1853 43176 99120 43456
rect 1853 42912 99991 43176
rect 1853 42632 99120 42912
rect 1853 42368 99991 42632
rect 1853 42088 99120 42368
rect 1853 41824 99991 42088
rect 1853 41544 99120 41824
rect 1853 41416 99991 41544
rect 1853 41136 99120 41416
rect 1853 40872 99991 41136
rect 1853 40592 99120 40872
rect 1853 40328 99991 40592
rect 1853 40048 99120 40328
rect 1853 39920 99991 40048
rect 1853 39640 99120 39920
rect 1853 39376 99991 39640
rect 1853 39096 99120 39376
rect 1853 38832 99991 39096
rect 1853 38552 99120 38832
rect 1853 38288 99991 38552
rect 1853 38008 99120 38288
rect 1853 37880 99991 38008
rect 1853 37600 99120 37880
rect 1853 37336 99991 37600
rect 1853 37056 99120 37336
rect 1853 36792 99991 37056
rect 1853 36512 99120 36792
rect 1853 36248 99991 36512
rect 1853 35968 99120 36248
rect 1853 35840 99991 35968
rect 1853 35560 99120 35840
rect 1853 35296 99991 35560
rect 1853 35016 99120 35296
rect 1853 34752 99991 35016
rect 1853 34472 99120 34752
rect 1853 34208 99991 34472
rect 1853 33928 99120 34208
rect 1853 33800 99991 33928
rect 1853 33520 99120 33800
rect 1853 33256 99991 33520
rect 1853 32976 99120 33256
rect 1853 32712 99991 32976
rect 1853 32432 99120 32712
rect 1853 32304 99991 32432
rect 1853 32024 99120 32304
rect 1853 31760 99991 32024
rect 1853 31480 99120 31760
rect 1853 31216 99991 31480
rect 1853 30936 99120 31216
rect 1853 30672 99991 30936
rect 1853 30392 99120 30672
rect 1853 30264 99991 30392
rect 1853 29984 99120 30264
rect 1853 29720 99991 29984
rect 1853 29440 99120 29720
rect 1853 29176 99991 29440
rect 1853 28896 99120 29176
rect 1853 28632 99991 28896
rect 1853 28352 99120 28632
rect 1853 28224 99991 28352
rect 1853 27944 99120 28224
rect 1853 27680 99991 27944
rect 1853 27400 99120 27680
rect 1853 27136 99991 27400
rect 1853 26856 99120 27136
rect 1853 26728 99991 26856
rect 1853 26448 99120 26728
rect 1853 26184 99991 26448
rect 1853 25904 99120 26184
rect 1853 25640 99991 25904
rect 1853 25360 99120 25640
rect 1853 25096 99991 25360
rect 1853 24816 99120 25096
rect 1853 24688 99991 24816
rect 1853 24408 99120 24688
rect 1853 24144 99991 24408
rect 1853 23864 99120 24144
rect 1853 23600 99991 23864
rect 1853 23320 99120 23600
rect 1853 23056 99991 23320
rect 1853 22776 99120 23056
rect 1853 22648 99991 22776
rect 1853 22368 99120 22648
rect 1853 22104 99991 22368
rect 1853 21824 99120 22104
rect 1853 21560 99991 21824
rect 1853 21280 99120 21560
rect 1853 21016 99991 21280
rect 1853 20736 99120 21016
rect 1853 20608 99991 20736
rect 1853 20328 99120 20608
rect 1853 20064 99991 20328
rect 1853 19784 99120 20064
rect 1853 19520 99991 19784
rect 1853 19240 99120 19520
rect 1853 19112 99991 19240
rect 1853 18832 99120 19112
rect 1853 18568 99991 18832
rect 1853 18288 99120 18568
rect 1853 18024 99991 18288
rect 1853 17744 99120 18024
rect 1853 17480 99991 17744
rect 1853 17200 99120 17480
rect 1853 17072 99991 17200
rect 1853 16792 99120 17072
rect 1853 16528 99991 16792
rect 1853 16248 99120 16528
rect 1853 15984 99991 16248
rect 1853 15704 99120 15984
rect 1853 15440 99991 15704
rect 1853 15160 99120 15440
rect 1853 15032 99991 15160
rect 1853 14752 99120 15032
rect 1853 14488 99991 14752
rect 1853 14208 99120 14488
rect 1853 13944 99991 14208
rect 1853 13664 99120 13944
rect 1853 13536 99991 13664
rect 1853 13256 99120 13536
rect 1853 12992 99991 13256
rect 1853 12712 99120 12992
rect 1853 12448 99991 12712
rect 1853 12168 99120 12448
rect 1853 11904 99991 12168
rect 1853 11624 99120 11904
rect 1853 11496 99991 11624
rect 1853 11216 99120 11496
rect 1853 10952 99991 11216
rect 1853 10672 99120 10952
rect 1853 10408 99991 10672
rect 1853 10128 99120 10408
rect 1853 9864 99991 10128
rect 1853 9584 99120 9864
rect 1853 9456 99991 9584
rect 1853 9176 99120 9456
rect 1853 8912 99991 9176
rect 1853 8632 99120 8912
rect 1853 8368 99991 8632
rect 1853 8088 99120 8368
rect 1853 7824 99991 8088
rect 1853 7544 99120 7824
rect 1853 7416 99991 7544
rect 1853 7136 99120 7416
rect 1853 6872 99991 7136
rect 1853 6592 99120 6872
rect 1853 6328 99991 6592
rect 1853 6048 99120 6328
rect 1853 5920 99991 6048
rect 1853 5640 99120 5920
rect 1853 5376 99991 5640
rect 1853 5096 99120 5376
rect 1853 4832 99991 5096
rect 1853 4552 99120 4832
rect 1853 4288 99991 4552
rect 1853 4008 99120 4288
rect 1853 3880 99991 4008
rect 1853 3600 99120 3880
rect 1853 3336 99991 3600
rect 1853 3056 99120 3336
rect 1853 2792 99991 3056
rect 1853 2512 99120 2792
rect 1853 2248 99991 2512
rect 1853 1968 99120 2248
rect 1853 1840 99991 1968
rect 1853 1560 99120 1840
rect 1853 1296 99991 1560
rect 1853 1016 99120 1296
rect 1853 752 99991 1016
rect 1853 472 99120 752
rect 1853 344 99991 472
rect 1853 171 99120 344
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 90955 3571 96288 75853
rect 96768 3571 99117 75853
<< labels >>
rlabel metal3 s 99200 4088 100000 4208 6 sram0_csb0
port 1 nsew signal output
rlabel metal3 s 99200 4632 100000 4752 6 sram0_csb1
port 2 nsew signal output
rlabel metal3 s 99200 7624 100000 7744 6 sram0_dout0[0]
port 3 nsew signal input
rlabel metal3 s 99200 44208 100000 44328 6 sram0_dout0[10]
port 4 nsew signal input
rlabel metal3 s 99200 46792 100000 46912 6 sram0_dout0[11]
port 5 nsew signal input
rlabel metal3 s 99200 49240 100000 49360 6 sram0_dout0[12]
port 6 nsew signal input
rlabel metal3 s 99200 51824 100000 51944 6 sram0_dout0[13]
port 7 nsew signal input
rlabel metal3 s 99200 54408 100000 54528 6 sram0_dout0[14]
port 8 nsew signal input
rlabel metal3 s 99200 56856 100000 56976 6 sram0_dout0[15]
port 9 nsew signal input
rlabel metal3 s 99200 59440 100000 59560 6 sram0_dout0[16]
port 10 nsew signal input
rlabel metal3 s 99200 62024 100000 62144 6 sram0_dout0[17]
port 11 nsew signal input
rlabel metal3 s 99200 64472 100000 64592 6 sram0_dout0[18]
port 12 nsew signal input
rlabel metal3 s 99200 67056 100000 67176 6 sram0_dout0[19]
port 13 nsew signal input
rlabel metal3 s 99200 11704 100000 11824 6 sram0_dout0[1]
port 14 nsew signal input
rlabel metal3 s 99200 69640 100000 69760 6 sram0_dout0[20]
port 15 nsew signal input
rlabel metal3 s 99200 72088 100000 72208 6 sram0_dout0[21]
port 16 nsew signal input
rlabel metal3 s 99200 74672 100000 74792 6 sram0_dout0[22]
port 17 nsew signal input
rlabel metal3 s 99200 77256 100000 77376 6 sram0_dout0[23]
port 18 nsew signal input
rlabel metal3 s 99200 79704 100000 79824 6 sram0_dout0[24]
port 19 nsew signal input
rlabel metal3 s 99200 82288 100000 82408 6 sram0_dout0[25]
port 20 nsew signal input
rlabel metal3 s 99200 84872 100000 84992 6 sram0_dout0[26]
port 21 nsew signal input
rlabel metal3 s 99200 87320 100000 87440 6 sram0_dout0[27]
port 22 nsew signal input
rlabel metal3 s 99200 89904 100000 90024 6 sram0_dout0[28]
port 23 nsew signal input
rlabel metal3 s 99200 92488 100000 92608 6 sram0_dout0[29]
port 24 nsew signal input
rlabel metal3 s 99200 15784 100000 15904 6 sram0_dout0[2]
port 25 nsew signal input
rlabel metal3 s 99200 94936 100000 95056 6 sram0_dout0[30]
port 26 nsew signal input
rlabel metal3 s 99200 97520 100000 97640 6 sram0_dout0[31]
port 27 nsew signal input
rlabel metal3 s 99200 19864 100000 19984 6 sram0_dout0[3]
port 28 nsew signal input
rlabel metal3 s 99200 23944 100000 24064 6 sram0_dout0[4]
port 29 nsew signal input
rlabel metal3 s 99200 27480 100000 27600 6 sram0_dout0[5]
port 30 nsew signal input
rlabel metal3 s 99200 31016 100000 31136 6 sram0_dout0[6]
port 31 nsew signal input
rlabel metal3 s 99200 34552 100000 34672 6 sram0_dout0[7]
port 32 nsew signal input
rlabel metal3 s 99200 38088 100000 38208 6 sram0_dout0[8]
port 33 nsew signal input
rlabel metal3 s 99200 41624 100000 41744 6 sram0_dout0[9]
port 34 nsew signal input
rlabel metal3 s 99200 8168 100000 8288 6 sram0_dout1[0]
port 35 nsew signal input
rlabel metal3 s 99200 44752 100000 44872 6 sram0_dout1[10]
port 36 nsew signal input
rlabel metal3 s 99200 47200 100000 47320 6 sram0_dout1[11]
port 37 nsew signal input
rlabel metal3 s 99200 49784 100000 49904 6 sram0_dout1[12]
port 38 nsew signal input
rlabel metal3 s 99200 52368 100000 52488 6 sram0_dout1[13]
port 39 nsew signal input
rlabel metal3 s 99200 54816 100000 54936 6 sram0_dout1[14]
port 40 nsew signal input
rlabel metal3 s 99200 57400 100000 57520 6 sram0_dout1[15]
port 41 nsew signal input
rlabel metal3 s 99200 59984 100000 60104 6 sram0_dout1[16]
port 42 nsew signal input
rlabel metal3 s 99200 62432 100000 62552 6 sram0_dout1[17]
port 43 nsew signal input
rlabel metal3 s 99200 65016 100000 65136 6 sram0_dout1[18]
port 44 nsew signal input
rlabel metal3 s 99200 67600 100000 67720 6 sram0_dout1[19]
port 45 nsew signal input
rlabel metal3 s 99200 12248 100000 12368 6 sram0_dout1[1]
port 46 nsew signal input
rlabel metal3 s 99200 70048 100000 70168 6 sram0_dout1[20]
port 47 nsew signal input
rlabel metal3 s 99200 72632 100000 72752 6 sram0_dout1[21]
port 48 nsew signal input
rlabel metal3 s 99200 75216 100000 75336 6 sram0_dout1[22]
port 49 nsew signal input
rlabel metal3 s 99200 77664 100000 77784 6 sram0_dout1[23]
port 50 nsew signal input
rlabel metal3 s 99200 80248 100000 80368 6 sram0_dout1[24]
port 51 nsew signal input
rlabel metal3 s 99200 82832 100000 82952 6 sram0_dout1[25]
port 52 nsew signal input
rlabel metal3 s 99200 85280 100000 85400 6 sram0_dout1[26]
port 53 nsew signal input
rlabel metal3 s 99200 87864 100000 87984 6 sram0_dout1[27]
port 54 nsew signal input
rlabel metal3 s 99200 90448 100000 90568 6 sram0_dout1[28]
port 55 nsew signal input
rlabel metal3 s 99200 92896 100000 93016 6 sram0_dout1[29]
port 56 nsew signal input
rlabel metal3 s 99200 16328 100000 16448 6 sram0_dout1[2]
port 57 nsew signal input
rlabel metal3 s 99200 95480 100000 95600 6 sram0_dout1[30]
port 58 nsew signal input
rlabel metal3 s 99200 98064 100000 98184 6 sram0_dout1[31]
port 59 nsew signal input
rlabel metal3 s 99200 20408 100000 20528 6 sram0_dout1[3]
port 60 nsew signal input
rlabel metal3 s 99200 24488 100000 24608 6 sram0_dout1[4]
port 61 nsew signal input
rlabel metal3 s 99200 28024 100000 28144 6 sram0_dout1[5]
port 62 nsew signal input
rlabel metal3 s 99200 31560 100000 31680 6 sram0_dout1[6]
port 63 nsew signal input
rlabel metal3 s 99200 35096 100000 35216 6 sram0_dout1[7]
port 64 nsew signal input
rlabel metal3 s 99200 38632 100000 38752 6 sram0_dout1[8]
port 65 nsew signal input
rlabel metal3 s 99200 42168 100000 42288 6 sram0_dout1[9]
port 66 nsew signal input
rlabel metal3 s 99200 5176 100000 5296 6 sram1_csb0
port 67 nsew signal output
rlabel metal3 s 99200 5720 100000 5840 6 sram1_csb1
port 68 nsew signal output
rlabel metal3 s 99200 8712 100000 8832 6 sram1_dout0[0]
port 69 nsew signal input
rlabel metal3 s 99200 45296 100000 45416 6 sram1_dout0[10]
port 70 nsew signal input
rlabel metal3 s 99200 47744 100000 47864 6 sram1_dout0[11]
port 71 nsew signal input
rlabel metal3 s 99200 50328 100000 50448 6 sram1_dout0[12]
port 72 nsew signal input
rlabel metal3 s 99200 52912 100000 53032 6 sram1_dout0[13]
port 73 nsew signal input
rlabel metal3 s 99200 55360 100000 55480 6 sram1_dout0[14]
port 74 nsew signal input
rlabel metal3 s 99200 57944 100000 58064 6 sram1_dout0[15]
port 75 nsew signal input
rlabel metal3 s 99200 60392 100000 60512 6 sram1_dout0[16]
port 76 nsew signal input
rlabel metal3 s 99200 62976 100000 63096 6 sram1_dout0[17]
port 77 nsew signal input
rlabel metal3 s 99200 65560 100000 65680 6 sram1_dout0[18]
port 78 nsew signal input
rlabel metal3 s 99200 68008 100000 68128 6 sram1_dout0[19]
port 79 nsew signal input
rlabel metal3 s 99200 12792 100000 12912 6 sram1_dout0[1]
port 80 nsew signal input
rlabel metal3 s 99200 70592 100000 70712 6 sram1_dout0[20]
port 81 nsew signal input
rlabel metal3 s 99200 73176 100000 73296 6 sram1_dout0[21]
port 82 nsew signal input
rlabel metal3 s 99200 75624 100000 75744 6 sram1_dout0[22]
port 83 nsew signal input
rlabel metal3 s 99200 78208 100000 78328 6 sram1_dout0[23]
port 84 nsew signal input
rlabel metal3 s 99200 80792 100000 80912 6 sram1_dout0[24]
port 85 nsew signal input
rlabel metal3 s 99200 83240 100000 83360 6 sram1_dout0[25]
port 86 nsew signal input
rlabel metal3 s 99200 85824 100000 85944 6 sram1_dout0[26]
port 87 nsew signal input
rlabel metal3 s 99200 88408 100000 88528 6 sram1_dout0[27]
port 88 nsew signal input
rlabel metal3 s 99200 90856 100000 90976 6 sram1_dout0[28]
port 89 nsew signal input
rlabel metal3 s 99200 93440 100000 93560 6 sram1_dout0[29]
port 90 nsew signal input
rlabel metal3 s 99200 16872 100000 16992 6 sram1_dout0[2]
port 91 nsew signal input
rlabel metal3 s 99200 96024 100000 96144 6 sram1_dout0[30]
port 92 nsew signal input
rlabel metal3 s 99200 98472 100000 98592 6 sram1_dout0[31]
port 93 nsew signal input
rlabel metal3 s 99200 20816 100000 20936 6 sram1_dout0[3]
port 94 nsew signal input
rlabel metal3 s 99200 24896 100000 25016 6 sram1_dout0[4]
port 95 nsew signal input
rlabel metal3 s 99200 28432 100000 28552 6 sram1_dout0[5]
port 96 nsew signal input
rlabel metal3 s 99200 32104 100000 32224 6 sram1_dout0[6]
port 97 nsew signal input
rlabel metal3 s 99200 35640 100000 35760 6 sram1_dout0[7]
port 98 nsew signal input
rlabel metal3 s 99200 39176 100000 39296 6 sram1_dout0[8]
port 99 nsew signal input
rlabel metal3 s 99200 42712 100000 42832 6 sram1_dout0[9]
port 100 nsew signal input
rlabel metal3 s 99200 9256 100000 9376 6 sram1_dout1[0]
port 101 nsew signal input
rlabel metal3 s 99200 45704 100000 45824 6 sram1_dout1[10]
port 102 nsew signal input
rlabel metal3 s 99200 48288 100000 48408 6 sram1_dout1[11]
port 103 nsew signal input
rlabel metal3 s 99200 50872 100000 50992 6 sram1_dout1[12]
port 104 nsew signal input
rlabel metal3 s 99200 53320 100000 53440 6 sram1_dout1[13]
port 105 nsew signal input
rlabel metal3 s 99200 55904 100000 56024 6 sram1_dout1[14]
port 106 nsew signal input
rlabel metal3 s 99200 58488 100000 58608 6 sram1_dout1[15]
port 107 nsew signal input
rlabel metal3 s 99200 60936 100000 61056 6 sram1_dout1[16]
port 108 nsew signal input
rlabel metal3 s 99200 63520 100000 63640 6 sram1_dout1[17]
port 109 nsew signal input
rlabel metal3 s 99200 66104 100000 66224 6 sram1_dout1[18]
port 110 nsew signal input
rlabel metal3 s 99200 68552 100000 68672 6 sram1_dout1[19]
port 111 nsew signal input
rlabel metal3 s 99200 13336 100000 13456 6 sram1_dout1[1]
port 112 nsew signal input
rlabel metal3 s 99200 71136 100000 71256 6 sram1_dout1[20]
port 113 nsew signal input
rlabel metal3 s 99200 73584 100000 73704 6 sram1_dout1[21]
port 114 nsew signal input
rlabel metal3 s 99200 76168 100000 76288 6 sram1_dout1[22]
port 115 nsew signal input
rlabel metal3 s 99200 78752 100000 78872 6 sram1_dout1[23]
port 116 nsew signal input
rlabel metal3 s 99200 81200 100000 81320 6 sram1_dout1[24]
port 117 nsew signal input
rlabel metal3 s 99200 83784 100000 83904 6 sram1_dout1[25]
port 118 nsew signal input
rlabel metal3 s 99200 86368 100000 86488 6 sram1_dout1[26]
port 119 nsew signal input
rlabel metal3 s 99200 88816 100000 88936 6 sram1_dout1[27]
port 120 nsew signal input
rlabel metal3 s 99200 91400 100000 91520 6 sram1_dout1[28]
port 121 nsew signal input
rlabel metal3 s 99200 93984 100000 94104 6 sram1_dout1[29]
port 122 nsew signal input
rlabel metal3 s 99200 17280 100000 17400 6 sram1_dout1[2]
port 123 nsew signal input
rlabel metal3 s 99200 96432 100000 96552 6 sram1_dout1[30]
port 124 nsew signal input
rlabel metal3 s 99200 99016 100000 99136 6 sram1_dout1[31]
port 125 nsew signal input
rlabel metal3 s 99200 21360 100000 21480 6 sram1_dout1[3]
port 126 nsew signal input
rlabel metal3 s 99200 25440 100000 25560 6 sram1_dout1[4]
port 127 nsew signal input
rlabel metal3 s 99200 28976 100000 29096 6 sram1_dout1[5]
port 128 nsew signal input
rlabel metal3 s 99200 32512 100000 32632 6 sram1_dout1[6]
port 129 nsew signal input
rlabel metal3 s 99200 36048 100000 36168 6 sram1_dout1[7]
port 130 nsew signal input
rlabel metal3 s 99200 39720 100000 39840 6 sram1_dout1[8]
port 131 nsew signal input
rlabel metal3 s 99200 43256 100000 43376 6 sram1_dout1[9]
port 132 nsew signal input
rlabel metal3 s 99200 9664 100000 9784 6 sram_addr0[0]
port 133 nsew signal output
rlabel metal3 s 99200 13744 100000 13864 6 sram_addr0[1]
port 134 nsew signal output
rlabel metal3 s 99200 17824 100000 17944 6 sram_addr0[2]
port 135 nsew signal output
rlabel metal3 s 99200 21904 100000 22024 6 sram_addr0[3]
port 136 nsew signal output
rlabel metal3 s 99200 25984 100000 26104 6 sram_addr0[4]
port 137 nsew signal output
rlabel metal3 s 99200 29520 100000 29640 6 sram_addr0[5]
port 138 nsew signal output
rlabel metal3 s 99200 33056 100000 33176 6 sram_addr0[6]
port 139 nsew signal output
rlabel metal3 s 99200 36592 100000 36712 6 sram_addr0[7]
port 140 nsew signal output
rlabel metal3 s 99200 40128 100000 40248 6 sram_addr0[8]
port 141 nsew signal output
rlabel metal3 s 99200 10208 100000 10328 6 sram_addr1[0]
port 142 nsew signal output
rlabel metal3 s 99200 14288 100000 14408 6 sram_addr1[1]
port 143 nsew signal output
rlabel metal3 s 99200 18368 100000 18488 6 sram_addr1[2]
port 144 nsew signal output
rlabel metal3 s 99200 22448 100000 22568 6 sram_addr1[3]
port 145 nsew signal output
rlabel metal3 s 99200 26528 100000 26648 6 sram_addr1[4]
port 146 nsew signal output
rlabel metal3 s 99200 30064 100000 30184 6 sram_addr1[5]
port 147 nsew signal output
rlabel metal3 s 99200 33600 100000 33720 6 sram_addr1[6]
port 148 nsew signal output
rlabel metal3 s 99200 37136 100000 37256 6 sram_addr1[7]
port 149 nsew signal output
rlabel metal3 s 99200 40672 100000 40792 6 sram_addr1[8]
port 150 nsew signal output
rlabel metal3 s 99200 6128 100000 6248 6 sram_clk0
port 151 nsew signal output
rlabel metal3 s 99200 6672 100000 6792 6 sram_clk1
port 152 nsew signal output
rlabel metal3 s 99200 10752 100000 10872 6 sram_din0[0]
port 153 nsew signal output
rlabel metal3 s 99200 46248 100000 46368 6 sram_din0[10]
port 154 nsew signal output
rlabel metal3 s 99200 48832 100000 48952 6 sram_din0[11]
port 155 nsew signal output
rlabel metal3 s 99200 51280 100000 51400 6 sram_din0[12]
port 156 nsew signal output
rlabel metal3 s 99200 53864 100000 53984 6 sram_din0[13]
port 157 nsew signal output
rlabel metal3 s 99200 56448 100000 56568 6 sram_din0[14]
port 158 nsew signal output
rlabel metal3 s 99200 58896 100000 59016 6 sram_din0[15]
port 159 nsew signal output
rlabel metal3 s 99200 61480 100000 61600 6 sram_din0[16]
port 160 nsew signal output
rlabel metal3 s 99200 64064 100000 64184 6 sram_din0[17]
port 161 nsew signal output
rlabel metal3 s 99200 66512 100000 66632 6 sram_din0[18]
port 162 nsew signal output
rlabel metal3 s 99200 69096 100000 69216 6 sram_din0[19]
port 163 nsew signal output
rlabel metal3 s 99200 14832 100000 14952 6 sram_din0[1]
port 164 nsew signal output
rlabel metal3 s 99200 71680 100000 71800 6 sram_din0[20]
port 165 nsew signal output
rlabel metal3 s 99200 74128 100000 74248 6 sram_din0[21]
port 166 nsew signal output
rlabel metal3 s 99200 76712 100000 76832 6 sram_din0[22]
port 167 nsew signal output
rlabel metal3 s 99200 79296 100000 79416 6 sram_din0[23]
port 168 nsew signal output
rlabel metal3 s 99200 81744 100000 81864 6 sram_din0[24]
port 169 nsew signal output
rlabel metal3 s 99200 84328 100000 84448 6 sram_din0[25]
port 170 nsew signal output
rlabel metal3 s 99200 86776 100000 86896 6 sram_din0[26]
port 171 nsew signal output
rlabel metal3 s 99200 89360 100000 89480 6 sram_din0[27]
port 172 nsew signal output
rlabel metal3 s 99200 91944 100000 92064 6 sram_din0[28]
port 173 nsew signal output
rlabel metal3 s 99200 94392 100000 94512 6 sram_din0[29]
port 174 nsew signal output
rlabel metal3 s 99200 18912 100000 19032 6 sram_din0[2]
port 175 nsew signal output
rlabel metal3 s 99200 96976 100000 97096 6 sram_din0[30]
port 176 nsew signal output
rlabel metal3 s 99200 99560 100000 99680 6 sram_din0[31]
port 177 nsew signal output
rlabel metal3 s 99200 22856 100000 22976 6 sram_din0[3]
port 178 nsew signal output
rlabel metal3 s 99200 26936 100000 27056 6 sram_din0[4]
port 179 nsew signal output
rlabel metal3 s 99200 30472 100000 30592 6 sram_din0[5]
port 180 nsew signal output
rlabel metal3 s 99200 34008 100000 34128 6 sram_din0[6]
port 181 nsew signal output
rlabel metal3 s 99200 37680 100000 37800 6 sram_din0[7]
port 182 nsew signal output
rlabel metal3 s 99200 41216 100000 41336 6 sram_din0[8]
port 183 nsew signal output
rlabel metal3 s 99200 43664 100000 43784 6 sram_din0[9]
port 184 nsew signal output
rlabel metal3 s 99200 7216 100000 7336 6 sram_web0
port 185 nsew signal output
rlabel metal3 s 99200 11296 100000 11416 6 sram_wmask0[0]
port 186 nsew signal output
rlabel metal3 s 99200 15240 100000 15360 6 sram_wmask0[1]
port 187 nsew signal output
rlabel metal3 s 99200 19320 100000 19440 6 sram_wmask0[2]
port 188 nsew signal output
rlabel metal3 s 99200 23400 100000 23520 6 sram_wmask0[3]
port 189 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 190 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 190 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 190 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 190 nsew power input
rlabel metal3 s 99200 1096 100000 1216 6 vga_b[0]
port 191 nsew signal output
rlabel metal3 s 99200 2592 100000 2712 6 vga_b[1]
port 192 nsew signal output
rlabel metal3 s 99200 1640 100000 1760 6 vga_g[0]
port 193 nsew signal output
rlabel metal3 s 99200 3136 100000 3256 6 vga_g[1]
port 194 nsew signal output
rlabel metal3 s 99200 144 100000 264 6 vga_hsync
port 195 nsew signal output
rlabel metal3 s 99200 2048 100000 2168 6 vga_r[0]
port 196 nsew signal output
rlabel metal3 s 99200 3680 100000 3800 6 vga_r[1]
port 197 nsew signal output
rlabel metal3 s 99200 552 100000 672 6 vga_vsync
port 198 nsew signal output
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 199 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 199 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 199 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_ack_o
port 200 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wb_adr_i[0]
port 201 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wb_adr_i[10]
port 202 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wb_adr_i[11]
port 203 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 wb_adr_i[12]
port 204 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 wb_adr_i[13]
port 205 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wb_adr_i[14]
port 206 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wb_adr_i[15]
port 207 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 wb_adr_i[16]
port 208 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wb_adr_i[17]
port 209 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 wb_adr_i[18]
port 210 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 wb_adr_i[19]
port 211 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wb_adr_i[1]
port 212 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 wb_adr_i[20]
port 213 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 wb_adr_i[21]
port 214 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 wb_adr_i[22]
port 215 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 wb_adr_i[23]
port 216 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wb_adr_i[2]
port 217 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wb_adr_i[3]
port 218 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wb_adr_i[4]
port 219 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wb_adr_i[5]
port 220 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wb_adr_i[6]
port 221 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wb_adr_i[7]
port 222 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wb_adr_i[8]
port 223 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wb_adr_i[9]
port 224 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_clk_i
port 225 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wb_cyc_i
port 226 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wb_data_i[0]
port 227 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wb_data_i[10]
port 228 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wb_data_i[11]
port 229 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wb_data_i[12]
port 230 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wb_data_i[13]
port 231 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wb_data_i[14]
port 232 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wb_data_i[15]
port 233 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 wb_data_i[16]
port 234 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 wb_data_i[17]
port 235 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wb_data_i[18]
port 236 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 wb_data_i[19]
port 237 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wb_data_i[1]
port 238 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 wb_data_i[20]
port 239 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 wb_data_i[21]
port 240 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 wb_data_i[22]
port 241 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 wb_data_i[23]
port 242 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 wb_data_i[24]
port 243 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 wb_data_i[25]
port 244 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 wb_data_i[26]
port 245 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 wb_data_i[27]
port 246 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 wb_data_i[28]
port 247 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 wb_data_i[29]
port 248 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wb_data_i[2]
port 249 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 wb_data_i[30]
port 250 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 wb_data_i[31]
port 251 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wb_data_i[3]
port 252 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wb_data_i[4]
port 253 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wb_data_i[5]
port 254 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wb_data_i[6]
port 255 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wb_data_i[7]
port 256 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wb_data_i[8]
port 257 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wb_data_i[9]
port 258 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wb_data_o[0]
port 259 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 wb_data_o[10]
port 260 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 wb_data_o[11]
port 261 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 wb_data_o[12]
port 262 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 wb_data_o[13]
port 263 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 wb_data_o[14]
port 264 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 wb_data_o[15]
port 265 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 wb_data_o[16]
port 266 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 wb_data_o[17]
port 267 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 wb_data_o[18]
port 268 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 wb_data_o[19]
port 269 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wb_data_o[1]
port 270 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 wb_data_o[20]
port 271 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 wb_data_o[21]
port 272 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 wb_data_o[22]
port 273 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 wb_data_o[23]
port 274 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 wb_data_o[24]
port 275 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 wb_data_o[25]
port 276 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 wb_data_o[26]
port 277 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 wb_data_o[27]
port 278 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 wb_data_o[28]
port 279 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 wb_data_o[29]
port 280 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wb_data_o[2]
port 281 nsew signal output
rlabel metal2 s 97446 0 97502 800 6 wb_data_o[30]
port 282 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 wb_data_o[31]
port 283 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wb_data_o[3]
port 284 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 wb_data_o[4]
port 285 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wb_data_o[5]
port 286 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 wb_data_o[6]
port 287 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wb_data_o[7]
port 288 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wb_data_o[8]
port 289 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 wb_data_o[9]
port 290 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 wb_error_o
port 291 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wb_rst_i
port 292 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wb_sel_i[0]
port 293 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wb_sel_i[1]
port 294 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wb_sel_i[2]
port 295 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wb_sel_i[3]
port 296 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wb_stall_o
port 297 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 wb_stb_i
port 298 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wb_we_i
port 299 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6592686
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Video/runs/Video/results/finishing/Video.magic.gds
string GDS_START 572064
<< end >>

