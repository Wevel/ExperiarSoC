VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO GPIO
  CLASS BLOCK ;
  FOREIGN GPIO ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END clk
  PIN gpio0_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1.400 200.000 2.000 ;
    END
  END gpio0_input[0]
  PIN gpio0_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 106.120 200.000 106.720 ;
    END
  END gpio0_input[10]
  PIN gpio0_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 117.000 200.000 117.600 ;
    END
  END gpio0_input[11]
  PIN gpio0_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 127.200 200.000 127.800 ;
    END
  END gpio0_input[12]
  PIN gpio0_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 138.080 200.000 138.680 ;
    END
  END gpio0_input[13]
  PIN gpio0_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 148.280 200.000 148.880 ;
    END
  END gpio0_input[14]
  PIN gpio0_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 159.160 200.000 159.760 ;
    END
  END gpio0_input[15]
  PIN gpio0_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 169.360 200.000 169.960 ;
    END
  END gpio0_input[16]
  PIN gpio0_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 180.240 200.000 180.840 ;
    END
  END gpio0_input[17]
  PIN gpio0_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 190.440 200.000 191.040 ;
    END
  END gpio0_input[18]
  PIN gpio0_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 11.600 200.000 12.200 ;
    END
  END gpio0_input[1]
  PIN gpio0_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 21.800 200.000 22.400 ;
    END
  END gpio0_input[2]
  PIN gpio0_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 32.680 200.000 33.280 ;
    END
  END gpio0_input[3]
  PIN gpio0_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 42.880 200.000 43.480 ;
    END
  END gpio0_input[4]
  PIN gpio0_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 53.760 200.000 54.360 ;
    END
  END gpio0_input[5]
  PIN gpio0_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 63.960 200.000 64.560 ;
    END
  END gpio0_input[6]
  PIN gpio0_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 74.840 200.000 75.440 ;
    END
  END gpio0_input[7]
  PIN gpio0_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 85.040 200.000 85.640 ;
    END
  END gpio0_input[8]
  PIN gpio0_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.920 200.000 96.520 ;
    END
  END gpio0_input[9]
  PIN gpio0_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 4.800 200.000 5.400 ;
    END
  END gpio0_oe[0]
  PIN gpio0_oe[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 109.520 200.000 110.120 ;
    END
  END gpio0_oe[10]
  PIN gpio0_oe[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 120.400 200.000 121.000 ;
    END
  END gpio0_oe[11]
  PIN gpio0_oe[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 130.600 200.000 131.200 ;
    END
  END gpio0_oe[12]
  PIN gpio0_oe[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 141.480 200.000 142.080 ;
    END
  END gpio0_oe[13]
  PIN gpio0_oe[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 151.680 200.000 152.280 ;
    END
  END gpio0_oe[14]
  PIN gpio0_oe[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 162.560 200.000 163.160 ;
    END
  END gpio0_oe[15]
  PIN gpio0_oe[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 172.760 200.000 173.360 ;
    END
  END gpio0_oe[16]
  PIN gpio0_oe[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 183.640 200.000 184.240 ;
    END
  END gpio0_oe[17]
  PIN gpio0_oe[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 193.840 200.000 194.440 ;
    END
  END gpio0_oe[18]
  PIN gpio0_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 15.000 200.000 15.600 ;
    END
  END gpio0_oe[1]
  PIN gpio0_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 25.880 200.000 26.480 ;
    END
  END gpio0_oe[2]
  PIN gpio0_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 36.080 200.000 36.680 ;
    END
  END gpio0_oe[3]
  PIN gpio0_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 46.960 200.000 47.560 ;
    END
  END gpio0_oe[4]
  PIN gpio0_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 57.160 200.000 57.760 ;
    END
  END gpio0_oe[5]
  PIN gpio0_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 68.040 200.000 68.640 ;
    END
  END gpio0_oe[6]
  PIN gpio0_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.240 200.000 78.840 ;
    END
  END gpio0_oe[7]
  PIN gpio0_oe[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 88.440 200.000 89.040 ;
    END
  END gpio0_oe[8]
  PIN gpio0_oe[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 99.320 200.000 99.920 ;
    END
  END gpio0_oe[9]
  PIN gpio0_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 8.200 200.000 8.800 ;
    END
  END gpio0_output[0]
  PIN gpio0_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 113.600 200.000 114.200 ;
    END
  END gpio0_output[10]
  PIN gpio0_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 123.800 200.000 124.400 ;
    END
  END gpio0_output[11]
  PIN gpio0_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 134.680 200.000 135.280 ;
    END
  END gpio0_output[12]
  PIN gpio0_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 144.880 200.000 145.480 ;
    END
  END gpio0_output[13]
  PIN gpio0_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 155.080 200.000 155.680 ;
    END
  END gpio0_output[14]
  PIN gpio0_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 165.960 200.000 166.560 ;
    END
  END gpio0_output[15]
  PIN gpio0_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.160 200.000 176.760 ;
    END
  END gpio0_output[16]
  PIN gpio0_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.040 200.000 187.640 ;
    END
  END gpio0_output[17]
  PIN gpio0_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 197.240 200.000 197.840 ;
    END
  END gpio0_output[18]
  PIN gpio0_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 18.400 200.000 19.000 ;
    END
  END gpio0_output[1]
  PIN gpio0_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 29.280 200.000 29.880 ;
    END
  END gpio0_output[2]
  PIN gpio0_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 39.480 200.000 40.080 ;
    END
  END gpio0_output[3]
  PIN gpio0_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 50.360 200.000 50.960 ;
    END
  END gpio0_output[4]
  PIN gpio0_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 60.560 200.000 61.160 ;
    END
  END gpio0_output[5]
  PIN gpio0_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 71.440 200.000 72.040 ;
    END
  END gpio0_output[6]
  PIN gpio0_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 81.640 200.000 82.240 ;
    END
  END gpio0_output[7]
  PIN gpio0_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 92.520 200.000 93.120 ;
    END
  END gpio0_output[8]
  PIN gpio0_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 102.720 200.000 103.320 ;
    END
  END gpio0_output[9]
  PIN gpio1_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END gpio1_input[0]
  PIN gpio1_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END gpio1_input[10]
  PIN gpio1_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END gpio1_input[11]
  PIN gpio1_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END gpio1_input[12]
  PIN gpio1_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END gpio1_input[13]
  PIN gpio1_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END gpio1_input[14]
  PIN gpio1_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END gpio1_input[15]
  PIN gpio1_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END gpio1_input[16]
  PIN gpio1_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END gpio1_input[17]
  PIN gpio1_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END gpio1_input[18]
  PIN gpio1_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END gpio1_input[1]
  PIN gpio1_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END gpio1_input[2]
  PIN gpio1_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END gpio1_input[3]
  PIN gpio1_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gpio1_input[4]
  PIN gpio1_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END gpio1_input[5]
  PIN gpio1_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END gpio1_input[6]
  PIN gpio1_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END gpio1_input[7]
  PIN gpio1_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END gpio1_input[8]
  PIN gpio1_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END gpio1_input[9]
  PIN gpio1_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END gpio1_oe[0]
  PIN gpio1_oe[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END gpio1_oe[10]
  PIN gpio1_oe[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END gpio1_oe[11]
  PIN gpio1_oe[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END gpio1_oe[12]
  PIN gpio1_oe[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END gpio1_oe[13]
  PIN gpio1_oe[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END gpio1_oe[14]
  PIN gpio1_oe[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END gpio1_oe[15]
  PIN gpio1_oe[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END gpio1_oe[16]
  PIN gpio1_oe[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END gpio1_oe[17]
  PIN gpio1_oe[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END gpio1_oe[18]
  PIN gpio1_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END gpio1_oe[1]
  PIN gpio1_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END gpio1_oe[2]
  PIN gpio1_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END gpio1_oe[3]
  PIN gpio1_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END gpio1_oe[4]
  PIN gpio1_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END gpio1_oe[5]
  PIN gpio1_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END gpio1_oe[6]
  PIN gpio1_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END gpio1_oe[7]
  PIN gpio1_oe[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END gpio1_oe[8]
  PIN gpio1_oe[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END gpio1_oe[9]
  PIN gpio1_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END gpio1_output[0]
  PIN gpio1_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END gpio1_output[10]
  PIN gpio1_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END gpio1_output[11]
  PIN gpio1_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END gpio1_output[12]
  PIN gpio1_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END gpio1_output[13]
  PIN gpio1_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END gpio1_output[14]
  PIN gpio1_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END gpio1_output[15]
  PIN gpio1_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END gpio1_output[16]
  PIN gpio1_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END gpio1_output[17]
  PIN gpio1_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END gpio1_output[18]
  PIN gpio1_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END gpio1_output[1]
  PIN gpio1_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END gpio1_output[2]
  PIN gpio1_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END gpio1_output[3]
  PIN gpio1_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END gpio1_output[4]
  PIN gpio1_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END gpio1_output[5]
  PIN gpio1_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END gpio1_output[6]
  PIN gpio1_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END gpio1_output[7]
  PIN gpio1_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END gpio1_output[8]
  PIN gpio1_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END gpio1_output[9]
  PIN peripheralBus_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END peripheralBus_address[0]
  PIN peripheralBus_address[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END peripheralBus_address[10]
  PIN peripheralBus_address[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END peripheralBus_address[11]
  PIN peripheralBus_address[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END peripheralBus_address[12]
  PIN peripheralBus_address[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END peripheralBus_address[13]
  PIN peripheralBus_address[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END peripheralBus_address[14]
  PIN peripheralBus_address[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END peripheralBus_address[15]
  PIN peripheralBus_address[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END peripheralBus_address[16]
  PIN peripheralBus_address[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END peripheralBus_address[17]
  PIN peripheralBus_address[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END peripheralBus_address[18]
  PIN peripheralBus_address[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END peripheralBus_address[19]
  PIN peripheralBus_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END peripheralBus_address[1]
  PIN peripheralBus_address[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END peripheralBus_address[20]
  PIN peripheralBus_address[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END peripheralBus_address[21]
  PIN peripheralBus_address[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END peripheralBus_address[22]
  PIN peripheralBus_address[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END peripheralBus_address[23]
  PIN peripheralBus_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END peripheralBus_address[2]
  PIN peripheralBus_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END peripheralBus_address[3]
  PIN peripheralBus_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END peripheralBus_address[4]
  PIN peripheralBus_address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END peripheralBus_address[5]
  PIN peripheralBus_address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END peripheralBus_address[6]
  PIN peripheralBus_address[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END peripheralBus_address[7]
  PIN peripheralBus_address[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END peripheralBus_address[8]
  PIN peripheralBus_address[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END peripheralBus_address[9]
  PIN peripheralBus_busy
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END peripheralBus_busy
  PIN peripheralBus_dataIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END peripheralBus_dataIn[0]
  PIN peripheralBus_dataIn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END peripheralBus_dataIn[10]
  PIN peripheralBus_dataIn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END peripheralBus_dataIn[11]
  PIN peripheralBus_dataIn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END peripheralBus_dataIn[12]
  PIN peripheralBus_dataIn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END peripheralBus_dataIn[13]
  PIN peripheralBus_dataIn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END peripheralBus_dataIn[14]
  PIN peripheralBus_dataIn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END peripheralBus_dataIn[15]
  PIN peripheralBus_dataIn[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END peripheralBus_dataIn[16]
  PIN peripheralBus_dataIn[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END peripheralBus_dataIn[17]
  PIN peripheralBus_dataIn[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END peripheralBus_dataIn[18]
  PIN peripheralBus_dataIn[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END peripheralBus_dataIn[19]
  PIN peripheralBus_dataIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END peripheralBus_dataIn[1]
  PIN peripheralBus_dataIn[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END peripheralBus_dataIn[20]
  PIN peripheralBus_dataIn[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END peripheralBus_dataIn[21]
  PIN peripheralBus_dataIn[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END peripheralBus_dataIn[22]
  PIN peripheralBus_dataIn[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END peripheralBus_dataIn[23]
  PIN peripheralBus_dataIn[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END peripheralBus_dataIn[24]
  PIN peripheralBus_dataIn[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END peripheralBus_dataIn[25]
  PIN peripheralBus_dataIn[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END peripheralBus_dataIn[26]
  PIN peripheralBus_dataIn[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END peripheralBus_dataIn[27]
  PIN peripheralBus_dataIn[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END peripheralBus_dataIn[28]
  PIN peripheralBus_dataIn[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END peripheralBus_dataIn[29]
  PIN peripheralBus_dataIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END peripheralBus_dataIn[2]
  PIN peripheralBus_dataIn[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END peripheralBus_dataIn[30]
  PIN peripheralBus_dataIn[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END peripheralBus_dataIn[31]
  PIN peripheralBus_dataIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END peripheralBus_dataIn[3]
  PIN peripheralBus_dataIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END peripheralBus_dataIn[4]
  PIN peripheralBus_dataIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END peripheralBus_dataIn[5]
  PIN peripheralBus_dataIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END peripheralBus_dataIn[6]
  PIN peripheralBus_dataIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END peripheralBus_dataIn[7]
  PIN peripheralBus_dataIn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END peripheralBus_dataIn[8]
  PIN peripheralBus_dataIn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END peripheralBus_dataIn[9]
  PIN peripheralBus_dataOut[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END peripheralBus_dataOut[0]
  PIN peripheralBus_dataOut[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END peripheralBus_dataOut[10]
  PIN peripheralBus_dataOut[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END peripheralBus_dataOut[11]
  PIN peripheralBus_dataOut[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END peripheralBus_dataOut[12]
  PIN peripheralBus_dataOut[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END peripheralBus_dataOut[13]
  PIN peripheralBus_dataOut[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END peripheralBus_dataOut[14]
  PIN peripheralBus_dataOut[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END peripheralBus_dataOut[15]
  PIN peripheralBus_dataOut[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END peripheralBus_dataOut[16]
  PIN peripheralBus_dataOut[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END peripheralBus_dataOut[17]
  PIN peripheralBus_dataOut[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END peripheralBus_dataOut[18]
  PIN peripheralBus_dataOut[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END peripheralBus_dataOut[19]
  PIN peripheralBus_dataOut[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END peripheralBus_dataOut[1]
  PIN peripheralBus_dataOut[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END peripheralBus_dataOut[20]
  PIN peripheralBus_dataOut[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END peripheralBus_dataOut[21]
  PIN peripheralBus_dataOut[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END peripheralBus_dataOut[22]
  PIN peripheralBus_dataOut[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END peripheralBus_dataOut[23]
  PIN peripheralBus_dataOut[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END peripheralBus_dataOut[24]
  PIN peripheralBus_dataOut[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END peripheralBus_dataOut[25]
  PIN peripheralBus_dataOut[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END peripheralBus_dataOut[26]
  PIN peripheralBus_dataOut[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END peripheralBus_dataOut[27]
  PIN peripheralBus_dataOut[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END peripheralBus_dataOut[28]
  PIN peripheralBus_dataOut[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END peripheralBus_dataOut[29]
  PIN peripheralBus_dataOut[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END peripheralBus_dataOut[2]
  PIN peripheralBus_dataOut[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END peripheralBus_dataOut[30]
  PIN peripheralBus_dataOut[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END peripheralBus_dataOut[31]
  PIN peripheralBus_dataOut[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END peripheralBus_dataOut[3]
  PIN peripheralBus_dataOut[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END peripheralBus_dataOut[4]
  PIN peripheralBus_dataOut[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END peripheralBus_dataOut[5]
  PIN peripheralBus_dataOut[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END peripheralBus_dataOut[6]
  PIN peripheralBus_dataOut[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END peripheralBus_dataOut[7]
  PIN peripheralBus_dataOut[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END peripheralBus_dataOut[8]
  PIN peripheralBus_dataOut[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END peripheralBus_dataOut[9]
  PIN peripheralBus_oe
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END peripheralBus_oe
  PIN peripheralBus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END peripheralBus_we
  PIN requestOutput
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 196.000 100.190 200.000 ;
    END
  END requestOutput
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 1.450 1.060 198.190 187.920 ;
      LAYER met2 ;
        RECT 1.480 195.720 99.630 198.405 ;
        RECT 100.470 195.720 198.160 198.405 ;
        RECT 1.480 4.280 198.160 195.720 ;
        RECT 2.030 0.835 4.410 4.280 ;
        RECT 5.250 0.835 7.630 4.280 ;
        RECT 8.470 0.835 11.310 4.280 ;
        RECT 12.150 0.835 14.530 4.280 ;
        RECT 15.370 0.835 17.750 4.280 ;
        RECT 18.590 0.835 21.430 4.280 ;
        RECT 22.270 0.835 24.650 4.280 ;
        RECT 25.490 0.835 27.870 4.280 ;
        RECT 28.710 0.835 31.550 4.280 ;
        RECT 32.390 0.835 34.770 4.280 ;
        RECT 35.610 0.835 38.450 4.280 ;
        RECT 39.290 0.835 41.670 4.280 ;
        RECT 42.510 0.835 44.890 4.280 ;
        RECT 45.730 0.835 48.570 4.280 ;
        RECT 49.410 0.835 51.790 4.280 ;
        RECT 52.630 0.835 55.010 4.280 ;
        RECT 55.850 0.835 58.690 4.280 ;
        RECT 59.530 0.835 61.910 4.280 ;
        RECT 62.750 0.835 65.590 4.280 ;
        RECT 66.430 0.835 68.810 4.280 ;
        RECT 69.650 0.835 72.030 4.280 ;
        RECT 72.870 0.835 75.710 4.280 ;
        RECT 76.550 0.835 78.930 4.280 ;
        RECT 79.770 0.835 82.150 4.280 ;
        RECT 82.990 0.835 85.830 4.280 ;
        RECT 86.670 0.835 89.050 4.280 ;
        RECT 89.890 0.835 92.730 4.280 ;
        RECT 93.570 0.835 95.950 4.280 ;
        RECT 96.790 0.835 99.170 4.280 ;
        RECT 100.010 0.835 102.850 4.280 ;
        RECT 103.690 0.835 106.070 4.280 ;
        RECT 106.910 0.835 109.290 4.280 ;
        RECT 110.130 0.835 112.970 4.280 ;
        RECT 113.810 0.835 116.190 4.280 ;
        RECT 117.030 0.835 119.870 4.280 ;
        RECT 120.710 0.835 123.090 4.280 ;
        RECT 123.930 0.835 126.310 4.280 ;
        RECT 127.150 0.835 129.990 4.280 ;
        RECT 130.830 0.835 133.210 4.280 ;
        RECT 134.050 0.835 136.430 4.280 ;
        RECT 137.270 0.835 140.110 4.280 ;
        RECT 140.950 0.835 143.330 4.280 ;
        RECT 144.170 0.835 147.010 4.280 ;
        RECT 147.850 0.835 150.230 4.280 ;
        RECT 151.070 0.835 153.450 4.280 ;
        RECT 154.290 0.835 157.130 4.280 ;
        RECT 157.970 0.835 160.350 4.280 ;
        RECT 161.190 0.835 163.570 4.280 ;
        RECT 164.410 0.835 167.250 4.280 ;
        RECT 168.090 0.835 170.470 4.280 ;
        RECT 171.310 0.835 174.150 4.280 ;
        RECT 174.990 0.835 177.370 4.280 ;
        RECT 178.210 0.835 180.590 4.280 ;
        RECT 181.430 0.835 184.270 4.280 ;
        RECT 185.110 0.835 187.490 4.280 ;
        RECT 188.330 0.835 190.710 4.280 ;
        RECT 191.550 0.835 194.390 4.280 ;
        RECT 195.230 0.835 197.610 4.280 ;
      LAYER met3 ;
        RECT 4.400 198.240 196.000 198.385 ;
        RECT 4.400 197.520 195.600 198.240 ;
        RECT 4.000 196.880 195.600 197.520 ;
        RECT 4.400 196.840 195.600 196.880 ;
        RECT 4.400 195.480 196.000 196.840 ;
        RECT 4.000 194.840 196.000 195.480 ;
        RECT 4.400 193.440 195.600 194.840 ;
        RECT 4.000 192.800 196.000 193.440 ;
        RECT 4.400 191.440 196.000 192.800 ;
        RECT 4.400 191.400 195.600 191.440 ;
        RECT 4.000 190.080 195.600 191.400 ;
        RECT 4.400 190.040 195.600 190.080 ;
        RECT 4.400 188.680 196.000 190.040 ;
        RECT 4.000 188.040 196.000 188.680 ;
        RECT 4.400 186.640 195.600 188.040 ;
        RECT 4.000 186.000 196.000 186.640 ;
        RECT 4.400 184.640 196.000 186.000 ;
        RECT 4.400 184.600 195.600 184.640 ;
        RECT 4.000 183.960 195.600 184.600 ;
        RECT 4.400 183.240 195.600 183.960 ;
        RECT 4.400 182.560 196.000 183.240 ;
        RECT 4.000 181.240 196.000 182.560 ;
        RECT 4.400 179.840 195.600 181.240 ;
        RECT 4.000 179.200 196.000 179.840 ;
        RECT 4.400 177.800 196.000 179.200 ;
        RECT 4.000 177.160 196.000 177.800 ;
        RECT 4.400 175.760 195.600 177.160 ;
        RECT 4.000 175.120 196.000 175.760 ;
        RECT 4.400 173.760 196.000 175.120 ;
        RECT 4.400 173.720 195.600 173.760 ;
        RECT 4.000 173.080 195.600 173.720 ;
        RECT 4.400 172.360 195.600 173.080 ;
        RECT 4.400 171.680 196.000 172.360 ;
        RECT 4.000 170.360 196.000 171.680 ;
        RECT 4.400 168.960 195.600 170.360 ;
        RECT 4.000 168.320 196.000 168.960 ;
        RECT 4.400 166.960 196.000 168.320 ;
        RECT 4.400 166.920 195.600 166.960 ;
        RECT 4.000 166.280 195.600 166.920 ;
        RECT 4.400 165.560 195.600 166.280 ;
        RECT 4.400 164.880 196.000 165.560 ;
        RECT 4.000 164.240 196.000 164.880 ;
        RECT 4.400 163.560 196.000 164.240 ;
        RECT 4.400 162.840 195.600 163.560 ;
        RECT 4.000 162.160 195.600 162.840 ;
        RECT 4.000 161.520 196.000 162.160 ;
        RECT 4.400 160.160 196.000 161.520 ;
        RECT 4.400 160.120 195.600 160.160 ;
        RECT 4.000 159.480 195.600 160.120 ;
        RECT 4.400 158.760 195.600 159.480 ;
        RECT 4.400 158.080 196.000 158.760 ;
        RECT 4.000 157.440 196.000 158.080 ;
        RECT 4.400 156.080 196.000 157.440 ;
        RECT 4.400 156.040 195.600 156.080 ;
        RECT 4.000 155.400 195.600 156.040 ;
        RECT 4.400 154.680 195.600 155.400 ;
        RECT 4.400 154.000 196.000 154.680 ;
        RECT 4.000 152.680 196.000 154.000 ;
        RECT 4.400 151.280 195.600 152.680 ;
        RECT 4.000 150.640 196.000 151.280 ;
        RECT 4.400 149.280 196.000 150.640 ;
        RECT 4.400 149.240 195.600 149.280 ;
        RECT 4.000 148.600 195.600 149.240 ;
        RECT 4.400 147.880 195.600 148.600 ;
        RECT 4.400 147.200 196.000 147.880 ;
        RECT 4.000 146.560 196.000 147.200 ;
        RECT 4.400 145.880 196.000 146.560 ;
        RECT 4.400 145.160 195.600 145.880 ;
        RECT 4.000 144.520 195.600 145.160 ;
        RECT 4.400 144.480 195.600 144.520 ;
        RECT 4.400 143.120 196.000 144.480 ;
        RECT 4.000 142.480 196.000 143.120 ;
        RECT 4.000 141.800 195.600 142.480 ;
        RECT 4.400 141.080 195.600 141.800 ;
        RECT 4.400 140.400 196.000 141.080 ;
        RECT 4.000 139.760 196.000 140.400 ;
        RECT 4.400 139.080 196.000 139.760 ;
        RECT 4.400 138.360 195.600 139.080 ;
        RECT 4.000 137.720 195.600 138.360 ;
        RECT 4.400 137.680 195.600 137.720 ;
        RECT 4.400 136.320 196.000 137.680 ;
        RECT 4.000 135.680 196.000 136.320 ;
        RECT 4.400 134.280 195.600 135.680 ;
        RECT 4.000 132.960 196.000 134.280 ;
        RECT 4.400 131.600 196.000 132.960 ;
        RECT 4.400 131.560 195.600 131.600 ;
        RECT 4.000 130.920 195.600 131.560 ;
        RECT 4.400 130.200 195.600 130.920 ;
        RECT 4.400 129.520 196.000 130.200 ;
        RECT 4.000 128.880 196.000 129.520 ;
        RECT 4.400 128.200 196.000 128.880 ;
        RECT 4.400 127.480 195.600 128.200 ;
        RECT 4.000 126.840 195.600 127.480 ;
        RECT 4.400 126.800 195.600 126.840 ;
        RECT 4.400 125.440 196.000 126.800 ;
        RECT 4.000 124.800 196.000 125.440 ;
        RECT 4.000 124.120 195.600 124.800 ;
        RECT 4.400 123.400 195.600 124.120 ;
        RECT 4.400 122.720 196.000 123.400 ;
        RECT 4.000 122.080 196.000 122.720 ;
        RECT 4.400 121.400 196.000 122.080 ;
        RECT 4.400 120.680 195.600 121.400 ;
        RECT 4.000 120.040 195.600 120.680 ;
        RECT 4.400 120.000 195.600 120.040 ;
        RECT 4.400 118.640 196.000 120.000 ;
        RECT 4.000 118.000 196.000 118.640 ;
        RECT 4.400 116.600 195.600 118.000 ;
        RECT 4.000 115.960 196.000 116.600 ;
        RECT 4.400 114.600 196.000 115.960 ;
        RECT 4.400 114.560 195.600 114.600 ;
        RECT 4.000 113.240 195.600 114.560 ;
        RECT 4.400 113.200 195.600 113.240 ;
        RECT 4.400 111.840 196.000 113.200 ;
        RECT 4.000 111.200 196.000 111.840 ;
        RECT 4.400 110.520 196.000 111.200 ;
        RECT 4.400 109.800 195.600 110.520 ;
        RECT 4.000 109.160 195.600 109.800 ;
        RECT 4.400 109.120 195.600 109.160 ;
        RECT 4.400 107.760 196.000 109.120 ;
        RECT 4.000 107.120 196.000 107.760 ;
        RECT 4.400 105.720 195.600 107.120 ;
        RECT 4.000 104.400 196.000 105.720 ;
        RECT 4.400 103.720 196.000 104.400 ;
        RECT 4.400 103.000 195.600 103.720 ;
        RECT 4.000 102.360 195.600 103.000 ;
        RECT 4.400 102.320 195.600 102.360 ;
        RECT 4.400 100.960 196.000 102.320 ;
        RECT 4.000 100.320 196.000 100.960 ;
        RECT 4.400 98.920 195.600 100.320 ;
        RECT 4.000 98.280 196.000 98.920 ;
        RECT 4.400 96.920 196.000 98.280 ;
        RECT 4.400 96.880 195.600 96.920 ;
        RECT 4.000 95.560 195.600 96.880 ;
        RECT 4.400 95.520 195.600 95.560 ;
        RECT 4.400 94.160 196.000 95.520 ;
        RECT 4.000 93.520 196.000 94.160 ;
        RECT 4.400 92.120 195.600 93.520 ;
        RECT 4.000 91.480 196.000 92.120 ;
        RECT 4.400 90.080 196.000 91.480 ;
        RECT 4.000 89.440 196.000 90.080 ;
        RECT 4.400 88.040 195.600 89.440 ;
        RECT 4.000 87.400 196.000 88.040 ;
        RECT 4.400 86.040 196.000 87.400 ;
        RECT 4.400 86.000 195.600 86.040 ;
        RECT 4.000 84.680 195.600 86.000 ;
        RECT 4.400 84.640 195.600 84.680 ;
        RECT 4.400 83.280 196.000 84.640 ;
        RECT 4.000 82.640 196.000 83.280 ;
        RECT 4.400 81.240 195.600 82.640 ;
        RECT 4.000 80.600 196.000 81.240 ;
        RECT 4.400 79.240 196.000 80.600 ;
        RECT 4.400 79.200 195.600 79.240 ;
        RECT 4.000 78.560 195.600 79.200 ;
        RECT 4.400 77.840 195.600 78.560 ;
        RECT 4.400 77.160 196.000 77.840 ;
        RECT 4.000 75.840 196.000 77.160 ;
        RECT 4.400 74.440 195.600 75.840 ;
        RECT 4.000 73.800 196.000 74.440 ;
        RECT 4.400 72.440 196.000 73.800 ;
        RECT 4.400 72.400 195.600 72.440 ;
        RECT 4.000 71.760 195.600 72.400 ;
        RECT 4.400 71.040 195.600 71.760 ;
        RECT 4.400 70.360 196.000 71.040 ;
        RECT 4.000 69.720 196.000 70.360 ;
        RECT 4.400 69.040 196.000 69.720 ;
        RECT 4.400 68.320 195.600 69.040 ;
        RECT 4.000 67.640 195.600 68.320 ;
        RECT 4.000 67.000 196.000 67.640 ;
        RECT 4.400 65.600 196.000 67.000 ;
        RECT 4.000 64.960 196.000 65.600 ;
        RECT 4.400 63.560 195.600 64.960 ;
        RECT 4.000 62.920 196.000 63.560 ;
        RECT 4.400 61.560 196.000 62.920 ;
        RECT 4.400 61.520 195.600 61.560 ;
        RECT 4.000 60.880 195.600 61.520 ;
        RECT 4.400 60.160 195.600 60.880 ;
        RECT 4.400 59.480 196.000 60.160 ;
        RECT 4.000 58.840 196.000 59.480 ;
        RECT 4.400 58.160 196.000 58.840 ;
        RECT 4.400 57.440 195.600 58.160 ;
        RECT 4.000 56.760 195.600 57.440 ;
        RECT 4.000 56.120 196.000 56.760 ;
        RECT 4.400 54.760 196.000 56.120 ;
        RECT 4.400 54.720 195.600 54.760 ;
        RECT 4.000 54.080 195.600 54.720 ;
        RECT 4.400 53.360 195.600 54.080 ;
        RECT 4.400 52.680 196.000 53.360 ;
        RECT 4.000 52.040 196.000 52.680 ;
        RECT 4.400 51.360 196.000 52.040 ;
        RECT 4.400 50.640 195.600 51.360 ;
        RECT 4.000 50.000 195.600 50.640 ;
        RECT 4.400 49.960 195.600 50.000 ;
        RECT 4.400 48.600 196.000 49.960 ;
        RECT 4.000 47.960 196.000 48.600 ;
        RECT 4.000 47.280 195.600 47.960 ;
        RECT 4.400 46.560 195.600 47.280 ;
        RECT 4.400 45.880 196.000 46.560 ;
        RECT 4.000 45.240 196.000 45.880 ;
        RECT 4.400 43.880 196.000 45.240 ;
        RECT 4.400 43.840 195.600 43.880 ;
        RECT 4.000 43.200 195.600 43.840 ;
        RECT 4.400 42.480 195.600 43.200 ;
        RECT 4.400 41.800 196.000 42.480 ;
        RECT 4.000 41.160 196.000 41.800 ;
        RECT 4.400 40.480 196.000 41.160 ;
        RECT 4.400 39.760 195.600 40.480 ;
        RECT 4.000 39.080 195.600 39.760 ;
        RECT 4.000 38.440 196.000 39.080 ;
        RECT 4.400 37.080 196.000 38.440 ;
        RECT 4.400 37.040 195.600 37.080 ;
        RECT 4.000 36.400 195.600 37.040 ;
        RECT 4.400 35.680 195.600 36.400 ;
        RECT 4.400 35.000 196.000 35.680 ;
        RECT 4.000 34.360 196.000 35.000 ;
        RECT 4.400 33.680 196.000 34.360 ;
        RECT 4.400 32.960 195.600 33.680 ;
        RECT 4.000 32.320 195.600 32.960 ;
        RECT 4.400 32.280 195.600 32.320 ;
        RECT 4.400 30.920 196.000 32.280 ;
        RECT 4.000 30.280 196.000 30.920 ;
        RECT 4.400 28.880 195.600 30.280 ;
        RECT 4.000 27.560 196.000 28.880 ;
        RECT 4.400 26.880 196.000 27.560 ;
        RECT 4.400 26.160 195.600 26.880 ;
        RECT 4.000 25.520 195.600 26.160 ;
        RECT 4.400 25.480 195.600 25.520 ;
        RECT 4.400 24.120 196.000 25.480 ;
        RECT 4.000 23.480 196.000 24.120 ;
        RECT 4.400 22.800 196.000 23.480 ;
        RECT 4.400 22.080 195.600 22.800 ;
        RECT 4.000 21.440 195.600 22.080 ;
        RECT 4.400 21.400 195.600 21.440 ;
        RECT 4.400 20.040 196.000 21.400 ;
        RECT 4.000 19.400 196.000 20.040 ;
        RECT 4.000 18.720 195.600 19.400 ;
        RECT 4.400 18.000 195.600 18.720 ;
        RECT 4.400 17.320 196.000 18.000 ;
        RECT 4.000 16.680 196.000 17.320 ;
        RECT 4.400 16.000 196.000 16.680 ;
        RECT 4.400 15.280 195.600 16.000 ;
        RECT 4.000 14.640 195.600 15.280 ;
        RECT 4.400 14.600 195.600 14.640 ;
        RECT 4.400 13.240 196.000 14.600 ;
        RECT 4.000 12.600 196.000 13.240 ;
        RECT 4.400 11.200 195.600 12.600 ;
        RECT 4.000 9.880 196.000 11.200 ;
        RECT 4.400 9.200 196.000 9.880 ;
        RECT 4.400 8.480 195.600 9.200 ;
        RECT 4.000 7.840 195.600 8.480 ;
        RECT 4.400 7.800 195.600 7.840 ;
        RECT 4.400 6.440 196.000 7.800 ;
        RECT 4.000 5.800 196.000 6.440 ;
        RECT 4.400 4.400 195.600 5.800 ;
        RECT 4.000 3.760 196.000 4.400 ;
        RECT 4.400 2.400 196.000 3.760 ;
        RECT 4.400 2.360 195.600 2.400 ;
        RECT 4.000 1.720 195.600 2.360 ;
        RECT 4.400 1.000 195.600 1.720 ;
        RECT 4.400 0.855 196.000 1.000 ;
  END
END GPIO
END LIBRARY

