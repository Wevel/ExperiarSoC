magic
tech sky130A
magscale 1 2
timestamp 1654558847
<< obsli1 >>
rect 1104 2159 118864 187697
<< obsm1 >>
rect 842 1436 119126 187808
<< metal2 >>
rect 754 189200 810 190000
rect 2318 189200 2374 190000
rect 3882 189200 3938 190000
rect 5446 189200 5502 190000
rect 7010 189200 7066 190000
rect 8574 189200 8630 190000
rect 10138 189200 10194 190000
rect 11794 189200 11850 190000
rect 13358 189200 13414 190000
rect 14922 189200 14978 190000
rect 16486 189200 16542 190000
rect 18050 189200 18106 190000
rect 19614 189200 19670 190000
rect 21270 189200 21326 190000
rect 22834 189200 22890 190000
rect 24398 189200 24454 190000
rect 25962 189200 26018 190000
rect 27526 189200 27582 190000
rect 29090 189200 29146 190000
rect 30746 189200 30802 190000
rect 32310 189200 32366 190000
rect 33874 189200 33930 190000
rect 35438 189200 35494 190000
rect 37002 189200 37058 190000
rect 38566 189200 38622 190000
rect 40130 189200 40186 190000
rect 41786 189200 41842 190000
rect 43350 189200 43406 190000
rect 44914 189200 44970 190000
rect 46478 189200 46534 190000
rect 48042 189200 48098 190000
rect 49606 189200 49662 190000
rect 51262 189200 51318 190000
rect 52826 189200 52882 190000
rect 54390 189200 54446 190000
rect 55954 189200 56010 190000
rect 57518 189200 57574 190000
rect 59082 189200 59138 190000
rect 60738 189200 60794 190000
rect 62302 189200 62358 190000
rect 63866 189200 63922 190000
rect 65430 189200 65486 190000
rect 66994 189200 67050 190000
rect 68558 189200 68614 190000
rect 70122 189200 70178 190000
rect 71778 189200 71834 190000
rect 73342 189200 73398 190000
rect 74906 189200 74962 190000
rect 76470 189200 76526 190000
rect 78034 189200 78090 190000
rect 79598 189200 79654 190000
rect 81254 189200 81310 190000
rect 82818 189200 82874 190000
rect 84382 189200 84438 190000
rect 85946 189200 86002 190000
rect 87510 189200 87566 190000
rect 89074 189200 89130 190000
rect 90730 189200 90786 190000
rect 92294 189200 92350 190000
rect 93858 189200 93914 190000
rect 95422 189200 95478 190000
rect 96986 189200 97042 190000
rect 98550 189200 98606 190000
rect 100114 189200 100170 190000
rect 101770 189200 101826 190000
rect 103334 189200 103390 190000
rect 104898 189200 104954 190000
rect 106462 189200 106518 190000
rect 108026 189200 108082 190000
rect 109590 189200 109646 190000
rect 111246 189200 111302 190000
rect 112810 189200 112866 190000
rect 114374 189200 114430 190000
rect 115938 189200 115994 190000
rect 117502 189200 117558 190000
rect 119066 189200 119122 190000
rect 846 0 902 800
rect 2594 0 2650 800
rect 4434 0 4490 800
rect 6274 0 6330 800
rect 8114 0 8170 800
rect 9862 0 9918 800
rect 11702 0 11758 800
rect 13542 0 13598 800
rect 15382 0 15438 800
rect 17130 0 17186 800
rect 18970 0 19026 800
rect 20810 0 20866 800
rect 22650 0 22706 800
rect 24398 0 24454 800
rect 26238 0 26294 800
rect 28078 0 28134 800
rect 29918 0 29974 800
rect 31666 0 31722 800
rect 33506 0 33562 800
rect 35346 0 35402 800
rect 37186 0 37242 800
rect 38934 0 38990 800
rect 40774 0 40830 800
rect 42614 0 42670 800
rect 44454 0 44510 800
rect 46202 0 46258 800
rect 48042 0 48098 800
rect 49882 0 49938 800
rect 51722 0 51778 800
rect 53470 0 53526 800
rect 55310 0 55366 800
rect 57150 0 57206 800
rect 58990 0 59046 800
rect 60830 0 60886 800
rect 62578 0 62634 800
rect 64418 0 64474 800
rect 66258 0 66314 800
rect 68098 0 68154 800
rect 69846 0 69902 800
rect 71686 0 71742 800
rect 73526 0 73582 800
rect 75366 0 75422 800
rect 77114 0 77170 800
rect 78954 0 79010 800
rect 80794 0 80850 800
rect 82634 0 82690 800
rect 84382 0 84438 800
rect 86222 0 86278 800
rect 88062 0 88118 800
rect 89902 0 89958 800
rect 91650 0 91706 800
rect 93490 0 93546 800
rect 95330 0 95386 800
rect 97170 0 97226 800
rect 98918 0 98974 800
rect 100758 0 100814 800
rect 102598 0 102654 800
rect 104438 0 104494 800
rect 106186 0 106242 800
rect 108026 0 108082 800
rect 109866 0 109922 800
rect 111706 0 111762 800
rect 113454 0 113510 800
rect 115294 0 115350 800
rect 117134 0 117190 800
rect 118974 0 119030 800
<< obsm2 >>
rect 866 189144 2262 189258
rect 2430 189144 3826 189258
rect 3994 189144 5390 189258
rect 5558 189144 6954 189258
rect 7122 189144 8518 189258
rect 8686 189144 10082 189258
rect 10250 189144 11738 189258
rect 11906 189144 13302 189258
rect 13470 189144 14866 189258
rect 15034 189144 16430 189258
rect 16598 189144 17994 189258
rect 18162 189144 19558 189258
rect 19726 189144 21214 189258
rect 21382 189144 22778 189258
rect 22946 189144 24342 189258
rect 24510 189144 25906 189258
rect 26074 189144 27470 189258
rect 27638 189144 29034 189258
rect 29202 189144 30690 189258
rect 30858 189144 32254 189258
rect 32422 189144 33818 189258
rect 33986 189144 35382 189258
rect 35550 189144 36946 189258
rect 37114 189144 38510 189258
rect 38678 189144 40074 189258
rect 40242 189144 41730 189258
rect 41898 189144 43294 189258
rect 43462 189144 44858 189258
rect 45026 189144 46422 189258
rect 46590 189144 47986 189258
rect 48154 189144 49550 189258
rect 49718 189144 51206 189258
rect 51374 189144 52770 189258
rect 52938 189144 54334 189258
rect 54502 189144 55898 189258
rect 56066 189144 57462 189258
rect 57630 189144 59026 189258
rect 59194 189144 60682 189258
rect 60850 189144 62246 189258
rect 62414 189144 63810 189258
rect 63978 189144 65374 189258
rect 65542 189144 66938 189258
rect 67106 189144 68502 189258
rect 68670 189144 70066 189258
rect 70234 189144 71722 189258
rect 71890 189144 73286 189258
rect 73454 189144 74850 189258
rect 75018 189144 76414 189258
rect 76582 189144 77978 189258
rect 78146 189144 79542 189258
rect 79710 189144 81198 189258
rect 81366 189144 82762 189258
rect 82930 189144 84326 189258
rect 84494 189144 85890 189258
rect 86058 189144 87454 189258
rect 87622 189144 89018 189258
rect 89186 189144 90674 189258
rect 90842 189144 92238 189258
rect 92406 189144 93802 189258
rect 93970 189144 95366 189258
rect 95534 189144 96930 189258
rect 97098 189144 98494 189258
rect 98662 189144 100058 189258
rect 100226 189144 101714 189258
rect 101882 189144 103278 189258
rect 103446 189144 104842 189258
rect 105010 189144 106406 189258
rect 106574 189144 107970 189258
rect 108138 189144 109534 189258
rect 109702 189144 111190 189258
rect 111358 189144 112754 189258
rect 112922 189144 114318 189258
rect 114486 189144 115882 189258
rect 116050 189144 117446 189258
rect 117614 189144 119010 189258
rect 848 856 119120 189144
rect 958 734 2538 856
rect 2706 734 4378 856
rect 4546 734 6218 856
rect 6386 734 8058 856
rect 8226 734 9806 856
rect 9974 734 11646 856
rect 11814 734 13486 856
rect 13654 734 15326 856
rect 15494 734 17074 856
rect 17242 734 18914 856
rect 19082 734 20754 856
rect 20922 734 22594 856
rect 22762 734 24342 856
rect 24510 734 26182 856
rect 26350 734 28022 856
rect 28190 734 29862 856
rect 30030 734 31610 856
rect 31778 734 33450 856
rect 33618 734 35290 856
rect 35458 734 37130 856
rect 37298 734 38878 856
rect 39046 734 40718 856
rect 40886 734 42558 856
rect 42726 734 44398 856
rect 44566 734 46146 856
rect 46314 734 47986 856
rect 48154 734 49826 856
rect 49994 734 51666 856
rect 51834 734 53414 856
rect 53582 734 55254 856
rect 55422 734 57094 856
rect 57262 734 58934 856
rect 59102 734 60774 856
rect 60942 734 62522 856
rect 62690 734 64362 856
rect 64530 734 66202 856
rect 66370 734 68042 856
rect 68210 734 69790 856
rect 69958 734 71630 856
rect 71798 734 73470 856
rect 73638 734 75310 856
rect 75478 734 77058 856
rect 77226 734 78898 856
rect 79066 734 80738 856
rect 80906 734 82578 856
rect 82746 734 84326 856
rect 84494 734 86166 856
rect 86334 734 88006 856
rect 88174 734 89846 856
rect 90014 734 91594 856
rect 91762 734 93434 856
rect 93602 734 95274 856
rect 95442 734 97114 856
rect 97282 734 98862 856
rect 99030 734 100702 856
rect 100870 734 102542 856
rect 102710 734 104382 856
rect 104550 734 106130 856
rect 106298 734 107970 856
rect 108138 734 109810 856
rect 109978 734 111650 856
rect 111818 734 113398 856
rect 113566 734 115238 856
rect 115406 734 117078 856
rect 117246 734 118918 856
rect 119086 734 119120 856
<< metal3 >>
rect 0 188912 800 189032
rect 0 187008 800 187128
rect 0 185104 800 185224
rect 0 183200 800 183320
rect 0 181296 800 181416
rect 0 179392 800 179512
rect 0 177488 800 177608
rect 0 175584 800 175704
rect 119200 174088 120000 174208
rect 0 173680 800 173800
rect 0 171776 800 171896
rect 0 169872 800 169992
rect 0 167968 800 168088
rect 0 166064 800 166184
rect 0 164160 800 164280
rect 0 162256 800 162376
rect 0 160352 800 160472
rect 0 158448 800 158568
rect 0 156544 800 156664
rect 0 154640 800 154760
rect 0 152736 800 152856
rect 0 150832 800 150952
rect 0 148928 800 149048
rect 0 147024 800 147144
rect 0 145120 800 145240
rect 0 143216 800 143336
rect 119200 142400 120000 142520
rect 0 141312 800 141432
rect 0 139408 800 139528
rect 0 137504 800 137624
rect 0 135600 800 135720
rect 0 133696 800 133816
rect 0 131792 800 131912
rect 0 129888 800 130008
rect 0 127984 800 128104
rect 0 126216 800 126336
rect 0 124312 800 124432
rect 0 122408 800 122528
rect 0 120504 800 120624
rect 0 118600 800 118720
rect 0 116696 800 116816
rect 0 114792 800 114912
rect 0 112888 800 113008
rect 0 110984 800 111104
rect 119200 110712 120000 110832
rect 0 109080 800 109200
rect 0 107176 800 107296
rect 0 105272 800 105392
rect 0 103368 800 103488
rect 0 101464 800 101584
rect 0 99560 800 99680
rect 0 97656 800 97776
rect 0 95752 800 95872
rect 0 93848 800 93968
rect 0 91944 800 92064
rect 0 90040 800 90160
rect 0 88136 800 88256
rect 0 86232 800 86352
rect 0 84328 800 84448
rect 0 82424 800 82544
rect 0 80520 800 80640
rect 119200 79024 120000 79144
rect 0 78616 800 78736
rect 0 76712 800 76832
rect 0 74808 800 74928
rect 0 72904 800 73024
rect 0 71000 800 71120
rect 0 69096 800 69216
rect 0 67192 800 67312
rect 0 65288 800 65408
rect 0 63520 800 63640
rect 0 61616 800 61736
rect 0 59712 800 59832
rect 0 57808 800 57928
rect 0 55904 800 56024
rect 0 54000 800 54120
rect 0 52096 800 52216
rect 0 50192 800 50312
rect 0 48288 800 48408
rect 119200 47336 120000 47456
rect 0 46384 800 46504
rect 0 44480 800 44600
rect 0 42576 800 42696
rect 0 40672 800 40792
rect 0 38768 800 38888
rect 0 36864 800 36984
rect 0 34960 800 35080
rect 0 33056 800 33176
rect 0 31152 800 31272
rect 0 29248 800 29368
rect 0 27344 800 27464
rect 0 25440 800 25560
rect 0 23536 800 23656
rect 0 21632 800 21752
rect 0 19728 800 19848
rect 0 17824 800 17944
rect 0 15920 800 16040
rect 119200 15784 120000 15904
rect 0 14016 800 14136
rect 0 12112 800 12232
rect 0 10208 800 10328
rect 0 8304 800 8424
rect 0 6400 800 6520
rect 0 4496 800 4616
rect 0 2592 800 2712
rect 0 824 800 944
<< obsm3 >>
rect 880 188832 119200 189005
rect 800 187208 119200 188832
rect 880 186928 119200 187208
rect 800 185304 119200 186928
rect 880 185024 119200 185304
rect 800 183400 119200 185024
rect 880 183120 119200 183400
rect 800 181496 119200 183120
rect 880 181216 119200 181496
rect 800 179592 119200 181216
rect 880 179312 119200 179592
rect 800 177688 119200 179312
rect 880 177408 119200 177688
rect 800 175784 119200 177408
rect 880 175504 119200 175784
rect 800 174288 119200 175504
rect 800 174008 119120 174288
rect 800 173880 119200 174008
rect 880 173600 119200 173880
rect 800 171976 119200 173600
rect 880 171696 119200 171976
rect 800 170072 119200 171696
rect 880 169792 119200 170072
rect 800 168168 119200 169792
rect 880 167888 119200 168168
rect 800 166264 119200 167888
rect 880 165984 119200 166264
rect 800 164360 119200 165984
rect 880 164080 119200 164360
rect 800 162456 119200 164080
rect 880 162176 119200 162456
rect 800 160552 119200 162176
rect 880 160272 119200 160552
rect 800 158648 119200 160272
rect 880 158368 119200 158648
rect 800 156744 119200 158368
rect 880 156464 119200 156744
rect 800 154840 119200 156464
rect 880 154560 119200 154840
rect 800 152936 119200 154560
rect 880 152656 119200 152936
rect 800 151032 119200 152656
rect 880 150752 119200 151032
rect 800 149128 119200 150752
rect 880 148848 119200 149128
rect 800 147224 119200 148848
rect 880 146944 119200 147224
rect 800 145320 119200 146944
rect 880 145040 119200 145320
rect 800 143416 119200 145040
rect 880 143136 119200 143416
rect 800 142600 119200 143136
rect 800 142320 119120 142600
rect 800 141512 119200 142320
rect 880 141232 119200 141512
rect 800 139608 119200 141232
rect 880 139328 119200 139608
rect 800 137704 119200 139328
rect 880 137424 119200 137704
rect 800 135800 119200 137424
rect 880 135520 119200 135800
rect 800 133896 119200 135520
rect 880 133616 119200 133896
rect 800 131992 119200 133616
rect 880 131712 119200 131992
rect 800 130088 119200 131712
rect 880 129808 119200 130088
rect 800 128184 119200 129808
rect 880 127904 119200 128184
rect 800 126416 119200 127904
rect 880 126136 119200 126416
rect 800 124512 119200 126136
rect 880 124232 119200 124512
rect 800 122608 119200 124232
rect 880 122328 119200 122608
rect 800 120704 119200 122328
rect 880 120424 119200 120704
rect 800 118800 119200 120424
rect 880 118520 119200 118800
rect 800 116896 119200 118520
rect 880 116616 119200 116896
rect 800 114992 119200 116616
rect 880 114712 119200 114992
rect 800 113088 119200 114712
rect 880 112808 119200 113088
rect 800 111184 119200 112808
rect 880 110912 119200 111184
rect 880 110904 119120 110912
rect 800 110632 119120 110904
rect 800 109280 119200 110632
rect 880 109000 119200 109280
rect 800 107376 119200 109000
rect 880 107096 119200 107376
rect 800 105472 119200 107096
rect 880 105192 119200 105472
rect 800 103568 119200 105192
rect 880 103288 119200 103568
rect 800 101664 119200 103288
rect 880 101384 119200 101664
rect 800 99760 119200 101384
rect 880 99480 119200 99760
rect 800 97856 119200 99480
rect 880 97576 119200 97856
rect 800 95952 119200 97576
rect 880 95672 119200 95952
rect 800 94048 119200 95672
rect 880 93768 119200 94048
rect 800 92144 119200 93768
rect 880 91864 119200 92144
rect 800 90240 119200 91864
rect 880 89960 119200 90240
rect 800 88336 119200 89960
rect 880 88056 119200 88336
rect 800 86432 119200 88056
rect 880 86152 119200 86432
rect 800 84528 119200 86152
rect 880 84248 119200 84528
rect 800 82624 119200 84248
rect 880 82344 119200 82624
rect 800 80720 119200 82344
rect 880 80440 119200 80720
rect 800 79224 119200 80440
rect 800 78944 119120 79224
rect 800 78816 119200 78944
rect 880 78536 119200 78816
rect 800 76912 119200 78536
rect 880 76632 119200 76912
rect 800 75008 119200 76632
rect 880 74728 119200 75008
rect 800 73104 119200 74728
rect 880 72824 119200 73104
rect 800 71200 119200 72824
rect 880 70920 119200 71200
rect 800 69296 119200 70920
rect 880 69016 119200 69296
rect 800 67392 119200 69016
rect 880 67112 119200 67392
rect 800 65488 119200 67112
rect 880 65208 119200 65488
rect 800 63720 119200 65208
rect 880 63440 119200 63720
rect 800 61816 119200 63440
rect 880 61536 119200 61816
rect 800 59912 119200 61536
rect 880 59632 119200 59912
rect 800 58008 119200 59632
rect 880 57728 119200 58008
rect 800 56104 119200 57728
rect 880 55824 119200 56104
rect 800 54200 119200 55824
rect 880 53920 119200 54200
rect 800 52296 119200 53920
rect 880 52016 119200 52296
rect 800 50392 119200 52016
rect 880 50112 119200 50392
rect 800 48488 119200 50112
rect 880 48208 119200 48488
rect 800 47536 119200 48208
rect 800 47256 119120 47536
rect 800 46584 119200 47256
rect 880 46304 119200 46584
rect 800 44680 119200 46304
rect 880 44400 119200 44680
rect 800 42776 119200 44400
rect 880 42496 119200 42776
rect 800 40872 119200 42496
rect 880 40592 119200 40872
rect 800 38968 119200 40592
rect 880 38688 119200 38968
rect 800 37064 119200 38688
rect 880 36784 119200 37064
rect 800 35160 119200 36784
rect 880 34880 119200 35160
rect 800 33256 119200 34880
rect 880 32976 119200 33256
rect 800 31352 119200 32976
rect 880 31072 119200 31352
rect 800 29448 119200 31072
rect 880 29168 119200 29448
rect 800 27544 119200 29168
rect 880 27264 119200 27544
rect 800 25640 119200 27264
rect 880 25360 119200 25640
rect 800 23736 119200 25360
rect 880 23456 119200 23736
rect 800 21832 119200 23456
rect 880 21552 119200 21832
rect 800 19928 119200 21552
rect 880 19648 119200 19928
rect 800 18024 119200 19648
rect 880 17744 119200 18024
rect 800 16120 119200 17744
rect 880 15984 119200 16120
rect 880 15840 119120 15984
rect 800 15704 119120 15840
rect 800 14216 119200 15704
rect 880 13936 119200 14216
rect 800 12312 119200 13936
rect 880 12032 119200 12312
rect 800 10408 119200 12032
rect 880 10128 119200 10408
rect 800 8504 119200 10128
rect 880 8224 119200 8504
rect 800 6600 119200 8224
rect 880 6320 119200 6600
rect 800 4696 119200 6320
rect 880 4416 119200 4696
rect 800 2792 119200 4416
rect 880 2512 119200 2792
rect 800 1024 119200 2512
rect 880 851 119200 1024
<< metal4 >>
rect 4208 2128 4528 187728
rect 19568 2128 19888 187728
rect 34928 2128 35248 187728
rect 50288 2128 50608 187728
rect 65648 2128 65968 187728
rect 81008 2128 81328 187728
rect 96368 2128 96688 187728
rect 111728 2128 112048 187728
<< obsm4 >>
rect 1715 2619 4128 186693
rect 4608 2619 19488 186693
rect 19968 2619 34848 186693
rect 35328 2619 50208 186693
rect 50688 2619 65568 186693
rect 66048 2619 80928 186693
rect 81408 2619 96288 186693
rect 96768 2619 111648 186693
rect 112128 2619 116045 186693
<< labels >>
rlabel metal2 s 73526 0 73582 800 6 flash_csb
port 1 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 flash_io0_read
port 2 nsew signal output
rlabel metal2 s 77114 0 77170 800 6 flash_io0_we
port 3 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 flash_io0_write
port 4 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 flash_io1_read
port 5 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 flash_io1_we
port 6 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 flash_io1_write
port 7 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 flash_sck
port 8 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 internal_uart_rx
port 9 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 internal_uart_tx
port 10 nsew signal output
rlabel metal2 s 754 189200 810 190000 6 io_in[0]
port 11 nsew signal input
rlabel metal2 s 16486 189200 16542 190000 6 io_in[10]
port 12 nsew signal input
rlabel metal2 s 18050 189200 18106 190000 6 io_in[11]
port 13 nsew signal input
rlabel metal2 s 19614 189200 19670 190000 6 io_in[12]
port 14 nsew signal input
rlabel metal2 s 21270 189200 21326 190000 6 io_in[13]
port 15 nsew signal input
rlabel metal2 s 22834 189200 22890 190000 6 io_in[14]
port 16 nsew signal input
rlabel metal2 s 24398 189200 24454 190000 6 io_in[15]
port 17 nsew signal input
rlabel metal2 s 25962 189200 26018 190000 6 io_in[16]
port 18 nsew signal input
rlabel metal2 s 27526 189200 27582 190000 6 io_in[17]
port 19 nsew signal input
rlabel metal2 s 29090 189200 29146 190000 6 io_in[18]
port 20 nsew signal input
rlabel metal2 s 30746 189200 30802 190000 6 io_in[19]
port 21 nsew signal input
rlabel metal2 s 2318 189200 2374 190000 6 io_in[1]
port 22 nsew signal input
rlabel metal2 s 32310 189200 32366 190000 6 io_in[20]
port 23 nsew signal input
rlabel metal2 s 33874 189200 33930 190000 6 io_in[21]
port 24 nsew signal input
rlabel metal2 s 35438 189200 35494 190000 6 io_in[22]
port 25 nsew signal input
rlabel metal2 s 37002 189200 37058 190000 6 io_in[23]
port 26 nsew signal input
rlabel metal2 s 38566 189200 38622 190000 6 io_in[24]
port 27 nsew signal input
rlabel metal2 s 40130 189200 40186 190000 6 io_in[25]
port 28 nsew signal input
rlabel metal2 s 41786 189200 41842 190000 6 io_in[26]
port 29 nsew signal input
rlabel metal2 s 43350 189200 43406 190000 6 io_in[27]
port 30 nsew signal input
rlabel metal2 s 44914 189200 44970 190000 6 io_in[28]
port 31 nsew signal input
rlabel metal2 s 46478 189200 46534 190000 6 io_in[29]
port 32 nsew signal input
rlabel metal2 s 3882 189200 3938 190000 6 io_in[2]
port 33 nsew signal input
rlabel metal2 s 48042 189200 48098 190000 6 io_in[30]
port 34 nsew signal input
rlabel metal2 s 49606 189200 49662 190000 6 io_in[31]
port 35 nsew signal input
rlabel metal2 s 51262 189200 51318 190000 6 io_in[32]
port 36 nsew signal input
rlabel metal2 s 52826 189200 52882 190000 6 io_in[33]
port 37 nsew signal input
rlabel metal2 s 54390 189200 54446 190000 6 io_in[34]
port 38 nsew signal input
rlabel metal2 s 55954 189200 56010 190000 6 io_in[35]
port 39 nsew signal input
rlabel metal2 s 57518 189200 57574 190000 6 io_in[36]
port 40 nsew signal input
rlabel metal2 s 59082 189200 59138 190000 6 io_in[37]
port 41 nsew signal input
rlabel metal2 s 5446 189200 5502 190000 6 io_in[3]
port 42 nsew signal input
rlabel metal2 s 7010 189200 7066 190000 6 io_in[4]
port 43 nsew signal input
rlabel metal2 s 8574 189200 8630 190000 6 io_in[5]
port 44 nsew signal input
rlabel metal2 s 10138 189200 10194 190000 6 io_in[6]
port 45 nsew signal input
rlabel metal2 s 11794 189200 11850 190000 6 io_in[7]
port 46 nsew signal input
rlabel metal2 s 13358 189200 13414 190000 6 io_in[8]
port 47 nsew signal input
rlabel metal2 s 14922 189200 14978 190000 6 io_in[9]
port 48 nsew signal input
rlabel metal2 s 846 0 902 800 6 io_oeb[0]
port 49 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 io_oeb[10]
port 50 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 io_oeb[11]
port 51 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 io_oeb[12]
port 52 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 io_oeb[13]
port 53 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 io_oeb[14]
port 54 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 io_oeb[15]
port 55 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 io_oeb[16]
port 56 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 io_oeb[17]
port 57 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 io_oeb[18]
port 58 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 io_oeb[19]
port 59 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 io_oeb[1]
port 60 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 io_oeb[20]
port 61 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 io_oeb[21]
port 62 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 io_oeb[22]
port 63 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 io_oeb[23]
port 64 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 io_oeb[24]
port 65 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 io_oeb[25]
port 66 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 io_oeb[26]
port 67 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 io_oeb[27]
port 68 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 io_oeb[28]
port 69 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 io_oeb[29]
port 70 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 io_oeb[2]
port 71 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 io_oeb[30]
port 72 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 io_oeb[31]
port 73 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 io_oeb[32]
port 74 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 io_oeb[33]
port 75 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 io_oeb[34]
port 76 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 io_oeb[35]
port 77 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 io_oeb[36]
port 78 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 io_oeb[37]
port 79 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 io_oeb[3]
port 80 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 io_oeb[4]
port 81 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 io_oeb[5]
port 82 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 io_oeb[6]
port 83 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 io_oeb[7]
port 84 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 io_oeb[8]
port 85 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 60738 189200 60794 190000 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 76470 189200 76526 190000 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 78034 189200 78090 190000 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 79598 189200 79654 190000 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 81254 189200 81310 190000 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 82818 189200 82874 190000 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 84382 189200 84438 190000 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 85946 189200 86002 190000 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 87510 189200 87566 190000 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 89074 189200 89130 190000 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 90730 189200 90786 190000 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 62302 189200 62358 190000 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 92294 189200 92350 190000 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 93858 189200 93914 190000 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 95422 189200 95478 190000 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 96986 189200 97042 190000 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 98550 189200 98606 190000 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 100114 189200 100170 190000 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 101770 189200 101826 190000 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 103334 189200 103390 190000 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 104898 189200 104954 190000 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 106462 189200 106518 190000 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 63866 189200 63922 190000 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 108026 189200 108082 190000 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 109590 189200 109646 190000 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 111246 189200 111302 190000 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 112810 189200 112866 190000 6 io_out[33]
port 113 nsew signal output
rlabel metal2 s 114374 189200 114430 190000 6 io_out[34]
port 114 nsew signal output
rlabel metal2 s 115938 189200 115994 190000 6 io_out[35]
port 115 nsew signal output
rlabel metal2 s 117502 189200 117558 190000 6 io_out[36]
port 116 nsew signal output
rlabel metal2 s 119066 189200 119122 190000 6 io_out[37]
port 117 nsew signal output
rlabel metal2 s 65430 189200 65486 190000 6 io_out[3]
port 118 nsew signal output
rlabel metal2 s 66994 189200 67050 190000 6 io_out[4]
port 119 nsew signal output
rlabel metal2 s 68558 189200 68614 190000 6 io_out[5]
port 120 nsew signal output
rlabel metal2 s 70122 189200 70178 190000 6 io_out[6]
port 121 nsew signal output
rlabel metal2 s 71778 189200 71834 190000 6 io_out[7]
port 122 nsew signal output
rlabel metal2 s 73342 189200 73398 190000 6 io_out[8]
port 123 nsew signal output
rlabel metal2 s 74906 189200 74962 190000 6 io_out[9]
port 124 nsew signal output
rlabel metal3 s 119200 79024 120000 79144 6 jtag_tck
port 125 nsew signal output
rlabel metal3 s 119200 110712 120000 110832 6 jtag_tdi
port 126 nsew signal output
rlabel metal3 s 119200 142400 120000 142520 6 jtag_tdo
port 127 nsew signal input
rlabel metal3 s 119200 174088 120000 174208 6 jtag_tms
port 128 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 peripheral_irq[0]
port 129 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 peripheral_irq[1]
port 130 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 peripheral_irq[2]
port 131 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 peripheral_irq[3]
port 132 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 peripheral_irq[4]
port 133 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 peripheral_irq[5]
port 134 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 peripheral_irq[6]
port 135 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 peripheral_irq[7]
port 136 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 peripheral_irq[8]
port 137 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 peripheral_irq[9]
port 138 nsew signal output
rlabel metal3 s 119200 15784 120000 15904 6 probe_blink[0]
port 139 nsew signal output
rlabel metal3 s 119200 47336 120000 47456 6 probe_blink[1]
port 140 nsew signal output
rlabel metal4 s 4208 2128 4528 187728 6 vccd1
port 141 nsew power input
rlabel metal4 s 34928 2128 35248 187728 6 vccd1
port 141 nsew power input
rlabel metal4 s 65648 2128 65968 187728 6 vccd1
port 141 nsew power input
rlabel metal4 s 96368 2128 96688 187728 6 vccd1
port 141 nsew power input
rlabel metal2 s 109866 0 109922 800 6 vga_b[0]
port 142 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 vga_b[1]
port 143 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 vga_g[0]
port 144 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 vga_g[1]
port 145 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 vga_hsync
port 146 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 vga_r[0]
port 147 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 vga_r[1]
port 148 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 vga_vsync
port 149 nsew signal input
rlabel metal4 s 19568 2128 19888 187728 6 vssd1
port 150 nsew ground input
rlabel metal4 s 50288 2128 50608 187728 6 vssd1
port 150 nsew ground input
rlabel metal4 s 81008 2128 81328 187728 6 vssd1
port 150 nsew ground input
rlabel metal4 s 111728 2128 112048 187728 6 vssd1
port 150 nsew ground input
rlabel metal3 s 0 824 800 944 6 wb_ack_o
port 151 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 wb_adr_i[0]
port 152 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 wb_adr_i[10]
port 153 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 wb_adr_i[11]
port 154 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 wb_adr_i[12]
port 155 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 wb_adr_i[13]
port 156 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 wb_adr_i[14]
port 157 nsew signal input
rlabel metal3 s 0 109080 800 109200 6 wb_adr_i[15]
port 158 nsew signal input
rlabel metal3 s 0 114792 800 114912 6 wb_adr_i[16]
port 159 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 wb_adr_i[17]
port 160 nsew signal input
rlabel metal3 s 0 126216 800 126336 6 wb_adr_i[18]
port 161 nsew signal input
rlabel metal3 s 0 131792 800 131912 6 wb_adr_i[19]
port 162 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 wb_adr_i[1]
port 163 nsew signal input
rlabel metal3 s 0 137504 800 137624 6 wb_adr_i[20]
port 164 nsew signal input
rlabel metal3 s 0 143216 800 143336 6 wb_adr_i[21]
port 165 nsew signal input
rlabel metal3 s 0 148928 800 149048 6 wb_adr_i[22]
port 166 nsew signal input
rlabel metal3 s 0 154640 800 154760 6 wb_adr_i[23]
port 167 nsew signal input
rlabel metal3 s 0 31152 800 31272 6 wb_adr_i[2]
port 168 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 wb_adr_i[3]
port 169 nsew signal input
rlabel metal3 s 0 46384 800 46504 6 wb_adr_i[4]
port 170 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 wb_adr_i[5]
port 171 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 wb_adr_i[6]
port 172 nsew signal input
rlabel metal3 s 0 63520 800 63640 6 wb_adr_i[7]
port 173 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 wb_adr_i[8]
port 174 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 wb_adr_i[9]
port 175 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 wb_clk_i
port 176 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 wb_cyc_i
port 177 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 wb_data_i[0]
port 178 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 wb_data_i[10]
port 179 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 wb_data_i[11]
port 180 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 wb_data_i[12]
port 181 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 wb_data_i[13]
port 182 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 wb_data_i[14]
port 183 nsew signal input
rlabel metal3 s 0 110984 800 111104 6 wb_data_i[15]
port 184 nsew signal input
rlabel metal3 s 0 116696 800 116816 6 wb_data_i[16]
port 185 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 wb_data_i[17]
port 186 nsew signal input
rlabel metal3 s 0 127984 800 128104 6 wb_data_i[18]
port 187 nsew signal input
rlabel metal3 s 0 133696 800 133816 6 wb_data_i[19]
port 188 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 wb_data_i[1]
port 189 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 wb_data_i[20]
port 190 nsew signal input
rlabel metal3 s 0 145120 800 145240 6 wb_data_i[21]
port 191 nsew signal input
rlabel metal3 s 0 150832 800 150952 6 wb_data_i[22]
port 192 nsew signal input
rlabel metal3 s 0 156544 800 156664 6 wb_data_i[23]
port 193 nsew signal input
rlabel metal3 s 0 160352 800 160472 6 wb_data_i[24]
port 194 nsew signal input
rlabel metal3 s 0 164160 800 164280 6 wb_data_i[25]
port 195 nsew signal input
rlabel metal3 s 0 167968 800 168088 6 wb_data_i[26]
port 196 nsew signal input
rlabel metal3 s 0 171776 800 171896 6 wb_data_i[27]
port 197 nsew signal input
rlabel metal3 s 0 175584 800 175704 6 wb_data_i[28]
port 198 nsew signal input
rlabel metal3 s 0 179392 800 179512 6 wb_data_i[29]
port 199 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 wb_data_i[2]
port 200 nsew signal input
rlabel metal3 s 0 183200 800 183320 6 wb_data_i[30]
port 201 nsew signal input
rlabel metal3 s 0 187008 800 187128 6 wb_data_i[31]
port 202 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 wb_data_i[3]
port 203 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 wb_data_i[4]
port 204 nsew signal input
rlabel metal3 s 0 54000 800 54120 6 wb_data_i[5]
port 205 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 wb_data_i[6]
port 206 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 wb_data_i[7]
port 207 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 wb_data_i[8]
port 208 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 wb_data_i[9]
port 209 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 wb_data_o[0]
port 210 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 wb_data_o[10]
port 211 nsew signal output
rlabel metal3 s 0 90040 800 90160 6 wb_data_o[11]
port 212 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 wb_data_o[12]
port 213 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 wb_data_o[13]
port 214 nsew signal output
rlabel metal3 s 0 107176 800 107296 6 wb_data_o[14]
port 215 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 wb_data_o[15]
port 216 nsew signal output
rlabel metal3 s 0 118600 800 118720 6 wb_data_o[16]
port 217 nsew signal output
rlabel metal3 s 0 124312 800 124432 6 wb_data_o[17]
port 218 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 wb_data_o[18]
port 219 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 wb_data_o[19]
port 220 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 wb_data_o[1]
port 221 nsew signal output
rlabel metal3 s 0 141312 800 141432 6 wb_data_o[20]
port 222 nsew signal output
rlabel metal3 s 0 147024 800 147144 6 wb_data_o[21]
port 223 nsew signal output
rlabel metal3 s 0 152736 800 152856 6 wb_data_o[22]
port 224 nsew signal output
rlabel metal3 s 0 158448 800 158568 6 wb_data_o[23]
port 225 nsew signal output
rlabel metal3 s 0 162256 800 162376 6 wb_data_o[24]
port 226 nsew signal output
rlabel metal3 s 0 166064 800 166184 6 wb_data_o[25]
port 227 nsew signal output
rlabel metal3 s 0 169872 800 169992 6 wb_data_o[26]
port 228 nsew signal output
rlabel metal3 s 0 173680 800 173800 6 wb_data_o[27]
port 229 nsew signal output
rlabel metal3 s 0 177488 800 177608 6 wb_data_o[28]
port 230 nsew signal output
rlabel metal3 s 0 181296 800 181416 6 wb_data_o[29]
port 231 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 wb_data_o[2]
port 232 nsew signal output
rlabel metal3 s 0 185104 800 185224 6 wb_data_o[30]
port 233 nsew signal output
rlabel metal3 s 0 188912 800 189032 6 wb_data_o[31]
port 234 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 wb_data_o[3]
port 235 nsew signal output
rlabel metal3 s 0 50192 800 50312 6 wb_data_o[4]
port 236 nsew signal output
rlabel metal3 s 0 55904 800 56024 6 wb_data_o[5]
port 237 nsew signal output
rlabel metal3 s 0 61616 800 61736 6 wb_data_o[6]
port 238 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 wb_data_o[7]
port 239 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 wb_data_o[8]
port 240 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 wb_data_o[9]
port 241 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 wb_error_o
port 242 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 wb_rst_i
port 243 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 wb_sel_i[0]
port 244 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 wb_sel_i[1]
port 245 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 wb_sel_i[2]
port 246 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 wb_sel_i[3]
port 247 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 wb_stall_o
port 248 nsew signal output
rlabel metal3 s 0 12112 800 12232 6 wb_stb_i
port 249 nsew signal input
rlabel metal3 s 0 14016 800 14136 6 wb_we_i
port 250 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 190000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 69323354
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripherals_Flat/runs/Peripherals_Flat/results/finishing/Peripherals.magic.gds
string GDS_START 1312988
<< end >>

