VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ExperiarCore
  CLASS BLOCK ;
  FOREIGN ExperiarCore ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 800.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END addr0[8]
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.280 4.000 505.880 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 509.360 4.000 509.960 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 521.600 4.000 522.200 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.760 4.000 530.360 ;
    END
  END addr1[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END clk0
  PIN clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.880 4.000 485.480 ;
    END
  END clk1
  PIN coreIndex[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 796.000 14.170 800.000 ;
    END
  END coreIndex[0]
  PIN coreIndex[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 796.000 26.590 800.000 ;
    END
  END coreIndex[1]
  PIN coreIndex[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 796.000 39.010 800.000 ;
    END
  END coreIndex[2]
  PIN coreIndex[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 796.000 51.430 800.000 ;
    END
  END coreIndex[3]
  PIN coreIndex[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 796.000 63.850 800.000 ;
    END
  END coreIndex[4]
  PIN coreIndex[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 796.000 76.270 800.000 ;
    END
  END coreIndex[5]
  PIN coreIndex[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 796.000 88.690 800.000 ;
    END
  END coreIndex[6]
  PIN coreIndex[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 796.000 101.110 800.000 ;
    END
  END coreIndex[7]
  PIN core_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 64.640 500.000 65.240 ;
    END
  END core_wb_ack_i
  PIN core_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 85.040 500.000 85.640 ;
    END
  END core_wb_adr_o[0]
  PIN core_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 200.640 500.000 201.240 ;
    END
  END core_wb_adr_o[10]
  PIN core_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.840 500.000 211.440 ;
    END
  END core_wb_adr_o[11]
  PIN core_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 221.040 500.000 221.640 ;
    END
  END core_wb_adr_o[12]
  PIN core_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 231.240 500.000 231.840 ;
    END
  END core_wb_adr_o[13]
  PIN core_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 241.440 500.000 242.040 ;
    END
  END core_wb_adr_o[14]
  PIN core_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 251.640 500.000 252.240 ;
    END
  END core_wb_adr_o[15]
  PIN core_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 261.840 500.000 262.440 ;
    END
  END core_wb_adr_o[16]
  PIN core_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 272.040 500.000 272.640 ;
    END
  END core_wb_adr_o[17]
  PIN core_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 282.240 500.000 282.840 ;
    END
  END core_wb_adr_o[18]
  PIN core_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 292.440 500.000 293.040 ;
    END
  END core_wb_adr_o[19]
  PIN core_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 98.640 500.000 99.240 ;
    END
  END core_wb_adr_o[1]
  PIN core_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 302.640 500.000 303.240 ;
    END
  END core_wb_adr_o[20]
  PIN core_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 312.840 500.000 313.440 ;
    END
  END core_wb_adr_o[21]
  PIN core_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 323.040 500.000 323.640 ;
    END
  END core_wb_adr_o[22]
  PIN core_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 333.240 500.000 333.840 ;
    END
  END core_wb_adr_o[23]
  PIN core_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 343.440 500.000 344.040 ;
    END
  END core_wb_adr_o[24]
  PIN core_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 353.640 500.000 354.240 ;
    END
  END core_wb_adr_o[25]
  PIN core_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 363.840 500.000 364.440 ;
    END
  END core_wb_adr_o[26]
  PIN core_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 374.040 500.000 374.640 ;
    END
  END core_wb_adr_o[27]
  PIN core_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 112.240 500.000 112.840 ;
    END
  END core_wb_adr_o[2]
  PIN core_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 125.840 500.000 126.440 ;
    END
  END core_wb_adr_o[3]
  PIN core_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 139.440 500.000 140.040 ;
    END
  END core_wb_adr_o[4]
  PIN core_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 149.640 500.000 150.240 ;
    END
  END core_wb_adr_o[5]
  PIN core_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 159.840 500.000 160.440 ;
    END
  END core_wb_adr_o[6]
  PIN core_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 170.040 500.000 170.640 ;
    END
  END core_wb_adr_o[7]
  PIN core_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 180.240 500.000 180.840 ;
    END
  END core_wb_adr_o[8]
  PIN core_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 190.440 500.000 191.040 ;
    END
  END core_wb_adr_o[9]
  PIN core_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 68.040 500.000 68.640 ;
    END
  END core_wb_cyc_o
  PIN core_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 88.440 500.000 89.040 ;
    END
  END core_wb_data_i[0]
  PIN core_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 204.040 500.000 204.640 ;
    END
  END core_wb_data_i[10]
  PIN core_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 214.240 500.000 214.840 ;
    END
  END core_wb_data_i[11]
  PIN core_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 224.440 500.000 225.040 ;
    END
  END core_wb_data_i[12]
  PIN core_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 234.640 500.000 235.240 ;
    END
  END core_wb_data_i[13]
  PIN core_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 244.840 500.000 245.440 ;
    END
  END core_wb_data_i[14]
  PIN core_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 255.040 500.000 255.640 ;
    END
  END core_wb_data_i[15]
  PIN core_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 265.240 500.000 265.840 ;
    END
  END core_wb_data_i[16]
  PIN core_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 275.440 500.000 276.040 ;
    END
  END core_wb_data_i[17]
  PIN core_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 285.640 500.000 286.240 ;
    END
  END core_wb_data_i[18]
  PIN core_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 295.840 500.000 296.440 ;
    END
  END core_wb_data_i[19]
  PIN core_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 102.040 500.000 102.640 ;
    END
  END core_wb_data_i[1]
  PIN core_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 306.040 500.000 306.640 ;
    END
  END core_wb_data_i[20]
  PIN core_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 316.240 500.000 316.840 ;
    END
  END core_wb_data_i[21]
  PIN core_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 326.440 500.000 327.040 ;
    END
  END core_wb_data_i[22]
  PIN core_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 336.640 500.000 337.240 ;
    END
  END core_wb_data_i[23]
  PIN core_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 346.840 500.000 347.440 ;
    END
  END core_wb_data_i[24]
  PIN core_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 357.040 500.000 357.640 ;
    END
  END core_wb_data_i[25]
  PIN core_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 367.240 500.000 367.840 ;
    END
  END core_wb_data_i[26]
  PIN core_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 377.440 500.000 378.040 ;
    END
  END core_wb_data_i[27]
  PIN core_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 384.240 500.000 384.840 ;
    END
  END core_wb_data_i[28]
  PIN core_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 391.040 500.000 391.640 ;
    END
  END core_wb_data_i[29]
  PIN core_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 115.640 500.000 116.240 ;
    END
  END core_wb_data_i[2]
  PIN core_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 397.840 500.000 398.440 ;
    END
  END core_wb_data_i[30]
  PIN core_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 404.640 500.000 405.240 ;
    END
  END core_wb_data_i[31]
  PIN core_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 129.240 500.000 129.840 ;
    END
  END core_wb_data_i[3]
  PIN core_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 142.840 500.000 143.440 ;
    END
  END core_wb_data_i[4]
  PIN core_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 153.040 500.000 153.640 ;
    END
  END core_wb_data_i[5]
  PIN core_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 163.240 500.000 163.840 ;
    END
  END core_wb_data_i[6]
  PIN core_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 173.440 500.000 174.040 ;
    END
  END core_wb_data_i[7]
  PIN core_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 183.640 500.000 184.240 ;
    END
  END core_wb_data_i[8]
  PIN core_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 193.840 500.000 194.440 ;
    END
  END core_wb_data_i[9]
  PIN core_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 91.840 500.000 92.440 ;
    END
  END core_wb_data_o[0]
  PIN core_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 207.440 500.000 208.040 ;
    END
  END core_wb_data_o[10]
  PIN core_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 217.640 500.000 218.240 ;
    END
  END core_wb_data_o[11]
  PIN core_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 227.840 500.000 228.440 ;
    END
  END core_wb_data_o[12]
  PIN core_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 238.040 500.000 238.640 ;
    END
  END core_wb_data_o[13]
  PIN core_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 248.240 500.000 248.840 ;
    END
  END core_wb_data_o[14]
  PIN core_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 258.440 500.000 259.040 ;
    END
  END core_wb_data_o[15]
  PIN core_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 268.640 500.000 269.240 ;
    END
  END core_wb_data_o[16]
  PIN core_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 278.840 500.000 279.440 ;
    END
  END core_wb_data_o[17]
  PIN core_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 289.040 500.000 289.640 ;
    END
  END core_wb_data_o[18]
  PIN core_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 299.240 500.000 299.840 ;
    END
  END core_wb_data_o[19]
  PIN core_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 105.440 500.000 106.040 ;
    END
  END core_wb_data_o[1]
  PIN core_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 309.440 500.000 310.040 ;
    END
  END core_wb_data_o[20]
  PIN core_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 319.640 500.000 320.240 ;
    END
  END core_wb_data_o[21]
  PIN core_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 329.840 500.000 330.440 ;
    END
  END core_wb_data_o[22]
  PIN core_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.040 500.000 340.640 ;
    END
  END core_wb_data_o[23]
  PIN core_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 350.240 500.000 350.840 ;
    END
  END core_wb_data_o[24]
  PIN core_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 360.440 500.000 361.040 ;
    END
  END core_wb_data_o[25]
  PIN core_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 370.640 500.000 371.240 ;
    END
  END core_wb_data_o[26]
  PIN core_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 380.840 500.000 381.440 ;
    END
  END core_wb_data_o[27]
  PIN core_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 387.640 500.000 388.240 ;
    END
  END core_wb_data_o[28]
  PIN core_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 394.440 500.000 395.040 ;
    END
  END core_wb_data_o[29]
  PIN core_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 119.040 500.000 119.640 ;
    END
  END core_wb_data_o[2]
  PIN core_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 401.240 500.000 401.840 ;
    END
  END core_wb_data_o[30]
  PIN core_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 408.040 500.000 408.640 ;
    END
  END core_wb_data_o[31]
  PIN core_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 132.640 500.000 133.240 ;
    END
  END core_wb_data_o[3]
  PIN core_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 146.240 500.000 146.840 ;
    END
  END core_wb_data_o[4]
  PIN core_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 156.440 500.000 157.040 ;
    END
  END core_wb_data_o[5]
  PIN core_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 166.640 500.000 167.240 ;
    END
  END core_wb_data_o[6]
  PIN core_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 176.840 500.000 177.440 ;
    END
  END core_wb_data_o[7]
  PIN core_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 187.040 500.000 187.640 ;
    END
  END core_wb_data_o[8]
  PIN core_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 197.240 500.000 197.840 ;
    END
  END core_wb_data_o[9]
  PIN core_wb_error_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 71.440 500.000 72.040 ;
    END
  END core_wb_error_i
  PIN core_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.240 500.000 95.840 ;
    END
  END core_wb_sel_o[0]
  PIN core_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 108.840 500.000 109.440 ;
    END
  END core_wb_sel_o[1]
  PIN core_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 122.440 500.000 123.040 ;
    END
  END core_wb_sel_o[2]
  PIN core_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 136.040 500.000 136.640 ;
    END
  END core_wb_sel_o[3]
  PIN core_wb_stall_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 74.840 500.000 75.440 ;
    END
  END core_wb_stall_i
  PIN core_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 78.240 500.000 78.840 ;
    END
  END core_wb_stb_o
  PIN core_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 81.640 500.000 82.240 ;
    END
  END core_wb_we_o
  PIN csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END csb0[0]
  PIN csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END csb0[1]
  PIN csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END csb1[0]
  PIN csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END csb1[1]
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END din0[9]
  PIN dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END dout0[32]
  PIN dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END dout0[33]
  PIN dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END dout0[34]
  PIN dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END dout0[35]
  PIN dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END dout0[36]
  PIN dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END dout0[37]
  PIN dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END dout0[38]
  PIN dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END dout0[39]
  PIN dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END dout0[3]
  PIN dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END dout0[40]
  PIN dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END dout0[41]
  PIN dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END dout0[42]
  PIN dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END dout0[43]
  PIN dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END dout0[44]
  PIN dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END dout0[45]
  PIN dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END dout0[46]
  PIN dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END dout0[47]
  PIN dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.600 4.000 420.200 ;
    END
  END dout0[48]
  PIN dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END dout0[49]
  PIN dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END dout0[4]
  PIN dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END dout0[50]
  PIN dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END dout0[51]
  PIN dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END dout0[52]
  PIN dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END dout0[53]
  PIN dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END dout0[54]
  PIN dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.160 4.000 448.760 ;
    END
  END dout0[55]
  PIN dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END dout0[56]
  PIN dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 456.320 4.000 456.920 ;
    END
  END dout0[57]
  PIN dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 460.400 4.000 461.000 ;
    END
  END dout0[58]
  PIN dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 464.480 4.000 465.080 ;
    END
  END dout0[59]
  PIN dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END dout0[5]
  PIN dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END dout0[60]
  PIN dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END dout0[61]
  PIN dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END dout0[62]
  PIN dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END dout0[63]
  PIN dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END dout0[9]
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.800 4.000 583.400 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.880 4.000 587.480 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.280 4.000 607.880 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 611.360 4.000 611.960 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 4.000 538.520 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 619.520 4.000 620.120 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.000 4.000 644.600 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.080 4.000 648.680 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.000 4.000 542.600 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END dout1[31]
  PIN dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END dout1[32]
  PIN dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END dout1[33]
  PIN dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 672.560 4.000 673.160 ;
    END
  END dout1[34]
  PIN dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END dout1[35]
  PIN dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END dout1[36]
  PIN dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END dout1[37]
  PIN dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END dout1[38]
  PIN dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.960 4.000 693.560 ;
    END
  END dout1[39]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.080 4.000 546.680 ;
    END
  END dout1[3]
  PIN dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END dout1[40]
  PIN dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.120 4.000 701.720 ;
    END
  END dout1[41]
  PIN dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.200 4.000 705.800 ;
    END
  END dout1[42]
  PIN dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.280 4.000 709.880 ;
    END
  END dout1[43]
  PIN dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 713.360 4.000 713.960 ;
    END
  END dout1[44]
  PIN dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END dout1[45]
  PIN dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 721.520 4.000 722.120 ;
    END
  END dout1[46]
  PIN dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END dout1[47]
  PIN dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.680 4.000 730.280 ;
    END
  END dout1[48]
  PIN dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.760 4.000 734.360 ;
    END
  END dout1[49]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END dout1[4]
  PIN dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END dout1[50]
  PIN dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.920 4.000 742.520 ;
    END
  END dout1[51]
  PIN dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.000 4.000 746.600 ;
    END
  END dout1[52]
  PIN dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.080 4.000 750.680 ;
    END
  END dout1[53]
  PIN dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.160 4.000 754.760 ;
    END
  END dout1[54]
  PIN dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END dout1[55]
  PIN dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 762.320 4.000 762.920 ;
    END
  END dout1[56]
  PIN dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 766.400 4.000 767.000 ;
    END
  END dout1[57]
  PIN dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 770.480 4.000 771.080 ;
    END
  END dout1[58]
  PIN dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 774.560 4.000 775.160 ;
    END
  END dout1[59]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END dout1[5]
  PIN dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END dout1[60]
  PIN dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.720 4.000 783.320 ;
    END
  END dout1[61]
  PIN dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.800 4.000 787.400 ;
    END
  END dout1[62]
  PIN dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.880 4.000 791.480 ;
    END
  END dout1[63]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 558.320 4.000 558.920 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 4.000 567.080 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END dout1[9]
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END irq[0]
  PIN irq[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END irq[10]
  PIN irq[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END irq[11]
  PIN irq[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END irq[12]
  PIN irq[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END irq[13]
  PIN irq[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END irq[14]
  PIN irq[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END irq[15]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END irq[2]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END irq[5]
  PIN irq[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END irq[6]
  PIN irq[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END irq[7]
  PIN irq[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END irq[8]
  PIN irq[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END irq[9]
  PIN jtag_tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END jtag_tms
  PIN localMemory_wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 411.440 500.000 412.040 ;
    END
  END localMemory_wb_ack_o
  PIN localMemory_wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 431.840 500.000 432.440 ;
    END
  END localMemory_wb_adr_i[0]
  PIN localMemory_wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 547.440 500.000 548.040 ;
    END
  END localMemory_wb_adr_i[10]
  PIN localMemory_wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 557.640 500.000 558.240 ;
    END
  END localMemory_wb_adr_i[11]
  PIN localMemory_wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 567.840 500.000 568.440 ;
    END
  END localMemory_wb_adr_i[12]
  PIN localMemory_wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 578.040 500.000 578.640 ;
    END
  END localMemory_wb_adr_i[13]
  PIN localMemory_wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 588.240 500.000 588.840 ;
    END
  END localMemory_wb_adr_i[14]
  PIN localMemory_wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 598.440 500.000 599.040 ;
    END
  END localMemory_wb_adr_i[15]
  PIN localMemory_wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 608.640 500.000 609.240 ;
    END
  END localMemory_wb_adr_i[16]
  PIN localMemory_wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 618.840 500.000 619.440 ;
    END
  END localMemory_wb_adr_i[17]
  PIN localMemory_wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 629.040 500.000 629.640 ;
    END
  END localMemory_wb_adr_i[18]
  PIN localMemory_wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 639.240 500.000 639.840 ;
    END
  END localMemory_wb_adr_i[19]
  PIN localMemory_wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 445.440 500.000 446.040 ;
    END
  END localMemory_wb_adr_i[1]
  PIN localMemory_wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 649.440 500.000 650.040 ;
    END
  END localMemory_wb_adr_i[20]
  PIN localMemory_wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 659.640 500.000 660.240 ;
    END
  END localMemory_wb_adr_i[21]
  PIN localMemory_wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 669.840 500.000 670.440 ;
    END
  END localMemory_wb_adr_i[22]
  PIN localMemory_wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 680.040 500.000 680.640 ;
    END
  END localMemory_wb_adr_i[23]
  PIN localMemory_wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 459.040 500.000 459.640 ;
    END
  END localMemory_wb_adr_i[2]
  PIN localMemory_wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 472.640 500.000 473.240 ;
    END
  END localMemory_wb_adr_i[3]
  PIN localMemory_wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 486.240 500.000 486.840 ;
    END
  END localMemory_wb_adr_i[4]
  PIN localMemory_wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 496.440 500.000 497.040 ;
    END
  END localMemory_wb_adr_i[5]
  PIN localMemory_wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 506.640 500.000 507.240 ;
    END
  END localMemory_wb_adr_i[6]
  PIN localMemory_wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 516.840 500.000 517.440 ;
    END
  END localMemory_wb_adr_i[7]
  PIN localMemory_wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 527.040 500.000 527.640 ;
    END
  END localMemory_wb_adr_i[8]
  PIN localMemory_wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 537.240 500.000 537.840 ;
    END
  END localMemory_wb_adr_i[9]
  PIN localMemory_wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 414.840 500.000 415.440 ;
    END
  END localMemory_wb_cyc_i
  PIN localMemory_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 435.240 500.000 435.840 ;
    END
  END localMemory_wb_data_i[0]
  PIN localMemory_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 550.840 500.000 551.440 ;
    END
  END localMemory_wb_data_i[10]
  PIN localMemory_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 561.040 500.000 561.640 ;
    END
  END localMemory_wb_data_i[11]
  PIN localMemory_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 571.240 500.000 571.840 ;
    END
  END localMemory_wb_data_i[12]
  PIN localMemory_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 581.440 500.000 582.040 ;
    END
  END localMemory_wb_data_i[13]
  PIN localMemory_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 591.640 500.000 592.240 ;
    END
  END localMemory_wb_data_i[14]
  PIN localMemory_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 601.840 500.000 602.440 ;
    END
  END localMemory_wb_data_i[15]
  PIN localMemory_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 612.040 500.000 612.640 ;
    END
  END localMemory_wb_data_i[16]
  PIN localMemory_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 622.240 500.000 622.840 ;
    END
  END localMemory_wb_data_i[17]
  PIN localMemory_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 632.440 500.000 633.040 ;
    END
  END localMemory_wb_data_i[18]
  PIN localMemory_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 642.640 500.000 643.240 ;
    END
  END localMemory_wb_data_i[19]
  PIN localMemory_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 448.840 500.000 449.440 ;
    END
  END localMemory_wb_data_i[1]
  PIN localMemory_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 652.840 500.000 653.440 ;
    END
  END localMemory_wb_data_i[20]
  PIN localMemory_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 663.040 500.000 663.640 ;
    END
  END localMemory_wb_data_i[21]
  PIN localMemory_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 673.240 500.000 673.840 ;
    END
  END localMemory_wb_data_i[22]
  PIN localMemory_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 683.440 500.000 684.040 ;
    END
  END localMemory_wb_data_i[23]
  PIN localMemory_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 690.240 500.000 690.840 ;
    END
  END localMemory_wb_data_i[24]
  PIN localMemory_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 697.040 500.000 697.640 ;
    END
  END localMemory_wb_data_i[25]
  PIN localMemory_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 703.840 500.000 704.440 ;
    END
  END localMemory_wb_data_i[26]
  PIN localMemory_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 710.640 500.000 711.240 ;
    END
  END localMemory_wb_data_i[27]
  PIN localMemory_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 717.440 500.000 718.040 ;
    END
  END localMemory_wb_data_i[28]
  PIN localMemory_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 724.240 500.000 724.840 ;
    END
  END localMemory_wb_data_i[29]
  PIN localMemory_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 462.440 500.000 463.040 ;
    END
  END localMemory_wb_data_i[2]
  PIN localMemory_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 731.040 500.000 731.640 ;
    END
  END localMemory_wb_data_i[30]
  PIN localMemory_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 737.840 500.000 738.440 ;
    END
  END localMemory_wb_data_i[31]
  PIN localMemory_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 476.040 500.000 476.640 ;
    END
  END localMemory_wb_data_i[3]
  PIN localMemory_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 489.640 500.000 490.240 ;
    END
  END localMemory_wb_data_i[4]
  PIN localMemory_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 499.840 500.000 500.440 ;
    END
  END localMemory_wb_data_i[5]
  PIN localMemory_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 510.040 500.000 510.640 ;
    END
  END localMemory_wb_data_i[6]
  PIN localMemory_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 520.240 500.000 520.840 ;
    END
  END localMemory_wb_data_i[7]
  PIN localMemory_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 530.440 500.000 531.040 ;
    END
  END localMemory_wb_data_i[8]
  PIN localMemory_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 540.640 500.000 541.240 ;
    END
  END localMemory_wb_data_i[9]
  PIN localMemory_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 438.640 500.000 439.240 ;
    END
  END localMemory_wb_data_o[0]
  PIN localMemory_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 554.240 500.000 554.840 ;
    END
  END localMemory_wb_data_o[10]
  PIN localMemory_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 564.440 500.000 565.040 ;
    END
  END localMemory_wb_data_o[11]
  PIN localMemory_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 574.640 500.000 575.240 ;
    END
  END localMemory_wb_data_o[12]
  PIN localMemory_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 584.840 500.000 585.440 ;
    END
  END localMemory_wb_data_o[13]
  PIN localMemory_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 595.040 500.000 595.640 ;
    END
  END localMemory_wb_data_o[14]
  PIN localMemory_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 605.240 500.000 605.840 ;
    END
  END localMemory_wb_data_o[15]
  PIN localMemory_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 615.440 500.000 616.040 ;
    END
  END localMemory_wb_data_o[16]
  PIN localMemory_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 625.640 500.000 626.240 ;
    END
  END localMemory_wb_data_o[17]
  PIN localMemory_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 635.840 500.000 636.440 ;
    END
  END localMemory_wb_data_o[18]
  PIN localMemory_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 646.040 500.000 646.640 ;
    END
  END localMemory_wb_data_o[19]
  PIN localMemory_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 452.240 500.000 452.840 ;
    END
  END localMemory_wb_data_o[1]
  PIN localMemory_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 656.240 500.000 656.840 ;
    END
  END localMemory_wb_data_o[20]
  PIN localMemory_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 666.440 500.000 667.040 ;
    END
  END localMemory_wb_data_o[21]
  PIN localMemory_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 676.640 500.000 677.240 ;
    END
  END localMemory_wb_data_o[22]
  PIN localMemory_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 686.840 500.000 687.440 ;
    END
  END localMemory_wb_data_o[23]
  PIN localMemory_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 693.640 500.000 694.240 ;
    END
  END localMemory_wb_data_o[24]
  PIN localMemory_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 700.440 500.000 701.040 ;
    END
  END localMemory_wb_data_o[25]
  PIN localMemory_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 707.240 500.000 707.840 ;
    END
  END localMemory_wb_data_o[26]
  PIN localMemory_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 714.040 500.000 714.640 ;
    END
  END localMemory_wb_data_o[27]
  PIN localMemory_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 720.840 500.000 721.440 ;
    END
  END localMemory_wb_data_o[28]
  PIN localMemory_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 727.640 500.000 728.240 ;
    END
  END localMemory_wb_data_o[29]
  PIN localMemory_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 465.840 500.000 466.440 ;
    END
  END localMemory_wb_data_o[2]
  PIN localMemory_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 734.440 500.000 735.040 ;
    END
  END localMemory_wb_data_o[30]
  PIN localMemory_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 741.240 500.000 741.840 ;
    END
  END localMemory_wb_data_o[31]
  PIN localMemory_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 479.440 500.000 480.040 ;
    END
  END localMemory_wb_data_o[3]
  PIN localMemory_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 493.040 500.000 493.640 ;
    END
  END localMemory_wb_data_o[4]
  PIN localMemory_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 503.240 500.000 503.840 ;
    END
  END localMemory_wb_data_o[5]
  PIN localMemory_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 513.440 500.000 514.040 ;
    END
  END localMemory_wb_data_o[6]
  PIN localMemory_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 523.640 500.000 524.240 ;
    END
  END localMemory_wb_data_o[7]
  PIN localMemory_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 533.840 500.000 534.440 ;
    END
  END localMemory_wb_data_o[8]
  PIN localMemory_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 544.040 500.000 544.640 ;
    END
  END localMemory_wb_data_o[9]
  PIN localMemory_wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 418.240 500.000 418.840 ;
    END
  END localMemory_wb_error_o
  PIN localMemory_wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 442.040 500.000 442.640 ;
    END
  END localMemory_wb_sel_i[0]
  PIN localMemory_wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 455.640 500.000 456.240 ;
    END
  END localMemory_wb_sel_i[1]
  PIN localMemory_wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 469.240 500.000 469.840 ;
    END
  END localMemory_wb_sel_i[2]
  PIN localMemory_wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 482.840 500.000 483.440 ;
    END
  END localMemory_wb_sel_i[3]
  PIN localMemory_wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 421.640 500.000 422.240 ;
    END
  END localMemory_wb_stall_o
  PIN localMemory_wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 425.040 500.000 425.640 ;
    END
  END localMemory_wb_stb_i
  PIN localMemory_wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 428.440 500.000 429.040 ;
    END
  END localMemory_wb_we_i
  PIN manufacturerID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 796.000 113.530 800.000 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 796.000 237.730 800.000 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 796.000 125.950 800.000 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 796.000 138.370 800.000 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 796.000 150.790 800.000 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 796.000 163.210 800.000 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 796.000 175.630 800.000 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 796.000 188.050 800.000 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 796.000 200.470 800.000 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 796.000 212.890 800.000 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 796.000 225.310 800.000 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 796.000 250.150 800.000 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 796.000 374.350 800.000 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 796.000 386.770 800.000 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 796.000 399.190 800.000 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 796.000 411.610 800.000 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 796.000 424.030 800.000 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 796.000 436.450 800.000 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 796.000 262.570 800.000 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 796.000 274.990 800.000 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 796.000 287.410 800.000 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 796.000 299.830 800.000 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 796.000 312.250 800.000 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 796.000 324.670 800.000 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 796.000 337.090 800.000 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 796.000 349.510 800.000 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 796.000 361.930 800.000 ;
    END
  END partID[9]
  PIN probe_env[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END probe_env[0]
  PIN probe_env[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END probe_env[1]
  PIN probe_jtagInstruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END probe_jtagInstruction[0]
  PIN probe_jtagInstruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END probe_jtagInstruction[1]
  PIN probe_jtagInstruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END probe_jtagInstruction[2]
  PIN probe_jtagInstruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END probe_jtagInstruction[3]
  PIN probe_jtagInstruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END probe_jtagInstruction[4]
  PIN probe_programCounter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END probe_programCounter[0]
  PIN probe_programCounter[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END probe_programCounter[10]
  PIN probe_programCounter[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END probe_programCounter[11]
  PIN probe_programCounter[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END probe_programCounter[12]
  PIN probe_programCounter[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END probe_programCounter[13]
  PIN probe_programCounter[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END probe_programCounter[14]
  PIN probe_programCounter[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END probe_programCounter[15]
  PIN probe_programCounter[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END probe_programCounter[16]
  PIN probe_programCounter[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END probe_programCounter[17]
  PIN probe_programCounter[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END probe_programCounter[18]
  PIN probe_programCounter[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END probe_programCounter[19]
  PIN probe_programCounter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END probe_programCounter[1]
  PIN probe_programCounter[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END probe_programCounter[20]
  PIN probe_programCounter[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END probe_programCounter[21]
  PIN probe_programCounter[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END probe_programCounter[22]
  PIN probe_programCounter[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END probe_programCounter[23]
  PIN probe_programCounter[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END probe_programCounter[24]
  PIN probe_programCounter[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END probe_programCounter[25]
  PIN probe_programCounter[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END probe_programCounter[26]
  PIN probe_programCounter[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END probe_programCounter[27]
  PIN probe_programCounter[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END probe_programCounter[28]
  PIN probe_programCounter[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END probe_programCounter[29]
  PIN probe_programCounter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END probe_programCounter[2]
  PIN probe_programCounter[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END probe_programCounter[30]
  PIN probe_programCounter[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END probe_programCounter[31]
  PIN probe_programCounter[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END probe_programCounter[3]
  PIN probe_programCounter[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END probe_programCounter[4]
  PIN probe_programCounter[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END probe_programCounter[5]
  PIN probe_programCounter[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END probe_programCounter[6]
  PIN probe_programCounter[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END probe_programCounter[7]
  PIN probe_programCounter[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END probe_programCounter[8]
  PIN probe_programCounter[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END probe_programCounter[9]
  PIN probe_state
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END probe_state
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 796.000 448.870 800.000 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 796.000 461.290 800.000 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 796.000 473.710 800.000 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 796.000 486.130 800.000 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 57.840 500.000 58.440 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 61.240 500.000 61.840 ;
    END
  END wb_rst_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 788.885 ;
      LAYER met1 ;
        RECT 0.990 4.460 499.950 793.520 ;
      LAYER met2 ;
        RECT 1.020 795.720 13.610 796.690 ;
        RECT 14.450 795.720 26.030 796.690 ;
        RECT 26.870 795.720 38.450 796.690 ;
        RECT 39.290 795.720 50.870 796.690 ;
        RECT 51.710 795.720 63.290 796.690 ;
        RECT 64.130 795.720 75.710 796.690 ;
        RECT 76.550 795.720 88.130 796.690 ;
        RECT 88.970 795.720 100.550 796.690 ;
        RECT 101.390 795.720 112.970 796.690 ;
        RECT 113.810 795.720 125.390 796.690 ;
        RECT 126.230 795.720 137.810 796.690 ;
        RECT 138.650 795.720 150.230 796.690 ;
        RECT 151.070 795.720 162.650 796.690 ;
        RECT 163.490 795.720 175.070 796.690 ;
        RECT 175.910 795.720 187.490 796.690 ;
        RECT 188.330 795.720 199.910 796.690 ;
        RECT 200.750 795.720 212.330 796.690 ;
        RECT 213.170 795.720 224.750 796.690 ;
        RECT 225.590 795.720 237.170 796.690 ;
        RECT 238.010 795.720 249.590 796.690 ;
        RECT 250.430 795.720 262.010 796.690 ;
        RECT 262.850 795.720 274.430 796.690 ;
        RECT 275.270 795.720 286.850 796.690 ;
        RECT 287.690 795.720 299.270 796.690 ;
        RECT 300.110 795.720 311.690 796.690 ;
        RECT 312.530 795.720 324.110 796.690 ;
        RECT 324.950 795.720 336.530 796.690 ;
        RECT 337.370 795.720 348.950 796.690 ;
        RECT 349.790 795.720 361.370 796.690 ;
        RECT 362.210 795.720 373.790 796.690 ;
        RECT 374.630 795.720 386.210 796.690 ;
        RECT 387.050 795.720 398.630 796.690 ;
        RECT 399.470 795.720 411.050 796.690 ;
        RECT 411.890 795.720 423.470 796.690 ;
        RECT 424.310 795.720 435.890 796.690 ;
        RECT 436.730 795.720 448.310 796.690 ;
        RECT 449.150 795.720 460.730 796.690 ;
        RECT 461.570 795.720 473.150 796.690 ;
        RECT 473.990 795.720 485.570 796.690 ;
        RECT 486.410 795.720 499.920 796.690 ;
        RECT 1.020 4.280 499.920 795.720 ;
        RECT 1.020 3.670 9.010 4.280 ;
        RECT 9.850 3.670 17.750 4.280 ;
        RECT 18.590 3.670 26.490 4.280 ;
        RECT 27.330 3.670 35.230 4.280 ;
        RECT 36.070 3.670 43.970 4.280 ;
        RECT 44.810 3.670 52.710 4.280 ;
        RECT 53.550 3.670 61.450 4.280 ;
        RECT 62.290 3.670 70.190 4.280 ;
        RECT 71.030 3.670 78.930 4.280 ;
        RECT 79.770 3.670 87.670 4.280 ;
        RECT 88.510 3.670 96.410 4.280 ;
        RECT 97.250 3.670 105.150 4.280 ;
        RECT 105.990 3.670 113.890 4.280 ;
        RECT 114.730 3.670 122.630 4.280 ;
        RECT 123.470 3.670 131.370 4.280 ;
        RECT 132.210 3.670 140.110 4.280 ;
        RECT 140.950 3.670 148.850 4.280 ;
        RECT 149.690 3.670 157.590 4.280 ;
        RECT 158.430 3.670 166.330 4.280 ;
        RECT 167.170 3.670 175.070 4.280 ;
        RECT 175.910 3.670 183.810 4.280 ;
        RECT 184.650 3.670 192.550 4.280 ;
        RECT 193.390 3.670 201.290 4.280 ;
        RECT 202.130 3.670 210.030 4.280 ;
        RECT 210.870 3.670 218.770 4.280 ;
        RECT 219.610 3.670 227.510 4.280 ;
        RECT 228.350 3.670 236.250 4.280 ;
        RECT 237.090 3.670 244.990 4.280 ;
        RECT 245.830 3.670 253.730 4.280 ;
        RECT 254.570 3.670 262.470 4.280 ;
        RECT 263.310 3.670 271.210 4.280 ;
        RECT 272.050 3.670 279.950 4.280 ;
        RECT 280.790 3.670 288.690 4.280 ;
        RECT 289.530 3.670 297.430 4.280 ;
        RECT 298.270 3.670 306.170 4.280 ;
        RECT 307.010 3.670 314.910 4.280 ;
        RECT 315.750 3.670 323.650 4.280 ;
        RECT 324.490 3.670 332.390 4.280 ;
        RECT 333.230 3.670 341.130 4.280 ;
        RECT 341.970 3.670 349.870 4.280 ;
        RECT 350.710 3.670 358.610 4.280 ;
        RECT 359.450 3.670 367.350 4.280 ;
        RECT 368.190 3.670 376.090 4.280 ;
        RECT 376.930 3.670 384.830 4.280 ;
        RECT 385.670 3.670 393.570 4.280 ;
        RECT 394.410 3.670 402.310 4.280 ;
        RECT 403.150 3.670 411.050 4.280 ;
        RECT 411.890 3.670 419.790 4.280 ;
        RECT 420.630 3.670 428.530 4.280 ;
        RECT 429.370 3.670 437.270 4.280 ;
        RECT 438.110 3.670 446.010 4.280 ;
        RECT 446.850 3.670 454.750 4.280 ;
        RECT 455.590 3.670 463.490 4.280 ;
        RECT 464.330 3.670 472.230 4.280 ;
        RECT 473.070 3.670 480.970 4.280 ;
        RECT 481.810 3.670 489.710 4.280 ;
        RECT 490.550 3.670 499.920 4.280 ;
      LAYER met3 ;
        RECT 4.400 790.480 499.035 791.345 ;
        RECT 1.190 787.800 499.035 790.480 ;
        RECT 4.400 786.400 499.035 787.800 ;
        RECT 1.190 783.720 499.035 786.400 ;
        RECT 4.400 782.320 499.035 783.720 ;
        RECT 1.190 779.640 499.035 782.320 ;
        RECT 4.400 778.240 499.035 779.640 ;
        RECT 1.190 775.560 499.035 778.240 ;
        RECT 4.400 774.160 499.035 775.560 ;
        RECT 1.190 771.480 499.035 774.160 ;
        RECT 4.400 770.080 499.035 771.480 ;
        RECT 1.190 767.400 499.035 770.080 ;
        RECT 4.400 766.000 499.035 767.400 ;
        RECT 1.190 763.320 499.035 766.000 ;
        RECT 4.400 761.920 499.035 763.320 ;
        RECT 1.190 759.240 499.035 761.920 ;
        RECT 4.400 757.840 499.035 759.240 ;
        RECT 1.190 755.160 499.035 757.840 ;
        RECT 4.400 753.760 499.035 755.160 ;
        RECT 1.190 751.080 499.035 753.760 ;
        RECT 4.400 749.680 499.035 751.080 ;
        RECT 1.190 747.000 499.035 749.680 ;
        RECT 4.400 745.600 499.035 747.000 ;
        RECT 1.190 742.920 499.035 745.600 ;
        RECT 4.400 742.240 499.035 742.920 ;
        RECT 4.400 741.520 495.600 742.240 ;
        RECT 1.190 740.840 495.600 741.520 ;
        RECT 1.190 738.840 499.035 740.840 ;
        RECT 4.400 737.440 495.600 738.840 ;
        RECT 1.190 735.440 499.035 737.440 ;
        RECT 1.190 734.760 495.600 735.440 ;
        RECT 4.400 734.040 495.600 734.760 ;
        RECT 4.400 733.360 499.035 734.040 ;
        RECT 1.190 732.040 499.035 733.360 ;
        RECT 1.190 730.680 495.600 732.040 ;
        RECT 4.400 730.640 495.600 730.680 ;
        RECT 4.400 729.280 499.035 730.640 ;
        RECT 1.190 728.640 499.035 729.280 ;
        RECT 1.190 727.240 495.600 728.640 ;
        RECT 1.190 726.600 499.035 727.240 ;
        RECT 4.400 725.240 499.035 726.600 ;
        RECT 4.400 725.200 495.600 725.240 ;
        RECT 1.190 723.840 495.600 725.200 ;
        RECT 1.190 722.520 499.035 723.840 ;
        RECT 4.400 721.840 499.035 722.520 ;
        RECT 4.400 721.120 495.600 721.840 ;
        RECT 1.190 720.440 495.600 721.120 ;
        RECT 1.190 718.440 499.035 720.440 ;
        RECT 4.400 717.040 495.600 718.440 ;
        RECT 1.190 715.040 499.035 717.040 ;
        RECT 1.190 714.360 495.600 715.040 ;
        RECT 4.400 713.640 495.600 714.360 ;
        RECT 4.400 712.960 499.035 713.640 ;
        RECT 1.190 711.640 499.035 712.960 ;
        RECT 1.190 710.280 495.600 711.640 ;
        RECT 4.400 710.240 495.600 710.280 ;
        RECT 4.400 708.880 499.035 710.240 ;
        RECT 1.190 708.240 499.035 708.880 ;
        RECT 1.190 706.840 495.600 708.240 ;
        RECT 1.190 706.200 499.035 706.840 ;
        RECT 4.400 704.840 499.035 706.200 ;
        RECT 4.400 704.800 495.600 704.840 ;
        RECT 1.190 703.440 495.600 704.800 ;
        RECT 1.190 702.120 499.035 703.440 ;
        RECT 4.400 701.440 499.035 702.120 ;
        RECT 4.400 700.720 495.600 701.440 ;
        RECT 1.190 700.040 495.600 700.720 ;
        RECT 1.190 698.040 499.035 700.040 ;
        RECT 4.400 696.640 495.600 698.040 ;
        RECT 1.190 694.640 499.035 696.640 ;
        RECT 1.190 693.960 495.600 694.640 ;
        RECT 4.400 693.240 495.600 693.960 ;
        RECT 4.400 692.560 499.035 693.240 ;
        RECT 1.190 691.240 499.035 692.560 ;
        RECT 1.190 689.880 495.600 691.240 ;
        RECT 4.400 689.840 495.600 689.880 ;
        RECT 4.400 688.480 499.035 689.840 ;
        RECT 1.190 687.840 499.035 688.480 ;
        RECT 1.190 686.440 495.600 687.840 ;
        RECT 1.190 685.800 499.035 686.440 ;
        RECT 4.400 684.440 499.035 685.800 ;
        RECT 4.400 684.400 495.600 684.440 ;
        RECT 1.190 683.040 495.600 684.400 ;
        RECT 1.190 681.720 499.035 683.040 ;
        RECT 4.400 681.040 499.035 681.720 ;
        RECT 4.400 680.320 495.600 681.040 ;
        RECT 1.190 679.640 495.600 680.320 ;
        RECT 1.190 677.640 499.035 679.640 ;
        RECT 4.400 676.240 495.600 677.640 ;
        RECT 1.190 674.240 499.035 676.240 ;
        RECT 1.190 673.560 495.600 674.240 ;
        RECT 4.400 672.840 495.600 673.560 ;
        RECT 4.400 672.160 499.035 672.840 ;
        RECT 1.190 670.840 499.035 672.160 ;
        RECT 1.190 669.480 495.600 670.840 ;
        RECT 4.400 669.440 495.600 669.480 ;
        RECT 4.400 668.080 499.035 669.440 ;
        RECT 1.190 667.440 499.035 668.080 ;
        RECT 1.190 666.040 495.600 667.440 ;
        RECT 1.190 665.400 499.035 666.040 ;
        RECT 4.400 664.040 499.035 665.400 ;
        RECT 4.400 664.000 495.600 664.040 ;
        RECT 1.190 662.640 495.600 664.000 ;
        RECT 1.190 661.320 499.035 662.640 ;
        RECT 4.400 660.640 499.035 661.320 ;
        RECT 4.400 659.920 495.600 660.640 ;
        RECT 1.190 659.240 495.600 659.920 ;
        RECT 1.190 657.240 499.035 659.240 ;
        RECT 4.400 655.840 495.600 657.240 ;
        RECT 1.190 653.840 499.035 655.840 ;
        RECT 1.190 653.160 495.600 653.840 ;
        RECT 4.400 652.440 495.600 653.160 ;
        RECT 4.400 651.760 499.035 652.440 ;
        RECT 1.190 650.440 499.035 651.760 ;
        RECT 1.190 649.080 495.600 650.440 ;
        RECT 4.400 649.040 495.600 649.080 ;
        RECT 4.400 647.680 499.035 649.040 ;
        RECT 1.190 647.040 499.035 647.680 ;
        RECT 1.190 645.640 495.600 647.040 ;
        RECT 1.190 645.000 499.035 645.640 ;
        RECT 4.400 643.640 499.035 645.000 ;
        RECT 4.400 643.600 495.600 643.640 ;
        RECT 1.190 642.240 495.600 643.600 ;
        RECT 1.190 640.920 499.035 642.240 ;
        RECT 4.400 640.240 499.035 640.920 ;
        RECT 4.400 639.520 495.600 640.240 ;
        RECT 1.190 638.840 495.600 639.520 ;
        RECT 1.190 636.840 499.035 638.840 ;
        RECT 4.400 635.440 495.600 636.840 ;
        RECT 1.190 633.440 499.035 635.440 ;
        RECT 1.190 632.760 495.600 633.440 ;
        RECT 4.400 632.040 495.600 632.760 ;
        RECT 4.400 631.360 499.035 632.040 ;
        RECT 1.190 630.040 499.035 631.360 ;
        RECT 1.190 628.680 495.600 630.040 ;
        RECT 4.400 628.640 495.600 628.680 ;
        RECT 4.400 627.280 499.035 628.640 ;
        RECT 1.190 626.640 499.035 627.280 ;
        RECT 1.190 625.240 495.600 626.640 ;
        RECT 1.190 624.600 499.035 625.240 ;
        RECT 4.400 623.240 499.035 624.600 ;
        RECT 4.400 623.200 495.600 623.240 ;
        RECT 1.190 621.840 495.600 623.200 ;
        RECT 1.190 620.520 499.035 621.840 ;
        RECT 4.400 619.840 499.035 620.520 ;
        RECT 4.400 619.120 495.600 619.840 ;
        RECT 1.190 618.440 495.600 619.120 ;
        RECT 1.190 616.440 499.035 618.440 ;
        RECT 4.400 615.040 495.600 616.440 ;
        RECT 1.190 613.040 499.035 615.040 ;
        RECT 1.190 612.360 495.600 613.040 ;
        RECT 4.400 611.640 495.600 612.360 ;
        RECT 4.400 610.960 499.035 611.640 ;
        RECT 1.190 609.640 499.035 610.960 ;
        RECT 1.190 608.280 495.600 609.640 ;
        RECT 4.400 608.240 495.600 608.280 ;
        RECT 4.400 606.880 499.035 608.240 ;
        RECT 1.190 606.240 499.035 606.880 ;
        RECT 1.190 604.840 495.600 606.240 ;
        RECT 1.190 604.200 499.035 604.840 ;
        RECT 4.400 602.840 499.035 604.200 ;
        RECT 4.400 602.800 495.600 602.840 ;
        RECT 1.190 601.440 495.600 602.800 ;
        RECT 1.190 600.120 499.035 601.440 ;
        RECT 4.400 599.440 499.035 600.120 ;
        RECT 4.400 598.720 495.600 599.440 ;
        RECT 1.190 598.040 495.600 598.720 ;
        RECT 1.190 596.040 499.035 598.040 ;
        RECT 4.400 594.640 495.600 596.040 ;
        RECT 1.190 592.640 499.035 594.640 ;
        RECT 1.190 591.960 495.600 592.640 ;
        RECT 4.400 591.240 495.600 591.960 ;
        RECT 4.400 590.560 499.035 591.240 ;
        RECT 1.190 589.240 499.035 590.560 ;
        RECT 1.190 587.880 495.600 589.240 ;
        RECT 4.400 587.840 495.600 587.880 ;
        RECT 4.400 586.480 499.035 587.840 ;
        RECT 1.190 585.840 499.035 586.480 ;
        RECT 1.190 584.440 495.600 585.840 ;
        RECT 1.190 583.800 499.035 584.440 ;
        RECT 4.400 582.440 499.035 583.800 ;
        RECT 4.400 582.400 495.600 582.440 ;
        RECT 1.190 581.040 495.600 582.400 ;
        RECT 1.190 579.720 499.035 581.040 ;
        RECT 4.400 579.040 499.035 579.720 ;
        RECT 4.400 578.320 495.600 579.040 ;
        RECT 1.190 577.640 495.600 578.320 ;
        RECT 1.190 575.640 499.035 577.640 ;
        RECT 4.400 574.240 495.600 575.640 ;
        RECT 1.190 572.240 499.035 574.240 ;
        RECT 1.190 571.560 495.600 572.240 ;
        RECT 4.400 570.840 495.600 571.560 ;
        RECT 4.400 570.160 499.035 570.840 ;
        RECT 1.190 568.840 499.035 570.160 ;
        RECT 1.190 567.480 495.600 568.840 ;
        RECT 4.400 567.440 495.600 567.480 ;
        RECT 4.400 566.080 499.035 567.440 ;
        RECT 1.190 565.440 499.035 566.080 ;
        RECT 1.190 564.040 495.600 565.440 ;
        RECT 1.190 563.400 499.035 564.040 ;
        RECT 4.400 562.040 499.035 563.400 ;
        RECT 4.400 562.000 495.600 562.040 ;
        RECT 1.190 560.640 495.600 562.000 ;
        RECT 1.190 559.320 499.035 560.640 ;
        RECT 4.400 558.640 499.035 559.320 ;
        RECT 4.400 557.920 495.600 558.640 ;
        RECT 1.190 557.240 495.600 557.920 ;
        RECT 1.190 555.240 499.035 557.240 ;
        RECT 4.400 553.840 495.600 555.240 ;
        RECT 1.190 551.840 499.035 553.840 ;
        RECT 1.190 551.160 495.600 551.840 ;
        RECT 4.400 550.440 495.600 551.160 ;
        RECT 4.400 549.760 499.035 550.440 ;
        RECT 1.190 548.440 499.035 549.760 ;
        RECT 1.190 547.080 495.600 548.440 ;
        RECT 4.400 547.040 495.600 547.080 ;
        RECT 4.400 545.680 499.035 547.040 ;
        RECT 1.190 545.040 499.035 545.680 ;
        RECT 1.190 543.640 495.600 545.040 ;
        RECT 1.190 543.000 499.035 543.640 ;
        RECT 4.400 541.640 499.035 543.000 ;
        RECT 4.400 541.600 495.600 541.640 ;
        RECT 1.190 540.240 495.600 541.600 ;
        RECT 1.190 538.920 499.035 540.240 ;
        RECT 4.400 538.240 499.035 538.920 ;
        RECT 4.400 537.520 495.600 538.240 ;
        RECT 1.190 536.840 495.600 537.520 ;
        RECT 1.190 534.840 499.035 536.840 ;
        RECT 4.400 533.440 495.600 534.840 ;
        RECT 1.190 531.440 499.035 533.440 ;
        RECT 1.190 530.760 495.600 531.440 ;
        RECT 4.400 530.040 495.600 530.760 ;
        RECT 4.400 529.360 499.035 530.040 ;
        RECT 1.190 528.040 499.035 529.360 ;
        RECT 1.190 526.680 495.600 528.040 ;
        RECT 4.400 526.640 495.600 526.680 ;
        RECT 4.400 525.280 499.035 526.640 ;
        RECT 1.190 524.640 499.035 525.280 ;
        RECT 1.190 523.240 495.600 524.640 ;
        RECT 1.190 522.600 499.035 523.240 ;
        RECT 4.400 521.240 499.035 522.600 ;
        RECT 4.400 521.200 495.600 521.240 ;
        RECT 1.190 519.840 495.600 521.200 ;
        RECT 1.190 518.520 499.035 519.840 ;
        RECT 4.400 517.840 499.035 518.520 ;
        RECT 4.400 517.120 495.600 517.840 ;
        RECT 1.190 516.440 495.600 517.120 ;
        RECT 1.190 514.440 499.035 516.440 ;
        RECT 4.400 513.040 495.600 514.440 ;
        RECT 1.190 511.040 499.035 513.040 ;
        RECT 1.190 510.360 495.600 511.040 ;
        RECT 4.400 509.640 495.600 510.360 ;
        RECT 4.400 508.960 499.035 509.640 ;
        RECT 1.190 507.640 499.035 508.960 ;
        RECT 1.190 506.280 495.600 507.640 ;
        RECT 4.400 506.240 495.600 506.280 ;
        RECT 4.400 504.880 499.035 506.240 ;
        RECT 1.190 504.240 499.035 504.880 ;
        RECT 1.190 502.840 495.600 504.240 ;
        RECT 1.190 502.200 499.035 502.840 ;
        RECT 4.400 500.840 499.035 502.200 ;
        RECT 4.400 500.800 495.600 500.840 ;
        RECT 1.190 499.440 495.600 500.800 ;
        RECT 1.190 498.120 499.035 499.440 ;
        RECT 4.400 497.440 499.035 498.120 ;
        RECT 4.400 496.720 495.600 497.440 ;
        RECT 1.190 496.040 495.600 496.720 ;
        RECT 1.190 494.040 499.035 496.040 ;
        RECT 4.400 492.640 495.600 494.040 ;
        RECT 1.190 490.640 499.035 492.640 ;
        RECT 1.190 489.960 495.600 490.640 ;
        RECT 4.400 489.240 495.600 489.960 ;
        RECT 4.400 488.560 499.035 489.240 ;
        RECT 1.190 487.240 499.035 488.560 ;
        RECT 1.190 485.880 495.600 487.240 ;
        RECT 4.400 485.840 495.600 485.880 ;
        RECT 4.400 484.480 499.035 485.840 ;
        RECT 1.190 483.840 499.035 484.480 ;
        RECT 1.190 482.440 495.600 483.840 ;
        RECT 1.190 481.800 499.035 482.440 ;
        RECT 4.400 480.440 499.035 481.800 ;
        RECT 4.400 480.400 495.600 480.440 ;
        RECT 1.190 479.040 495.600 480.400 ;
        RECT 1.190 477.720 499.035 479.040 ;
        RECT 4.400 477.040 499.035 477.720 ;
        RECT 4.400 476.320 495.600 477.040 ;
        RECT 1.190 475.640 495.600 476.320 ;
        RECT 1.190 473.640 499.035 475.640 ;
        RECT 4.400 472.240 495.600 473.640 ;
        RECT 1.190 470.240 499.035 472.240 ;
        RECT 1.190 469.560 495.600 470.240 ;
        RECT 4.400 468.840 495.600 469.560 ;
        RECT 4.400 468.160 499.035 468.840 ;
        RECT 1.190 466.840 499.035 468.160 ;
        RECT 1.190 465.480 495.600 466.840 ;
        RECT 4.400 465.440 495.600 465.480 ;
        RECT 4.400 464.080 499.035 465.440 ;
        RECT 1.190 463.440 499.035 464.080 ;
        RECT 1.190 462.040 495.600 463.440 ;
        RECT 1.190 461.400 499.035 462.040 ;
        RECT 4.400 460.040 499.035 461.400 ;
        RECT 4.400 460.000 495.600 460.040 ;
        RECT 1.190 458.640 495.600 460.000 ;
        RECT 1.190 457.320 499.035 458.640 ;
        RECT 4.400 456.640 499.035 457.320 ;
        RECT 4.400 455.920 495.600 456.640 ;
        RECT 1.190 455.240 495.600 455.920 ;
        RECT 1.190 453.240 499.035 455.240 ;
        RECT 4.400 451.840 495.600 453.240 ;
        RECT 1.190 449.840 499.035 451.840 ;
        RECT 1.190 449.160 495.600 449.840 ;
        RECT 4.400 448.440 495.600 449.160 ;
        RECT 4.400 447.760 499.035 448.440 ;
        RECT 1.190 446.440 499.035 447.760 ;
        RECT 1.190 445.080 495.600 446.440 ;
        RECT 4.400 445.040 495.600 445.080 ;
        RECT 4.400 443.680 499.035 445.040 ;
        RECT 1.190 443.040 499.035 443.680 ;
        RECT 1.190 441.640 495.600 443.040 ;
        RECT 1.190 441.000 499.035 441.640 ;
        RECT 4.400 439.640 499.035 441.000 ;
        RECT 4.400 439.600 495.600 439.640 ;
        RECT 1.190 438.240 495.600 439.600 ;
        RECT 1.190 436.920 499.035 438.240 ;
        RECT 4.400 436.240 499.035 436.920 ;
        RECT 4.400 435.520 495.600 436.240 ;
        RECT 1.190 434.840 495.600 435.520 ;
        RECT 1.190 432.840 499.035 434.840 ;
        RECT 4.400 431.440 495.600 432.840 ;
        RECT 1.190 429.440 499.035 431.440 ;
        RECT 1.190 428.760 495.600 429.440 ;
        RECT 4.400 428.040 495.600 428.760 ;
        RECT 4.400 427.360 499.035 428.040 ;
        RECT 1.190 426.040 499.035 427.360 ;
        RECT 1.190 424.680 495.600 426.040 ;
        RECT 4.400 424.640 495.600 424.680 ;
        RECT 4.400 423.280 499.035 424.640 ;
        RECT 1.190 422.640 499.035 423.280 ;
        RECT 1.190 421.240 495.600 422.640 ;
        RECT 1.190 420.600 499.035 421.240 ;
        RECT 4.400 419.240 499.035 420.600 ;
        RECT 4.400 419.200 495.600 419.240 ;
        RECT 1.190 417.840 495.600 419.200 ;
        RECT 1.190 416.520 499.035 417.840 ;
        RECT 4.400 415.840 499.035 416.520 ;
        RECT 4.400 415.120 495.600 415.840 ;
        RECT 1.190 414.440 495.600 415.120 ;
        RECT 1.190 412.440 499.035 414.440 ;
        RECT 4.400 411.040 495.600 412.440 ;
        RECT 1.190 409.040 499.035 411.040 ;
        RECT 1.190 408.360 495.600 409.040 ;
        RECT 4.400 407.640 495.600 408.360 ;
        RECT 4.400 406.960 499.035 407.640 ;
        RECT 1.190 405.640 499.035 406.960 ;
        RECT 1.190 404.280 495.600 405.640 ;
        RECT 4.400 404.240 495.600 404.280 ;
        RECT 4.400 402.880 499.035 404.240 ;
        RECT 1.190 402.240 499.035 402.880 ;
        RECT 1.190 400.840 495.600 402.240 ;
        RECT 1.190 400.200 499.035 400.840 ;
        RECT 4.400 398.840 499.035 400.200 ;
        RECT 4.400 398.800 495.600 398.840 ;
        RECT 1.190 397.440 495.600 398.800 ;
        RECT 1.190 396.120 499.035 397.440 ;
        RECT 4.400 395.440 499.035 396.120 ;
        RECT 4.400 394.720 495.600 395.440 ;
        RECT 1.190 394.040 495.600 394.720 ;
        RECT 1.190 392.040 499.035 394.040 ;
        RECT 4.400 390.640 495.600 392.040 ;
        RECT 1.190 388.640 499.035 390.640 ;
        RECT 1.190 387.960 495.600 388.640 ;
        RECT 4.400 387.240 495.600 387.960 ;
        RECT 4.400 386.560 499.035 387.240 ;
        RECT 1.190 385.240 499.035 386.560 ;
        RECT 1.190 383.880 495.600 385.240 ;
        RECT 4.400 383.840 495.600 383.880 ;
        RECT 4.400 382.480 499.035 383.840 ;
        RECT 1.190 381.840 499.035 382.480 ;
        RECT 1.190 380.440 495.600 381.840 ;
        RECT 1.190 379.800 499.035 380.440 ;
        RECT 4.400 378.440 499.035 379.800 ;
        RECT 4.400 378.400 495.600 378.440 ;
        RECT 1.190 377.040 495.600 378.400 ;
        RECT 1.190 375.720 499.035 377.040 ;
        RECT 4.400 375.040 499.035 375.720 ;
        RECT 4.400 374.320 495.600 375.040 ;
        RECT 1.190 373.640 495.600 374.320 ;
        RECT 1.190 371.640 499.035 373.640 ;
        RECT 4.400 370.240 495.600 371.640 ;
        RECT 1.190 368.240 499.035 370.240 ;
        RECT 1.190 367.560 495.600 368.240 ;
        RECT 4.400 366.840 495.600 367.560 ;
        RECT 4.400 366.160 499.035 366.840 ;
        RECT 1.190 364.840 499.035 366.160 ;
        RECT 1.190 363.480 495.600 364.840 ;
        RECT 4.400 363.440 495.600 363.480 ;
        RECT 4.400 362.080 499.035 363.440 ;
        RECT 1.190 361.440 499.035 362.080 ;
        RECT 1.190 360.040 495.600 361.440 ;
        RECT 1.190 359.400 499.035 360.040 ;
        RECT 4.400 358.040 499.035 359.400 ;
        RECT 4.400 358.000 495.600 358.040 ;
        RECT 1.190 356.640 495.600 358.000 ;
        RECT 1.190 355.320 499.035 356.640 ;
        RECT 4.400 354.640 499.035 355.320 ;
        RECT 4.400 353.920 495.600 354.640 ;
        RECT 1.190 353.240 495.600 353.920 ;
        RECT 1.190 351.240 499.035 353.240 ;
        RECT 4.400 349.840 495.600 351.240 ;
        RECT 1.190 347.840 499.035 349.840 ;
        RECT 1.190 347.160 495.600 347.840 ;
        RECT 4.400 346.440 495.600 347.160 ;
        RECT 4.400 345.760 499.035 346.440 ;
        RECT 1.190 344.440 499.035 345.760 ;
        RECT 1.190 343.080 495.600 344.440 ;
        RECT 4.400 343.040 495.600 343.080 ;
        RECT 4.400 341.680 499.035 343.040 ;
        RECT 1.190 341.040 499.035 341.680 ;
        RECT 1.190 339.640 495.600 341.040 ;
        RECT 1.190 339.000 499.035 339.640 ;
        RECT 4.400 337.640 499.035 339.000 ;
        RECT 4.400 337.600 495.600 337.640 ;
        RECT 1.190 336.240 495.600 337.600 ;
        RECT 1.190 334.920 499.035 336.240 ;
        RECT 4.400 334.240 499.035 334.920 ;
        RECT 4.400 333.520 495.600 334.240 ;
        RECT 1.190 332.840 495.600 333.520 ;
        RECT 1.190 330.840 499.035 332.840 ;
        RECT 4.400 329.440 495.600 330.840 ;
        RECT 1.190 327.440 499.035 329.440 ;
        RECT 1.190 326.760 495.600 327.440 ;
        RECT 4.400 326.040 495.600 326.760 ;
        RECT 4.400 325.360 499.035 326.040 ;
        RECT 1.190 324.040 499.035 325.360 ;
        RECT 1.190 322.680 495.600 324.040 ;
        RECT 4.400 322.640 495.600 322.680 ;
        RECT 4.400 321.280 499.035 322.640 ;
        RECT 1.190 320.640 499.035 321.280 ;
        RECT 1.190 319.240 495.600 320.640 ;
        RECT 1.190 318.600 499.035 319.240 ;
        RECT 4.400 317.240 499.035 318.600 ;
        RECT 4.400 317.200 495.600 317.240 ;
        RECT 1.190 315.840 495.600 317.200 ;
        RECT 1.190 314.520 499.035 315.840 ;
        RECT 4.400 313.840 499.035 314.520 ;
        RECT 4.400 313.120 495.600 313.840 ;
        RECT 1.190 312.440 495.600 313.120 ;
        RECT 1.190 310.440 499.035 312.440 ;
        RECT 4.400 309.040 495.600 310.440 ;
        RECT 1.190 307.040 499.035 309.040 ;
        RECT 1.190 306.360 495.600 307.040 ;
        RECT 4.400 305.640 495.600 306.360 ;
        RECT 4.400 304.960 499.035 305.640 ;
        RECT 1.190 303.640 499.035 304.960 ;
        RECT 1.190 302.280 495.600 303.640 ;
        RECT 4.400 302.240 495.600 302.280 ;
        RECT 4.400 300.880 499.035 302.240 ;
        RECT 1.190 300.240 499.035 300.880 ;
        RECT 1.190 298.840 495.600 300.240 ;
        RECT 1.190 298.200 499.035 298.840 ;
        RECT 4.400 296.840 499.035 298.200 ;
        RECT 4.400 296.800 495.600 296.840 ;
        RECT 1.190 295.440 495.600 296.800 ;
        RECT 1.190 294.120 499.035 295.440 ;
        RECT 4.400 293.440 499.035 294.120 ;
        RECT 4.400 292.720 495.600 293.440 ;
        RECT 1.190 292.040 495.600 292.720 ;
        RECT 1.190 290.040 499.035 292.040 ;
        RECT 4.400 288.640 495.600 290.040 ;
        RECT 1.190 286.640 499.035 288.640 ;
        RECT 1.190 285.960 495.600 286.640 ;
        RECT 4.400 285.240 495.600 285.960 ;
        RECT 4.400 284.560 499.035 285.240 ;
        RECT 1.190 283.240 499.035 284.560 ;
        RECT 1.190 281.880 495.600 283.240 ;
        RECT 4.400 281.840 495.600 281.880 ;
        RECT 4.400 280.480 499.035 281.840 ;
        RECT 1.190 279.840 499.035 280.480 ;
        RECT 1.190 278.440 495.600 279.840 ;
        RECT 1.190 277.800 499.035 278.440 ;
        RECT 4.400 276.440 499.035 277.800 ;
        RECT 4.400 276.400 495.600 276.440 ;
        RECT 1.190 275.040 495.600 276.400 ;
        RECT 1.190 273.720 499.035 275.040 ;
        RECT 4.400 273.040 499.035 273.720 ;
        RECT 4.400 272.320 495.600 273.040 ;
        RECT 1.190 271.640 495.600 272.320 ;
        RECT 1.190 269.640 499.035 271.640 ;
        RECT 4.400 268.240 495.600 269.640 ;
        RECT 1.190 266.240 499.035 268.240 ;
        RECT 1.190 265.560 495.600 266.240 ;
        RECT 4.400 264.840 495.600 265.560 ;
        RECT 4.400 264.160 499.035 264.840 ;
        RECT 1.190 262.840 499.035 264.160 ;
        RECT 1.190 261.480 495.600 262.840 ;
        RECT 4.400 261.440 495.600 261.480 ;
        RECT 4.400 260.080 499.035 261.440 ;
        RECT 1.190 259.440 499.035 260.080 ;
        RECT 1.190 258.040 495.600 259.440 ;
        RECT 1.190 257.400 499.035 258.040 ;
        RECT 4.400 256.040 499.035 257.400 ;
        RECT 4.400 256.000 495.600 256.040 ;
        RECT 1.190 254.640 495.600 256.000 ;
        RECT 1.190 253.320 499.035 254.640 ;
        RECT 4.400 252.640 499.035 253.320 ;
        RECT 4.400 251.920 495.600 252.640 ;
        RECT 1.190 251.240 495.600 251.920 ;
        RECT 1.190 249.240 499.035 251.240 ;
        RECT 4.400 247.840 495.600 249.240 ;
        RECT 1.190 245.840 499.035 247.840 ;
        RECT 1.190 245.160 495.600 245.840 ;
        RECT 4.400 244.440 495.600 245.160 ;
        RECT 4.400 243.760 499.035 244.440 ;
        RECT 1.190 242.440 499.035 243.760 ;
        RECT 1.190 241.080 495.600 242.440 ;
        RECT 4.400 241.040 495.600 241.080 ;
        RECT 4.400 239.680 499.035 241.040 ;
        RECT 1.190 239.040 499.035 239.680 ;
        RECT 1.190 237.640 495.600 239.040 ;
        RECT 1.190 237.000 499.035 237.640 ;
        RECT 4.400 235.640 499.035 237.000 ;
        RECT 4.400 235.600 495.600 235.640 ;
        RECT 1.190 234.240 495.600 235.600 ;
        RECT 1.190 232.920 499.035 234.240 ;
        RECT 4.400 232.240 499.035 232.920 ;
        RECT 4.400 231.520 495.600 232.240 ;
        RECT 1.190 230.840 495.600 231.520 ;
        RECT 1.190 228.840 499.035 230.840 ;
        RECT 4.400 227.440 495.600 228.840 ;
        RECT 1.190 225.440 499.035 227.440 ;
        RECT 1.190 224.760 495.600 225.440 ;
        RECT 4.400 224.040 495.600 224.760 ;
        RECT 4.400 223.360 499.035 224.040 ;
        RECT 1.190 222.040 499.035 223.360 ;
        RECT 1.190 220.680 495.600 222.040 ;
        RECT 4.400 220.640 495.600 220.680 ;
        RECT 4.400 219.280 499.035 220.640 ;
        RECT 1.190 218.640 499.035 219.280 ;
        RECT 1.190 217.240 495.600 218.640 ;
        RECT 1.190 216.600 499.035 217.240 ;
        RECT 4.400 215.240 499.035 216.600 ;
        RECT 4.400 215.200 495.600 215.240 ;
        RECT 1.190 213.840 495.600 215.200 ;
        RECT 1.190 212.520 499.035 213.840 ;
        RECT 4.400 211.840 499.035 212.520 ;
        RECT 4.400 211.120 495.600 211.840 ;
        RECT 1.190 210.440 495.600 211.120 ;
        RECT 1.190 208.440 499.035 210.440 ;
        RECT 4.400 207.040 495.600 208.440 ;
        RECT 1.190 205.040 499.035 207.040 ;
        RECT 1.190 204.360 495.600 205.040 ;
        RECT 4.400 203.640 495.600 204.360 ;
        RECT 4.400 202.960 499.035 203.640 ;
        RECT 1.190 201.640 499.035 202.960 ;
        RECT 1.190 200.280 495.600 201.640 ;
        RECT 4.400 200.240 495.600 200.280 ;
        RECT 4.400 198.880 499.035 200.240 ;
        RECT 1.190 198.240 499.035 198.880 ;
        RECT 1.190 196.840 495.600 198.240 ;
        RECT 1.190 196.200 499.035 196.840 ;
        RECT 4.400 194.840 499.035 196.200 ;
        RECT 4.400 194.800 495.600 194.840 ;
        RECT 1.190 193.440 495.600 194.800 ;
        RECT 1.190 192.120 499.035 193.440 ;
        RECT 4.400 191.440 499.035 192.120 ;
        RECT 4.400 190.720 495.600 191.440 ;
        RECT 1.190 190.040 495.600 190.720 ;
        RECT 1.190 188.040 499.035 190.040 ;
        RECT 4.400 186.640 495.600 188.040 ;
        RECT 1.190 184.640 499.035 186.640 ;
        RECT 1.190 183.960 495.600 184.640 ;
        RECT 4.400 183.240 495.600 183.960 ;
        RECT 4.400 182.560 499.035 183.240 ;
        RECT 1.190 181.240 499.035 182.560 ;
        RECT 1.190 179.880 495.600 181.240 ;
        RECT 4.400 179.840 495.600 179.880 ;
        RECT 4.400 178.480 499.035 179.840 ;
        RECT 1.190 177.840 499.035 178.480 ;
        RECT 1.190 176.440 495.600 177.840 ;
        RECT 1.190 175.800 499.035 176.440 ;
        RECT 4.400 174.440 499.035 175.800 ;
        RECT 4.400 174.400 495.600 174.440 ;
        RECT 1.190 173.040 495.600 174.400 ;
        RECT 1.190 171.720 499.035 173.040 ;
        RECT 4.400 171.040 499.035 171.720 ;
        RECT 4.400 170.320 495.600 171.040 ;
        RECT 1.190 169.640 495.600 170.320 ;
        RECT 1.190 167.640 499.035 169.640 ;
        RECT 4.400 166.240 495.600 167.640 ;
        RECT 1.190 164.240 499.035 166.240 ;
        RECT 1.190 163.560 495.600 164.240 ;
        RECT 4.400 162.840 495.600 163.560 ;
        RECT 4.400 162.160 499.035 162.840 ;
        RECT 1.190 160.840 499.035 162.160 ;
        RECT 1.190 159.480 495.600 160.840 ;
        RECT 4.400 159.440 495.600 159.480 ;
        RECT 4.400 158.080 499.035 159.440 ;
        RECT 1.190 157.440 499.035 158.080 ;
        RECT 1.190 156.040 495.600 157.440 ;
        RECT 1.190 155.400 499.035 156.040 ;
        RECT 4.400 154.040 499.035 155.400 ;
        RECT 4.400 154.000 495.600 154.040 ;
        RECT 1.190 152.640 495.600 154.000 ;
        RECT 1.190 151.320 499.035 152.640 ;
        RECT 4.400 150.640 499.035 151.320 ;
        RECT 4.400 149.920 495.600 150.640 ;
        RECT 1.190 149.240 495.600 149.920 ;
        RECT 1.190 147.240 499.035 149.240 ;
        RECT 4.400 145.840 495.600 147.240 ;
        RECT 1.190 143.840 499.035 145.840 ;
        RECT 1.190 143.160 495.600 143.840 ;
        RECT 4.400 142.440 495.600 143.160 ;
        RECT 4.400 141.760 499.035 142.440 ;
        RECT 1.190 140.440 499.035 141.760 ;
        RECT 1.190 139.080 495.600 140.440 ;
        RECT 4.400 139.040 495.600 139.080 ;
        RECT 4.400 137.680 499.035 139.040 ;
        RECT 1.190 137.040 499.035 137.680 ;
        RECT 1.190 135.640 495.600 137.040 ;
        RECT 1.190 135.000 499.035 135.640 ;
        RECT 4.400 133.640 499.035 135.000 ;
        RECT 4.400 133.600 495.600 133.640 ;
        RECT 1.190 132.240 495.600 133.600 ;
        RECT 1.190 130.920 499.035 132.240 ;
        RECT 4.400 130.240 499.035 130.920 ;
        RECT 4.400 129.520 495.600 130.240 ;
        RECT 1.190 128.840 495.600 129.520 ;
        RECT 1.190 126.840 499.035 128.840 ;
        RECT 4.400 125.440 495.600 126.840 ;
        RECT 1.190 123.440 499.035 125.440 ;
        RECT 1.190 122.760 495.600 123.440 ;
        RECT 4.400 122.040 495.600 122.760 ;
        RECT 4.400 121.360 499.035 122.040 ;
        RECT 1.190 120.040 499.035 121.360 ;
        RECT 1.190 118.680 495.600 120.040 ;
        RECT 4.400 118.640 495.600 118.680 ;
        RECT 4.400 117.280 499.035 118.640 ;
        RECT 1.190 116.640 499.035 117.280 ;
        RECT 1.190 115.240 495.600 116.640 ;
        RECT 1.190 114.600 499.035 115.240 ;
        RECT 4.400 113.240 499.035 114.600 ;
        RECT 4.400 113.200 495.600 113.240 ;
        RECT 1.190 111.840 495.600 113.200 ;
        RECT 1.190 110.520 499.035 111.840 ;
        RECT 4.400 109.840 499.035 110.520 ;
        RECT 4.400 109.120 495.600 109.840 ;
        RECT 1.190 108.440 495.600 109.120 ;
        RECT 1.190 106.440 499.035 108.440 ;
        RECT 4.400 105.040 495.600 106.440 ;
        RECT 1.190 103.040 499.035 105.040 ;
        RECT 1.190 102.360 495.600 103.040 ;
        RECT 4.400 101.640 495.600 102.360 ;
        RECT 4.400 100.960 499.035 101.640 ;
        RECT 1.190 99.640 499.035 100.960 ;
        RECT 1.190 98.280 495.600 99.640 ;
        RECT 4.400 98.240 495.600 98.280 ;
        RECT 4.400 96.880 499.035 98.240 ;
        RECT 1.190 96.240 499.035 96.880 ;
        RECT 1.190 94.840 495.600 96.240 ;
        RECT 1.190 94.200 499.035 94.840 ;
        RECT 4.400 92.840 499.035 94.200 ;
        RECT 4.400 92.800 495.600 92.840 ;
        RECT 1.190 91.440 495.600 92.800 ;
        RECT 1.190 90.120 499.035 91.440 ;
        RECT 4.400 89.440 499.035 90.120 ;
        RECT 4.400 88.720 495.600 89.440 ;
        RECT 1.190 88.040 495.600 88.720 ;
        RECT 1.190 86.040 499.035 88.040 ;
        RECT 4.400 84.640 495.600 86.040 ;
        RECT 1.190 82.640 499.035 84.640 ;
        RECT 1.190 81.960 495.600 82.640 ;
        RECT 4.400 81.240 495.600 81.960 ;
        RECT 4.400 80.560 499.035 81.240 ;
        RECT 1.190 79.240 499.035 80.560 ;
        RECT 1.190 77.880 495.600 79.240 ;
        RECT 4.400 77.840 495.600 77.880 ;
        RECT 4.400 76.480 499.035 77.840 ;
        RECT 1.190 75.840 499.035 76.480 ;
        RECT 1.190 74.440 495.600 75.840 ;
        RECT 1.190 73.800 499.035 74.440 ;
        RECT 4.400 72.440 499.035 73.800 ;
        RECT 4.400 72.400 495.600 72.440 ;
        RECT 1.190 71.040 495.600 72.400 ;
        RECT 1.190 69.720 499.035 71.040 ;
        RECT 4.400 69.040 499.035 69.720 ;
        RECT 4.400 68.320 495.600 69.040 ;
        RECT 1.190 67.640 495.600 68.320 ;
        RECT 1.190 65.640 499.035 67.640 ;
        RECT 4.400 64.240 495.600 65.640 ;
        RECT 1.190 62.240 499.035 64.240 ;
        RECT 1.190 61.560 495.600 62.240 ;
        RECT 4.400 60.840 495.600 61.560 ;
        RECT 4.400 60.160 499.035 60.840 ;
        RECT 1.190 58.840 499.035 60.160 ;
        RECT 1.190 57.480 495.600 58.840 ;
        RECT 4.400 57.440 495.600 57.480 ;
        RECT 4.400 56.080 499.035 57.440 ;
        RECT 1.190 53.400 499.035 56.080 ;
        RECT 4.400 52.000 499.035 53.400 ;
        RECT 1.190 49.320 499.035 52.000 ;
        RECT 4.400 47.920 499.035 49.320 ;
        RECT 1.190 45.240 499.035 47.920 ;
        RECT 4.400 43.840 499.035 45.240 ;
        RECT 1.190 41.160 499.035 43.840 ;
        RECT 4.400 39.760 499.035 41.160 ;
        RECT 1.190 37.080 499.035 39.760 ;
        RECT 4.400 35.680 499.035 37.080 ;
        RECT 1.190 33.000 499.035 35.680 ;
        RECT 4.400 31.600 499.035 33.000 ;
        RECT 1.190 28.920 499.035 31.600 ;
        RECT 4.400 27.520 499.035 28.920 ;
        RECT 1.190 24.840 499.035 27.520 ;
        RECT 4.400 23.440 499.035 24.840 ;
        RECT 1.190 20.760 499.035 23.440 ;
        RECT 4.400 19.360 499.035 20.760 ;
        RECT 1.190 16.680 499.035 19.360 ;
        RECT 4.400 15.280 499.035 16.680 ;
        RECT 1.190 12.600 499.035 15.280 ;
        RECT 4.400 11.200 499.035 12.600 ;
        RECT 1.190 8.520 499.035 11.200 ;
        RECT 4.400 7.655 499.035 8.520 ;
      LAYER met4 ;
        RECT 1.215 11.735 20.640 780.465 ;
        RECT 23.040 11.735 97.440 780.465 ;
        RECT 99.840 11.735 174.240 780.465 ;
        RECT 176.640 11.735 251.040 780.465 ;
        RECT 253.440 11.735 327.840 780.465 ;
        RECT 330.240 11.735 404.640 780.465 ;
        RECT 407.040 11.735 481.440 780.465 ;
        RECT 483.840 11.735 494.665 780.465 ;
  END
END ExperiarCore
END LIBRARY

