magic
tech sky130A
magscale 1 2
timestamp 1653062883
<< obsli1 >>
rect 1104 2159 118864 37553
<< obsm1 >>
rect 382 1368 118864 37584
<< metal2 >>
rect 2042 39200 2098 40000
rect 6090 39200 6146 40000
rect 10230 39200 10286 40000
rect 14370 39200 14426 40000
rect 18510 39200 18566 40000
rect 22650 39200 22706 40000
rect 26790 39200 26846 40000
rect 30930 39200 30986 40000
rect 35070 39200 35126 40000
rect 39210 39200 39266 40000
rect 43350 39200 43406 40000
rect 47490 39200 47546 40000
rect 51630 39200 51686 40000
rect 55770 39200 55826 40000
rect 59910 39200 59966 40000
rect 64050 39200 64106 40000
rect 68190 39200 68246 40000
rect 72330 39200 72386 40000
rect 76470 39200 76526 40000
rect 80610 39200 80666 40000
rect 84750 39200 84806 40000
rect 88890 39200 88946 40000
rect 93030 39200 93086 40000
rect 97170 39200 97226 40000
rect 101310 39200 101366 40000
rect 105450 39200 105506 40000
rect 109590 39200 109646 40000
rect 113730 39200 113786 40000
rect 117870 39200 117926 40000
rect 386 0 442 800
rect 1122 0 1178 800
rect 1950 0 2006 800
rect 2778 0 2834 800
rect 3514 0 3570 800
rect 4342 0 4398 800
rect 5170 0 5226 800
rect 5906 0 5962 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8298 0 8354 800
rect 9126 0 9182 800
rect 9954 0 10010 800
rect 10782 0 10838 800
rect 11518 0 11574 800
rect 12346 0 12402 800
rect 13174 0 13230 800
rect 13910 0 13966 800
rect 14738 0 14794 800
rect 15566 0 15622 800
rect 16302 0 16358 800
rect 17130 0 17186 800
rect 17958 0 18014 800
rect 18694 0 18750 800
rect 19522 0 19578 800
rect 20350 0 20406 800
rect 21178 0 21234 800
rect 21914 0 21970 800
rect 22742 0 22798 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 25134 0 25190 800
rect 25962 0 26018 800
rect 26698 0 26754 800
rect 27526 0 27582 800
rect 28354 0 28410 800
rect 29090 0 29146 800
rect 29918 0 29974 800
rect 30746 0 30802 800
rect 31574 0 31630 800
rect 32310 0 32366 800
rect 33138 0 33194 800
rect 33966 0 34022 800
rect 34702 0 34758 800
rect 35530 0 35586 800
rect 36358 0 36414 800
rect 37094 0 37150 800
rect 37922 0 37978 800
rect 38750 0 38806 800
rect 39486 0 39542 800
rect 40314 0 40370 800
rect 41142 0 41198 800
rect 41970 0 42026 800
rect 42706 0 42762 800
rect 43534 0 43590 800
rect 44362 0 44418 800
rect 45098 0 45154 800
rect 45926 0 45982 800
rect 46754 0 46810 800
rect 47490 0 47546 800
rect 48318 0 48374 800
rect 49146 0 49202 800
rect 49882 0 49938 800
rect 50710 0 50766 800
rect 51538 0 51594 800
rect 52366 0 52422 800
rect 53102 0 53158 800
rect 53930 0 53986 800
rect 54758 0 54814 800
rect 55494 0 55550 800
rect 56322 0 56378 800
rect 57150 0 57206 800
rect 57886 0 57942 800
rect 58714 0 58770 800
rect 59542 0 59598 800
rect 60370 0 60426 800
rect 61106 0 61162 800
rect 61934 0 61990 800
rect 62762 0 62818 800
rect 63498 0 63554 800
rect 64326 0 64382 800
rect 65154 0 65210 800
rect 65890 0 65946 800
rect 66718 0 66774 800
rect 67546 0 67602 800
rect 68282 0 68338 800
rect 69110 0 69166 800
rect 69938 0 69994 800
rect 70766 0 70822 800
rect 71502 0 71558 800
rect 72330 0 72386 800
rect 73158 0 73214 800
rect 73894 0 73950 800
rect 74722 0 74778 800
rect 75550 0 75606 800
rect 76286 0 76342 800
rect 77114 0 77170 800
rect 77942 0 77998 800
rect 78678 0 78734 800
rect 79506 0 79562 800
rect 80334 0 80390 800
rect 81162 0 81218 800
rect 81898 0 81954 800
rect 82726 0 82782 800
rect 83554 0 83610 800
rect 84290 0 84346 800
rect 85118 0 85174 800
rect 85946 0 86002 800
rect 86682 0 86738 800
rect 87510 0 87566 800
rect 88338 0 88394 800
rect 89074 0 89130 800
rect 89902 0 89958 800
rect 90730 0 90786 800
rect 91558 0 91614 800
rect 92294 0 92350 800
rect 93122 0 93178 800
rect 93950 0 94006 800
rect 94686 0 94742 800
rect 95514 0 95570 800
rect 96342 0 96398 800
rect 97078 0 97134 800
rect 97906 0 97962 800
rect 98734 0 98790 800
rect 99470 0 99526 800
rect 100298 0 100354 800
rect 101126 0 101182 800
rect 101954 0 102010 800
rect 102690 0 102746 800
rect 103518 0 103574 800
rect 104346 0 104402 800
rect 105082 0 105138 800
rect 105910 0 105966 800
rect 106738 0 106794 800
rect 107474 0 107530 800
rect 108302 0 108358 800
rect 109130 0 109186 800
rect 109866 0 109922 800
rect 110694 0 110750 800
rect 111522 0 111578 800
rect 112350 0 112406 800
rect 113086 0 113142 800
rect 113914 0 113970 800
rect 114742 0 114798 800
rect 115478 0 115534 800
rect 116306 0 116362 800
rect 117134 0 117190 800
rect 117870 0 117926 800
rect 118698 0 118754 800
rect 119526 0 119582 800
<< obsm2 >>
rect 388 39144 1986 39273
rect 2154 39144 6034 39273
rect 6202 39144 10174 39273
rect 10342 39144 14314 39273
rect 14482 39144 18454 39273
rect 18622 39144 22594 39273
rect 22762 39144 26734 39273
rect 26902 39144 30874 39273
rect 31042 39144 35014 39273
rect 35182 39144 39154 39273
rect 39322 39144 43294 39273
rect 43462 39144 47434 39273
rect 47602 39144 51574 39273
rect 51742 39144 55714 39273
rect 55882 39144 59854 39273
rect 60022 39144 63994 39273
rect 64162 39144 68134 39273
rect 68302 39144 72274 39273
rect 72442 39144 76414 39273
rect 76582 39144 80554 39273
rect 80722 39144 84694 39273
rect 84862 39144 88834 39273
rect 89002 39144 92974 39273
rect 93142 39144 97114 39273
rect 97282 39144 101254 39273
rect 101422 39144 105394 39273
rect 105562 39144 109534 39273
rect 109702 39144 113674 39273
rect 113842 39144 117814 39273
rect 117982 39144 118202 39273
rect 388 856 118202 39144
rect 498 711 1066 856
rect 1234 711 1894 856
rect 2062 711 2722 856
rect 2890 711 3458 856
rect 3626 711 4286 856
rect 4454 711 5114 856
rect 5282 711 5850 856
rect 6018 711 6678 856
rect 6846 711 7506 856
rect 7674 711 8242 856
rect 8410 711 9070 856
rect 9238 711 9898 856
rect 10066 711 10726 856
rect 10894 711 11462 856
rect 11630 711 12290 856
rect 12458 711 13118 856
rect 13286 711 13854 856
rect 14022 711 14682 856
rect 14850 711 15510 856
rect 15678 711 16246 856
rect 16414 711 17074 856
rect 17242 711 17902 856
rect 18070 711 18638 856
rect 18806 711 19466 856
rect 19634 711 20294 856
rect 20462 711 21122 856
rect 21290 711 21858 856
rect 22026 711 22686 856
rect 22854 711 23514 856
rect 23682 711 24250 856
rect 24418 711 25078 856
rect 25246 711 25906 856
rect 26074 711 26642 856
rect 26810 711 27470 856
rect 27638 711 28298 856
rect 28466 711 29034 856
rect 29202 711 29862 856
rect 30030 711 30690 856
rect 30858 711 31518 856
rect 31686 711 32254 856
rect 32422 711 33082 856
rect 33250 711 33910 856
rect 34078 711 34646 856
rect 34814 711 35474 856
rect 35642 711 36302 856
rect 36470 711 37038 856
rect 37206 711 37866 856
rect 38034 711 38694 856
rect 38862 711 39430 856
rect 39598 711 40258 856
rect 40426 711 41086 856
rect 41254 711 41914 856
rect 42082 711 42650 856
rect 42818 711 43478 856
rect 43646 711 44306 856
rect 44474 711 45042 856
rect 45210 711 45870 856
rect 46038 711 46698 856
rect 46866 711 47434 856
rect 47602 711 48262 856
rect 48430 711 49090 856
rect 49258 711 49826 856
rect 49994 711 50654 856
rect 50822 711 51482 856
rect 51650 711 52310 856
rect 52478 711 53046 856
rect 53214 711 53874 856
rect 54042 711 54702 856
rect 54870 711 55438 856
rect 55606 711 56266 856
rect 56434 711 57094 856
rect 57262 711 57830 856
rect 57998 711 58658 856
rect 58826 711 59486 856
rect 59654 711 60314 856
rect 60482 711 61050 856
rect 61218 711 61878 856
rect 62046 711 62706 856
rect 62874 711 63442 856
rect 63610 711 64270 856
rect 64438 711 65098 856
rect 65266 711 65834 856
rect 66002 711 66662 856
rect 66830 711 67490 856
rect 67658 711 68226 856
rect 68394 711 69054 856
rect 69222 711 69882 856
rect 70050 711 70710 856
rect 70878 711 71446 856
rect 71614 711 72274 856
rect 72442 711 73102 856
rect 73270 711 73838 856
rect 74006 711 74666 856
rect 74834 711 75494 856
rect 75662 711 76230 856
rect 76398 711 77058 856
rect 77226 711 77886 856
rect 78054 711 78622 856
rect 78790 711 79450 856
rect 79618 711 80278 856
rect 80446 711 81106 856
rect 81274 711 81842 856
rect 82010 711 82670 856
rect 82838 711 83498 856
rect 83666 711 84234 856
rect 84402 711 85062 856
rect 85230 711 85890 856
rect 86058 711 86626 856
rect 86794 711 87454 856
rect 87622 711 88282 856
rect 88450 711 89018 856
rect 89186 711 89846 856
rect 90014 711 90674 856
rect 90842 711 91502 856
rect 91670 711 92238 856
rect 92406 711 93066 856
rect 93234 711 93894 856
rect 94062 711 94630 856
rect 94798 711 95458 856
rect 95626 711 96286 856
rect 96454 711 97022 856
rect 97190 711 97850 856
rect 98018 711 98678 856
rect 98846 711 99414 856
rect 99582 711 100242 856
rect 100410 711 101070 856
rect 101238 711 101898 856
rect 102066 711 102634 856
rect 102802 711 103462 856
rect 103630 711 104290 856
rect 104458 711 105026 856
rect 105194 711 105854 856
rect 106022 711 106682 856
rect 106850 711 107418 856
rect 107586 711 108246 856
rect 108414 711 109074 856
rect 109242 711 109810 856
rect 109978 711 110638 856
rect 110806 711 111466 856
rect 111634 711 112294 856
rect 112462 711 113030 856
rect 113198 711 113858 856
rect 114026 711 114686 856
rect 114854 711 115422 856
rect 115590 711 116250 856
rect 116418 711 117078 856
rect 117246 711 117814 856
rect 117982 711 118202 856
<< metal3 >>
rect 0 39040 800 39160
rect 119200 39176 120000 39296
rect 119200 37816 120000 37936
rect 0 37408 800 37528
rect 119200 36320 120000 36440
rect 0 35776 800 35896
rect 119200 34960 120000 35080
rect 0 34144 800 34264
rect 119200 33464 120000 33584
rect 0 32376 800 32496
rect 119200 32104 120000 32224
rect 0 30744 800 30864
rect 119200 30608 120000 30728
rect 0 29112 800 29232
rect 119200 29248 120000 29368
rect 119200 27752 120000 27872
rect 0 27480 800 27600
rect 119200 26392 120000 26512
rect 0 25712 800 25832
rect 119200 24896 120000 25016
rect 0 24080 800 24200
rect 119200 23536 120000 23656
rect 0 22448 800 22568
rect 119200 22040 120000 22160
rect 0 20816 800 20936
rect 119200 20680 120000 20800
rect 0 19048 800 19168
rect 119200 19184 120000 19304
rect 119200 17824 120000 17944
rect 0 17416 800 17536
rect 119200 16328 120000 16448
rect 0 15784 800 15904
rect 119200 14968 120000 15088
rect 0 14152 800 14272
rect 119200 13472 120000 13592
rect 0 12384 800 12504
rect 119200 12112 120000 12232
rect 0 10752 800 10872
rect 119200 10616 120000 10736
rect 0 9120 800 9240
rect 119200 9256 120000 9376
rect 119200 7760 120000 7880
rect 0 7488 800 7608
rect 119200 6400 120000 6520
rect 0 5720 800 5840
rect 119200 4904 120000 5024
rect 0 4088 800 4208
rect 119200 3544 120000 3664
rect 0 2456 800 2576
rect 119200 2048 120000 2168
rect 0 824 800 944
rect 119200 688 120000 808
<< obsm3 >>
rect 800 39240 119120 39269
rect 880 39096 119120 39240
rect 880 38960 119200 39096
rect 800 38016 119200 38960
rect 800 37736 119120 38016
rect 800 37608 119200 37736
rect 880 37328 119200 37608
rect 800 36520 119200 37328
rect 800 36240 119120 36520
rect 800 35976 119200 36240
rect 880 35696 119200 35976
rect 800 35160 119200 35696
rect 800 34880 119120 35160
rect 800 34344 119200 34880
rect 880 34064 119200 34344
rect 800 33664 119200 34064
rect 800 33384 119120 33664
rect 800 32576 119200 33384
rect 880 32304 119200 32576
rect 880 32296 119120 32304
rect 800 32024 119120 32296
rect 800 30944 119200 32024
rect 880 30808 119200 30944
rect 880 30664 119120 30808
rect 800 30528 119120 30664
rect 800 29448 119200 30528
rect 800 29312 119120 29448
rect 880 29168 119120 29312
rect 880 29032 119200 29168
rect 800 27952 119200 29032
rect 800 27680 119120 27952
rect 880 27672 119120 27680
rect 880 27400 119200 27672
rect 800 26592 119200 27400
rect 800 26312 119120 26592
rect 800 25912 119200 26312
rect 880 25632 119200 25912
rect 800 25096 119200 25632
rect 800 24816 119120 25096
rect 800 24280 119200 24816
rect 880 24000 119200 24280
rect 800 23736 119200 24000
rect 800 23456 119120 23736
rect 800 22648 119200 23456
rect 880 22368 119200 22648
rect 800 22240 119200 22368
rect 800 21960 119120 22240
rect 800 21016 119200 21960
rect 880 20880 119200 21016
rect 880 20736 119120 20880
rect 800 20600 119120 20736
rect 800 19384 119200 20600
rect 800 19248 119120 19384
rect 880 19104 119120 19248
rect 880 18968 119200 19104
rect 800 18024 119200 18968
rect 800 17744 119120 18024
rect 800 17616 119200 17744
rect 880 17336 119200 17616
rect 800 16528 119200 17336
rect 800 16248 119120 16528
rect 800 15984 119200 16248
rect 880 15704 119200 15984
rect 800 15168 119200 15704
rect 800 14888 119120 15168
rect 800 14352 119200 14888
rect 880 14072 119200 14352
rect 800 13672 119200 14072
rect 800 13392 119120 13672
rect 800 12584 119200 13392
rect 880 12312 119200 12584
rect 880 12304 119120 12312
rect 800 12032 119120 12304
rect 800 10952 119200 12032
rect 880 10816 119200 10952
rect 880 10672 119120 10816
rect 800 10536 119120 10672
rect 800 9456 119200 10536
rect 800 9320 119120 9456
rect 880 9176 119120 9320
rect 880 9040 119200 9176
rect 800 7960 119200 9040
rect 800 7688 119120 7960
rect 880 7680 119120 7688
rect 880 7408 119200 7680
rect 800 6600 119200 7408
rect 800 6320 119120 6600
rect 800 5920 119200 6320
rect 880 5640 119200 5920
rect 800 5104 119200 5640
rect 800 4824 119120 5104
rect 800 4288 119200 4824
rect 880 4008 119200 4288
rect 800 3744 119200 4008
rect 800 3464 119120 3744
rect 800 2656 119200 3464
rect 880 2376 119200 2656
rect 800 2248 119200 2376
rect 800 1968 119120 2248
rect 800 1024 119200 1968
rect 880 888 119200 1024
rect 880 744 119120 888
rect 800 715 119120 744
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
rect 65648 2128 65968 37584
rect 81008 2128 81328 37584
rect 96368 2128 96688 37584
rect 111728 2128 112048 37584
<< labels >>
rlabel metal2 s 2042 39200 2098 40000 6 flash_csb
port 1 nsew signal output
rlabel metal2 s 6090 39200 6146 40000 6 flash_io0_read
port 2 nsew signal input
rlabel metal2 s 10230 39200 10286 40000 6 flash_io0_we
port 3 nsew signal output
rlabel metal2 s 14370 39200 14426 40000 6 flash_io0_write
port 4 nsew signal output
rlabel metal2 s 18510 39200 18566 40000 6 flash_io1_read
port 5 nsew signal input
rlabel metal2 s 22650 39200 22706 40000 6 flash_io1_we
port 6 nsew signal output
rlabel metal2 s 26790 39200 26846 40000 6 flash_io1_write
port 7 nsew signal output
rlabel metal2 s 30930 39200 30986 40000 6 flash_sck
port 8 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 sram_addr0[0]
port 9 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 sram_addr0[1]
port 10 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 sram_addr0[2]
port 11 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 sram_addr0[3]
port 12 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 sram_addr0[4]
port 13 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 sram_addr0[5]
port 14 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 sram_addr0[6]
port 15 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 sram_addr0[7]
port 16 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 sram_addr0[8]
port 17 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 sram_addr1[0]
port 18 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 sram_addr1[1]
port 19 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 sram_addr1[2]
port 20 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 sram_addr1[3]
port 21 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 sram_addr1[4]
port 22 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 sram_addr1[5]
port 23 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 sram_addr1[6]
port 24 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 sram_addr1[7]
port 25 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 sram_addr1[8]
port 26 nsew signal output
rlabel metal2 s 386 0 442 800 6 sram_clk0
port 27 nsew signal output
rlabel metal2 s 1122 0 1178 800 6 sram_clk1
port 28 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 sram_csb0
port 29 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 sram_csb1
port 30 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 sram_din0[0]
port 31 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 sram_din0[10]
port 32 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 sram_din0[11]
port 33 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 sram_din0[12]
port 34 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 sram_din0[13]
port 35 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 sram_din0[14]
port 36 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 sram_din0[15]
port 37 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 sram_din0[16]
port 38 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 sram_din0[17]
port 39 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 sram_din0[18]
port 40 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 sram_din0[19]
port 41 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 sram_din0[1]
port 42 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 sram_din0[20]
port 43 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 sram_din0[21]
port 44 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 sram_din0[22]
port 45 nsew signal output
rlabel metal2 s 77114 0 77170 800 6 sram_din0[23]
port 46 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 sram_din0[24]
port 47 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 sram_din0[25]
port 48 nsew signal output
rlabel metal2 s 84290 0 84346 800 6 sram_din0[26]
port 49 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 sram_din0[27]
port 50 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 sram_din0[28]
port 51 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 sram_din0[29]
port 52 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 sram_din0[2]
port 53 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 sram_din0[30]
port 54 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 sram_din0[31]
port 55 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 sram_din0[3]
port 56 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 sram_din0[4]
port 57 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 sram_din0[5]
port 58 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 sram_din0[6]
port 59 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 sram_din0[7]
port 60 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 sram_din0[8]
port 61 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 sram_din0[9]
port 62 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 sram_dout0[0]
port 63 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 sram_dout0[10]
port 64 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 sram_dout0[11]
port 65 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 sram_dout0[12]
port 66 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 sram_dout0[13]
port 67 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 sram_dout0[14]
port 68 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 sram_dout0[15]
port 69 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 sram_dout0[16]
port 70 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 sram_dout0[17]
port 71 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 sram_dout0[18]
port 72 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 sram_dout0[19]
port 73 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 sram_dout0[1]
port 74 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 sram_dout0[20]
port 75 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 sram_dout0[21]
port 76 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 sram_dout0[22]
port 77 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 sram_dout0[23]
port 78 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 sram_dout0[24]
port 79 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 sram_dout0[25]
port 80 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 sram_dout0[26]
port 81 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 sram_dout0[27]
port 82 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 sram_dout0[28]
port 83 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 sram_dout0[29]
port 84 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 sram_dout0[2]
port 85 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 sram_dout0[30]
port 86 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 sram_dout0[31]
port 87 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 sram_dout0[3]
port 88 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 sram_dout0[4]
port 89 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 sram_dout0[5]
port 90 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 sram_dout0[6]
port 91 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 sram_dout0[7]
port 92 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 sram_dout0[8]
port 93 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 sram_dout0[9]
port 94 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 sram_dout1[0]
port 95 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 sram_dout1[10]
port 96 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 sram_dout1[11]
port 97 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 sram_dout1[12]
port 98 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 sram_dout1[13]
port 99 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 sram_dout1[14]
port 100 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 sram_dout1[15]
port 101 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 sram_dout1[16]
port 102 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 sram_dout1[17]
port 103 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 sram_dout1[18]
port 104 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 sram_dout1[19]
port 105 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 sram_dout1[1]
port 106 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 sram_dout1[20]
port 107 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 sram_dout1[21]
port 108 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 sram_dout1[22]
port 109 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 sram_dout1[23]
port 110 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 sram_dout1[24]
port 111 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 sram_dout1[25]
port 112 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 sram_dout1[26]
port 113 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 sram_dout1[27]
port 114 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 sram_dout1[28]
port 115 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 sram_dout1[29]
port 116 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 sram_dout1[2]
port 117 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 sram_dout1[30]
port 118 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 sram_dout1[31]
port 119 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 sram_dout1[3]
port 120 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 sram_dout1[4]
port 121 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 sram_dout1[5]
port 122 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 sram_dout1[6]
port 123 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 sram_dout1[7]
port 124 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 sram_dout1[8]
port 125 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 sram_dout1[9]
port 126 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 sram_web0
port 127 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 sram_wmask0[0]
port 128 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 sram_wmask0[1]
port 129 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 sram_wmask0[2]
port 130 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 sram_wmask0[3]
port 131 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 37584 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 133 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 133 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 37584 6 vssd1
port 133 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 37584 6 vssd1
port 133 nsew ground bidirectional
rlabel metal3 s 119200 688 120000 808 6 wb_ack_o
port 134 nsew signal output
rlabel metal2 s 98734 0 98790 800 6 wb_adr_i[0]
port 135 nsew signal input
rlabel metal3 s 119200 17824 120000 17944 6 wb_adr_i[10]
port 136 nsew signal input
rlabel metal3 s 119200 20680 120000 20800 6 wb_adr_i[11]
port 137 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_adr_i[12]
port 138 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 wb_adr_i[13]
port 139 nsew signal input
rlabel metal2 s 76470 39200 76526 40000 6 wb_adr_i[14]
port 140 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wb_adr_i[15]
port 141 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 wb_adr_i[16]
port 142 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 wb_adr_i[17]
port 143 nsew signal input
rlabel metal3 s 119200 29248 120000 29368 6 wb_adr_i[18]
port 144 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 wb_adr_i[19]
port 145 nsew signal input
rlabel metal3 s 119200 9256 120000 9376 6 wb_adr_i[1]
port 146 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 wb_adr_i[20]
port 147 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 wb_adr_i[21]
port 148 nsew signal input
rlabel metal2 s 93030 39200 93086 40000 6 wb_adr_i[22]
port 149 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 wb_adr_i[23]
port 150 nsew signal input
rlabel metal2 s 51630 39200 51686 40000 6 wb_adr_i[2]
port 151 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 wb_adr_i[3]
port 152 nsew signal input
rlabel metal3 s 119200 12112 120000 12232 6 wb_adr_i[4]
port 153 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 wb_adr_i[5]
port 154 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 wb_adr_i[6]
port 155 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 wb_adr_i[7]
port 156 nsew signal input
rlabel metal3 s 119200 14968 120000 15088 6 wb_adr_i[8]
port 157 nsew signal input
rlabel metal2 s 68190 39200 68246 40000 6 wb_adr_i[9]
port 158 nsew signal input
rlabel metal3 s 0 824 800 944 6 wb_clk_i
port 159 nsew signal input
rlabel metal3 s 119200 2048 120000 2168 6 wb_cyc_i
port 160 nsew signal input
rlabel metal2 s 43350 39200 43406 40000 6 wb_data_i[0]
port 161 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 wb_data_i[10]
port 162 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 wb_data_i[11]
port 163 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 wb_data_i[12]
port 164 nsew signal input
rlabel metal3 s 119200 24896 120000 25016 6 wb_data_i[13]
port 165 nsew signal input
rlabel metal2 s 80610 39200 80666 40000 6 wb_data_i[14]
port 166 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 wb_data_i[15]
port 167 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 wb_data_i[16]
port 168 nsew signal input
rlabel metal3 s 119200 27752 120000 27872 6 wb_data_i[17]
port 169 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 wb_data_i[18]
port 170 nsew signal input
rlabel metal3 s 119200 30608 120000 30728 6 wb_data_i[19]
port 171 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 wb_data_i[1]
port 172 nsew signal input
rlabel metal2 s 88890 39200 88946 40000 6 wb_data_i[20]
port 173 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 wb_data_i[21]
port 174 nsew signal input
rlabel metal2 s 97170 39200 97226 40000 6 wb_data_i[22]
port 175 nsew signal input
rlabel metal3 s 119200 32104 120000 32224 6 wb_data_i[23]
port 176 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 wb_data_i[24]
port 177 nsew signal input
rlabel metal2 s 101310 39200 101366 40000 6 wb_data_i[25]
port 178 nsew signal input
rlabel metal2 s 105450 39200 105506 40000 6 wb_data_i[26]
port 179 nsew signal input
rlabel metal3 s 119200 36320 120000 36440 6 wb_data_i[27]
port 180 nsew signal input
rlabel metal3 s 119200 37816 120000 37936 6 wb_data_i[28]
port 181 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 wb_data_i[29]
port 182 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 wb_data_i[2]
port 183 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 wb_data_i[30]
port 184 nsew signal input
rlabel metal2 s 113730 39200 113786 40000 6 wb_data_i[31]
port 185 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 wb_data_i[3]
port 186 nsew signal input
rlabel metal3 s 119200 13472 120000 13592 6 wb_data_i[4]
port 187 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 wb_data_i[5]
port 188 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wb_data_i[6]
port 189 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 wb_data_i[7]
port 190 nsew signal input
rlabel metal3 s 119200 16328 120000 16448 6 wb_data_i[8]
port 191 nsew signal input
rlabel metal2 s 72330 39200 72386 40000 6 wb_data_i[9]
port 192 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 wb_data_o[0]
port 193 nsew signal output
rlabel metal3 s 119200 19184 120000 19304 6 wb_data_o[10]
port 194 nsew signal output
rlabel metal3 s 119200 22040 120000 22160 6 wb_data_o[11]
port 195 nsew signal output
rlabel metal3 s 119200 23536 120000 23656 6 wb_data_o[12]
port 196 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 wb_data_o[13]
port 197 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 wb_data_o[14]
port 198 nsew signal output
rlabel metal3 s 119200 26392 120000 26512 6 wb_data_o[15]
port 199 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 wb_data_o[16]
port 200 nsew signal output
rlabel metal2 s 84750 39200 84806 40000 6 wb_data_o[17]
port 201 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 wb_data_o[18]
port 202 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 wb_data_o[19]
port 203 nsew signal output
rlabel metal2 s 47490 39200 47546 40000 6 wb_data_o[1]
port 204 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 wb_data_o[20]
port 205 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 wb_data_o[21]
port 206 nsew signal output
rlabel metal2 s 114742 0 114798 800 6 wb_data_o[22]
port 207 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 wb_data_o[23]
port 208 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 wb_data_o[24]
port 209 nsew signal output
rlabel metal3 s 119200 33464 120000 33584 6 wb_data_o[25]
port 210 nsew signal output
rlabel metal3 s 119200 34960 120000 35080 6 wb_data_o[26]
port 211 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 wb_data_o[27]
port 212 nsew signal output
rlabel metal3 s 119200 39176 120000 39296 6 wb_data_o[28]
port 213 nsew signal output
rlabel metal3 s 0 39040 800 39160 6 wb_data_o[29]
port 214 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 wb_data_o[2]
port 215 nsew signal output
rlabel metal2 s 109590 39200 109646 40000 6 wb_data_o[30]
port 216 nsew signal output
rlabel metal2 s 117870 39200 117926 40000 6 wb_data_o[31]
port 217 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 wb_data_o[3]
port 218 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 wb_data_o[4]
port 219 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 wb_data_o[5]
port 220 nsew signal output
rlabel metal2 s 55770 39200 55826 40000 6 wb_data_o[6]
port 221 nsew signal output
rlabel metal2 s 59910 39200 59966 40000 6 wb_data_o[7]
port 222 nsew signal output
rlabel metal2 s 64050 39200 64106 40000 6 wb_data_o[8]
port 223 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 wb_data_o[9]
port 224 nsew signal output
rlabel metal2 s 35070 39200 35126 40000 6 wb_error_o
port 225 nsew signal output
rlabel metal3 s 119200 3544 120000 3664 6 wb_rst_i
port 226 nsew signal input
rlabel metal3 s 119200 7760 120000 7880 6 wb_sel_i[0]
port 227 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 wb_sel_i[1]
port 228 nsew signal input
rlabel metal3 s 119200 10616 120000 10736 6 wb_sel_i[2]
port 229 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 wb_sel_i[3]
port 230 nsew signal input
rlabel metal3 s 119200 4904 120000 5024 6 wb_stall_o
port 231 nsew signal output
rlabel metal2 s 39210 39200 39266 40000 6 wb_stb_i
port 232 nsew signal input
rlabel metal3 s 119200 6400 120000 6520 6 wb_we_i
port 233 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1868304
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Flash/runs/Flash/results/signoff/Flash.magic.gds
string GDS_START 198456
<< end >>

