VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO WishboneInterconnect
  CLASS BLOCK ;
  FOREIGN WishboneInterconnect ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 1000.000 ;
  PIN master0_wb_ack_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END master0_wb_ack_i
  PIN master0_wb_adr_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END master0_wb_adr_o[0]
  PIN master0_wb_adr_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END master0_wb_adr_o[10]
  PIN master0_wb_adr_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END master0_wb_adr_o[11]
  PIN master0_wb_adr_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END master0_wb_adr_o[12]
  PIN master0_wb_adr_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END master0_wb_adr_o[13]
  PIN master0_wb_adr_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END master0_wb_adr_o[14]
  PIN master0_wb_adr_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END master0_wb_adr_o[15]
  PIN master0_wb_adr_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END master0_wb_adr_o[16]
  PIN master0_wb_adr_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END master0_wb_adr_o[17]
  PIN master0_wb_adr_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END master0_wb_adr_o[18]
  PIN master0_wb_adr_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END master0_wb_adr_o[19]
  PIN master0_wb_adr_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END master0_wb_adr_o[1]
  PIN master0_wb_adr_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END master0_wb_adr_o[20]
  PIN master0_wb_adr_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END master0_wb_adr_o[21]
  PIN master0_wb_adr_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END master0_wb_adr_o[22]
  PIN master0_wb_adr_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END master0_wb_adr_o[23]
  PIN master0_wb_adr_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END master0_wb_adr_o[24]
  PIN master0_wb_adr_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END master0_wb_adr_o[25]
  PIN master0_wb_adr_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END master0_wb_adr_o[26]
  PIN master0_wb_adr_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END master0_wb_adr_o[27]
  PIN master0_wb_adr_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END master0_wb_adr_o[2]
  PIN master0_wb_adr_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END master0_wb_adr_o[3]
  PIN master0_wb_adr_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END master0_wb_adr_o[4]
  PIN master0_wb_adr_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END master0_wb_adr_o[5]
  PIN master0_wb_adr_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END master0_wb_adr_o[6]
  PIN master0_wb_adr_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END master0_wb_adr_o[7]
  PIN master0_wb_adr_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END master0_wb_adr_o[8]
  PIN master0_wb_adr_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END master0_wb_adr_o[9]
  PIN master0_wb_cyc_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END master0_wb_cyc_o
  PIN master0_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END master0_wb_data_i[0]
  PIN master0_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END master0_wb_data_i[10]
  PIN master0_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END master0_wb_data_i[11]
  PIN master0_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END master0_wb_data_i[12]
  PIN master0_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END master0_wb_data_i[13]
  PIN master0_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END master0_wb_data_i[14]
  PIN master0_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END master0_wb_data_i[15]
  PIN master0_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END master0_wb_data_i[16]
  PIN master0_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END master0_wb_data_i[17]
  PIN master0_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END master0_wb_data_i[18]
  PIN master0_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END master0_wb_data_i[19]
  PIN master0_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END master0_wb_data_i[1]
  PIN master0_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END master0_wb_data_i[20]
  PIN master0_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END master0_wb_data_i[21]
  PIN master0_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END master0_wb_data_i[22]
  PIN master0_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END master0_wb_data_i[23]
  PIN master0_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END master0_wb_data_i[24]
  PIN master0_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END master0_wb_data_i[25]
  PIN master0_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END master0_wb_data_i[26]
  PIN master0_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END master0_wb_data_i[27]
  PIN master0_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END master0_wb_data_i[28]
  PIN master0_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END master0_wb_data_i[29]
  PIN master0_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END master0_wb_data_i[2]
  PIN master0_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END master0_wb_data_i[30]
  PIN master0_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END master0_wb_data_i[31]
  PIN master0_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END master0_wb_data_i[3]
  PIN master0_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END master0_wb_data_i[4]
  PIN master0_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END master0_wb_data_i[5]
  PIN master0_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END master0_wb_data_i[6]
  PIN master0_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END master0_wb_data_i[7]
  PIN master0_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END master0_wb_data_i[8]
  PIN master0_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END master0_wb_data_i[9]
  PIN master0_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END master0_wb_data_o[0]
  PIN master0_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END master0_wb_data_o[10]
  PIN master0_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END master0_wb_data_o[11]
  PIN master0_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END master0_wb_data_o[12]
  PIN master0_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END master0_wb_data_o[13]
  PIN master0_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END master0_wb_data_o[14]
  PIN master0_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END master0_wb_data_o[15]
  PIN master0_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END master0_wb_data_o[16]
  PIN master0_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END master0_wb_data_o[17]
  PIN master0_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END master0_wb_data_o[18]
  PIN master0_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END master0_wb_data_o[19]
  PIN master0_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END master0_wb_data_o[1]
  PIN master0_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END master0_wb_data_o[20]
  PIN master0_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END master0_wb_data_o[21]
  PIN master0_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END master0_wb_data_o[22]
  PIN master0_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END master0_wb_data_o[23]
  PIN master0_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END master0_wb_data_o[24]
  PIN master0_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END master0_wb_data_o[25]
  PIN master0_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END master0_wb_data_o[26]
  PIN master0_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END master0_wb_data_o[27]
  PIN master0_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END master0_wb_data_o[28]
  PIN master0_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END master0_wb_data_o[29]
  PIN master0_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END master0_wb_data_o[2]
  PIN master0_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END master0_wb_data_o[30]
  PIN master0_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END master0_wb_data_o[31]
  PIN master0_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END master0_wb_data_o[3]
  PIN master0_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END master0_wb_data_o[4]
  PIN master0_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END master0_wb_data_o[5]
  PIN master0_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END master0_wb_data_o[6]
  PIN master0_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END master0_wb_data_o[7]
  PIN master0_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END master0_wb_data_o[8]
  PIN master0_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END master0_wb_data_o[9]
  PIN master0_wb_error_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END master0_wb_error_i
  PIN master0_wb_sel_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END master0_wb_sel_o[0]
  PIN master0_wb_sel_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END master0_wb_sel_o[1]
  PIN master0_wb_sel_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END master0_wb_sel_o[2]
  PIN master0_wb_sel_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END master0_wb_sel_o[3]
  PIN master0_wb_stall_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END master0_wb_stall_i
  PIN master0_wb_stb_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END master0_wb_stb_o
  PIN master0_wb_we_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END master0_wb_we_o
  PIN master1_wb_ack_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END master1_wb_ack_i
  PIN master1_wb_adr_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END master1_wb_adr_o[0]
  PIN master1_wb_adr_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 600.480 4.000 601.080 ;
    END
  END master1_wb_adr_o[10]
  PIN master1_wb_adr_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END master1_wb_adr_o[11]
  PIN master1_wb_adr_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END master1_wb_adr_o[12]
  PIN master1_wb_adr_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END master1_wb_adr_o[13]
  PIN master1_wb_adr_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END master1_wb_adr_o[14]
  PIN master1_wb_adr_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END master1_wb_adr_o[15]
  PIN master1_wb_adr_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 645.360 4.000 645.960 ;
    END
  END master1_wb_adr_o[16]
  PIN master1_wb_adr_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END master1_wb_adr_o[17]
  PIN master1_wb_adr_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END master1_wb_adr_o[18]
  PIN master1_wb_adr_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END master1_wb_adr_o[19]
  PIN master1_wb_adr_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END master1_wb_adr_o[1]
  PIN master1_wb_adr_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.280 4.000 675.880 ;
    END
  END master1_wb_adr_o[20]
  PIN master1_wb_adr_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END master1_wb_adr_o[21]
  PIN master1_wb_adr_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END master1_wb_adr_o[22]
  PIN master1_wb_adr_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 698.400 4.000 699.000 ;
    END
  END master1_wb_adr_o[23]
  PIN master1_wb_adr_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END master1_wb_adr_o[24]
  PIN master1_wb_adr_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 713.360 4.000 713.960 ;
    END
  END master1_wb_adr_o[25]
  PIN master1_wb_adr_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END master1_wb_adr_o[26]
  PIN master1_wb_adr_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 728.320 4.000 728.920 ;
    END
  END master1_wb_adr_o[27]
  PIN master1_wb_adr_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END master1_wb_adr_o[2]
  PIN master1_wb_adr_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END master1_wb_adr_o[3]
  PIN master1_wb_adr_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END master1_wb_adr_o[4]
  PIN master1_wb_adr_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END master1_wb_adr_o[5]
  PIN master1_wb_adr_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END master1_wb_adr_o[6]
  PIN master1_wb_adr_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END master1_wb_adr_o[7]
  PIN master1_wb_adr_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END master1_wb_adr_o[8]
  PIN master1_wb_adr_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END master1_wb_adr_o[9]
  PIN master1_wb_cyc_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END master1_wb_cyc_o
  PIN master1_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END master1_wb_data_i[0]
  PIN master1_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END master1_wb_data_i[10]
  PIN master1_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END master1_wb_data_i[11]
  PIN master1_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.160 4.000 618.760 ;
    END
  END master1_wb_data_i[12]
  PIN master1_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END master1_wb_data_i[13]
  PIN master1_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.120 4.000 633.720 ;
    END
  END master1_wb_data_i[14]
  PIN master1_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END master1_wb_data_i[15]
  PIN master1_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.080 4.000 648.680 ;
    END
  END master1_wb_data_i[16]
  PIN master1_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END master1_wb_data_i[17]
  PIN master1_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END master1_wb_data_i[18]
  PIN master1_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END master1_wb_data_i[19]
  PIN master1_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END master1_wb_data_i[1]
  PIN master1_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END master1_wb_data_i[20]
  PIN master1_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END master1_wb_data_i[21]
  PIN master1_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.960 4.000 693.560 ;
    END
  END master1_wb_data_i[22]
  PIN master1_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END master1_wb_data_i[23]
  PIN master1_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.920 4.000 708.520 ;
    END
  END master1_wb_data_i[24]
  PIN master1_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END master1_wb_data_i[25]
  PIN master1_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END master1_wb_data_i[26]
  PIN master1_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END master1_wb_data_i[27]
  PIN master1_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END master1_wb_data_i[28]
  PIN master1_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 740.560 4.000 741.160 ;
    END
  END master1_wb_data_i[29]
  PIN master1_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 4.000 538.520 ;
    END
  END master1_wb_data_i[2]
  PIN master1_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 4.000 745.920 ;
    END
  END master1_wb_data_i[30]
  PIN master1_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.760 4.000 751.360 ;
    END
  END master1_wb_data_i[31]
  PIN master1_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END master1_wb_data_i[3]
  PIN master1_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 558.320 4.000 558.920 ;
    END
  END master1_wb_data_i[4]
  PIN master1_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END master1_wb_data_i[5]
  PIN master1_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END master1_wb_data_i[6]
  PIN master1_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END master1_wb_data_i[7]
  PIN master1_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END master1_wb_data_i[8]
  PIN master1_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END master1_wb_data_i[9]
  PIN master1_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END master1_wb_data_o[0]
  PIN master1_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END master1_wb_data_o[10]
  PIN master1_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 4.000 613.320 ;
    END
  END master1_wb_data_o[11]
  PIN master1_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.880 4.000 621.480 ;
    END
  END master1_wb_data_o[12]
  PIN master1_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END master1_wb_data_o[13]
  PIN master1_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END master1_wb_data_o[14]
  PIN master1_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END master1_wb_data_o[15]
  PIN master1_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END master1_wb_data_o[16]
  PIN master1_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END master1_wb_data_o[17]
  PIN master1_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.760 4.000 666.360 ;
    END
  END master1_wb_data_o[18]
  PIN master1_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END master1_wb_data_o[19]
  PIN master1_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END master1_wb_data_o[1]
  PIN master1_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END master1_wb_data_o[20]
  PIN master1_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END master1_wb_data_o[21]
  PIN master1_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.680 4.000 696.280 ;
    END
  END master1_wb_data_o[22]
  PIN master1_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END master1_wb_data_o[23]
  PIN master1_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END master1_wb_data_o[24]
  PIN master1_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END master1_wb_data_o[25]
  PIN master1_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END master1_wb_data_o[26]
  PIN master1_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END master1_wb_data_o[27]
  PIN master1_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END master1_wb_data_o[28]
  PIN master1_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END master1_wb_data_o[29]
  PIN master1_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END master1_wb_data_o[2]
  PIN master1_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END master1_wb_data_o[30]
  PIN master1_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.800 4.000 753.400 ;
    END
  END master1_wb_data_o[31]
  PIN master1_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END master1_wb_data_o[3]
  PIN master1_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 560.360 4.000 560.960 ;
    END
  END master1_wb_data_o[4]
  PIN master1_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END master1_wb_data_o[5]
  PIN master1_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END master1_wb_data_o[6]
  PIN master1_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.800 4.000 583.400 ;
    END
  END master1_wb_data_o[7]
  PIN master1_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END master1_wb_data_o[8]
  PIN master1_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.760 4.000 598.360 ;
    END
  END master1_wb_data_o[9]
  PIN master1_wb_error_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.280 4.000 505.880 ;
    END
  END master1_wb_error_i
  PIN master1_wb_sel_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.960 4.000 523.560 ;
    END
  END master1_wb_sel_o[0]
  PIN master1_wb_sel_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END master1_wb_sel_o[1]
  PIN master1_wb_sel_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END master1_wb_sel_o[2]
  PIN master1_wb_sel_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END master1_wb_sel_o[3]
  PIN master1_wb_stall_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END master1_wb_stall_i
  PIN master1_wb_stb_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.720 4.000 511.320 ;
    END
  END master1_wb_stb_o
  PIN master1_wb_we_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END master1_wb_we_o
  PIN master2_wb_ack_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END master2_wb_ack_i
  PIN master2_wb_adr_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END master2_wb_adr_o[0]
  PIN master2_wb_adr_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END master2_wb_adr_o[10]
  PIN master2_wb_adr_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END master2_wb_adr_o[11]
  PIN master2_wb_adr_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END master2_wb_adr_o[12]
  PIN master2_wb_adr_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END master2_wb_adr_o[13]
  PIN master2_wb_adr_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END master2_wb_adr_o[14]
  PIN master2_wb_adr_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END master2_wb_adr_o[15]
  PIN master2_wb_adr_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END master2_wb_adr_o[16]
  PIN master2_wb_adr_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END master2_wb_adr_o[17]
  PIN master2_wb_adr_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END master2_wb_adr_o[18]
  PIN master2_wb_adr_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END master2_wb_adr_o[19]
  PIN master2_wb_adr_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END master2_wb_adr_o[1]
  PIN master2_wb_adr_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END master2_wb_adr_o[20]
  PIN master2_wb_adr_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END master2_wb_adr_o[21]
  PIN master2_wb_adr_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END master2_wb_adr_o[22]
  PIN master2_wb_adr_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.720 4.000 443.320 ;
    END
  END master2_wb_adr_o[23]
  PIN master2_wb_adr_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END master2_wb_adr_o[24]
  PIN master2_wb_adr_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END master2_wb_adr_o[25]
  PIN master2_wb_adr_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END master2_wb_adr_o[26]
  PIN master2_wb_adr_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END master2_wb_adr_o[27]
  PIN master2_wb_adr_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END master2_wb_adr_o[2]
  PIN master2_wb_adr_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END master2_wb_adr_o[3]
  PIN master2_wb_adr_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END master2_wb_adr_o[4]
  PIN master2_wb_adr_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END master2_wb_adr_o[5]
  PIN master2_wb_adr_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END master2_wb_adr_o[6]
  PIN master2_wb_adr_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END master2_wb_adr_o[7]
  PIN master2_wb_adr_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END master2_wb_adr_o[8]
  PIN master2_wb_adr_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END master2_wb_adr_o[9]
  PIN master2_wb_cyc_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END master2_wb_cyc_o
  PIN master2_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END master2_wb_data_i[0]
  PIN master2_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END master2_wb_data_i[10]
  PIN master2_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END master2_wb_data_i[11]
  PIN master2_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END master2_wb_data_i[12]
  PIN master2_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END master2_wb_data_i[13]
  PIN master2_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END master2_wb_data_i[14]
  PIN master2_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END master2_wb_data_i[15]
  PIN master2_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END master2_wb_data_i[16]
  PIN master2_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.560 4.000 401.160 ;
    END
  END master2_wb_data_i[17]
  PIN master2_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END master2_wb_data_i[18]
  PIN master2_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END master2_wb_data_i[19]
  PIN master2_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END master2_wb_data_i[1]
  PIN master2_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END master2_wb_data_i[20]
  PIN master2_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END master2_wb_data_i[21]
  PIN master2_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END master2_wb_data_i[22]
  PIN master2_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END master2_wb_data_i[23]
  PIN master2_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END master2_wb_data_i[24]
  PIN master2_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 460.400 4.000 461.000 ;
    END
  END master2_wb_data_i[25]
  PIN master2_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END master2_wb_data_i[26]
  PIN master2_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 475.360 4.000 475.960 ;
    END
  END master2_wb_data_i[27]
  PIN master2_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END master2_wb_data_i[28]
  PIN master2_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END master2_wb_data_i[29]
  PIN master2_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END master2_wb_data_i[2]
  PIN master2_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 490.320 4.000 490.920 ;
    END
  END master2_wb_data_i[30]
  PIN master2_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.760 4.000 496.360 ;
    END
  END master2_wb_data_i[31]
  PIN master2_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END master2_wb_data_i[3]
  PIN master2_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END master2_wb_data_i[4]
  PIN master2_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END master2_wb_data_i[5]
  PIN master2_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END master2_wb_data_i[6]
  PIN master2_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END master2_wb_data_i[7]
  PIN master2_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END master2_wb_data_i[8]
  PIN master2_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END master2_wb_data_i[9]
  PIN master2_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END master2_wb_data_o[0]
  PIN master2_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END master2_wb_data_o[10]
  PIN master2_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END master2_wb_data_o[11]
  PIN master2_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END master2_wb_data_o[12]
  PIN master2_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END master2_wb_data_o[13]
  PIN master2_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END master2_wb_data_o[14]
  PIN master2_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.320 4.000 388.920 ;
    END
  END master2_wb_data_o[15]
  PIN master2_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END master2_wb_data_o[16]
  PIN master2_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END master2_wb_data_o[17]
  PIN master2_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END master2_wb_data_o[18]
  PIN master2_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END master2_wb_data_o[19]
  PIN master2_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END master2_wb_data_o[1]
  PIN master2_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END master2_wb_data_o[20]
  PIN master2_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END master2_wb_data_o[21]
  PIN master2_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END master2_wb_data_o[22]
  PIN master2_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.160 4.000 448.760 ;
    END
  END master2_wb_data_o[23]
  PIN master2_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END master2_wb_data_o[24]
  PIN master2_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END master2_wb_data_o[25]
  PIN master2_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END master2_wb_data_o[26]
  PIN master2_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END master2_wb_data_o[27]
  PIN master2_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END master2_wb_data_o[28]
  PIN master2_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END master2_wb_data_o[29]
  PIN master2_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END master2_wb_data_o[2]
  PIN master2_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END master2_wb_data_o[30]
  PIN master2_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END master2_wb_data_o[31]
  PIN master2_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END master2_wb_data_o[3]
  PIN master2_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END master2_wb_data_o[4]
  PIN master2_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END master2_wb_data_o[5]
  PIN master2_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END master2_wb_data_o[6]
  PIN master2_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END master2_wb_data_o[7]
  PIN master2_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END master2_wb_data_o[8]
  PIN master2_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END master2_wb_data_o[9]
  PIN master2_wb_error_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END master2_wb_error_i
  PIN master2_wb_sel_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END master2_wb_sel_o[0]
  PIN master2_wb_sel_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END master2_wb_sel_o[1]
  PIN master2_wb_sel_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END master2_wb_sel_o[2]
  PIN master2_wb_sel_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END master2_wb_sel_o[3]
  PIN master2_wb_stall_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END master2_wb_stall_i
  PIN master2_wb_stb_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END master2_wb_stb_o
  PIN master2_wb_we_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END master2_wb_we_o
  PIN probe_master0_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END probe_master0_currentSlave[0]
  PIN probe_master0_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END probe_master0_currentSlave[1]
  PIN probe_master1_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END probe_master1_currentSlave[0]
  PIN probe_master1_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END probe_master1_currentSlave[1]
  PIN probe_master2_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END probe_master2_currentSlave[0]
  PIN probe_master2_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END probe_master2_currentSlave[1]
  PIN probe_master3_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END probe_master3_currentSlave[0]
  PIN probe_master3_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END probe_master3_currentSlave[1]
  PIN probe_slave0_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END probe_slave0_currentMaster[0]
  PIN probe_slave0_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END probe_slave0_currentMaster[1]
  PIN probe_slave1_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END probe_slave1_currentMaster[0]
  PIN probe_slave1_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END probe_slave1_currentMaster[1]
  PIN probe_slave2_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END probe_slave2_currentMaster[0]
  PIN probe_slave2_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END probe_slave2_currentMaster[1]
  PIN probe_slave3_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END probe_slave3_currentMaster[0]
  PIN probe_slave3_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END probe_slave3_currentMaster[1]
  PIN slave0_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.520 4.000 756.120 ;
    END
  END slave0_wb_ack_o
  PIN slave0_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 770.480 4.000 771.080 ;
    END
  END slave0_wb_adr_i[0]
  PIN slave0_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 855.480 4.000 856.080 ;
    END
  END slave0_wb_adr_i[10]
  PIN slave0_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.960 4.000 863.560 ;
    END
  END slave0_wb_adr_i[11]
  PIN slave0_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END slave0_wb_adr_i[12]
  PIN slave0_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.920 4.000 878.520 ;
    END
  END slave0_wb_adr_i[13]
  PIN slave0_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 885.400 4.000 886.000 ;
    END
  END slave0_wb_adr_i[14]
  PIN slave0_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.880 4.000 893.480 ;
    END
  END slave0_wb_adr_i[15]
  PIN slave0_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 900.360 4.000 900.960 ;
    END
  END slave0_wb_adr_i[16]
  PIN slave0_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END slave0_wb_adr_i[17]
  PIN slave0_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 915.320 4.000 915.920 ;
    END
  END slave0_wb_adr_i[18]
  PIN slave0_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.800 4.000 923.400 ;
    END
  END slave0_wb_adr_i[19]
  PIN slave0_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END slave0_wb_adr_i[1]
  PIN slave0_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END slave0_wb_adr_i[20]
  PIN slave0_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END slave0_wb_adr_i[21]
  PIN slave0_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.920 4.000 946.520 ;
    END
  END slave0_wb_adr_i[22]
  PIN slave0_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 953.400 4.000 954.000 ;
    END
  END slave0_wb_adr_i[23]
  PIN slave0_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.880 4.000 791.480 ;
    END
  END slave0_wb_adr_i[2]
  PIN slave0_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 800.400 4.000 801.000 ;
    END
  END slave0_wb_adr_i[3]
  PIN slave0_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 4.000 811.200 ;
    END
  END slave0_wb_adr_i[4]
  PIN slave0_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.080 4.000 818.680 ;
    END
  END slave0_wb_adr_i[5]
  PIN slave0_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END slave0_wb_adr_i[6]
  PIN slave0_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END slave0_wb_adr_i[7]
  PIN slave0_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END slave0_wb_adr_i[8]
  PIN slave0_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.000 4.000 848.600 ;
    END
  END slave0_wb_adr_i[9]
  PIN slave0_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END slave0_wb_cyc_i
  PIN slave0_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END slave0_wb_data_i[0]
  PIN slave0_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.200 4.000 858.800 ;
    END
  END slave0_wb_data_i[10]
  PIN slave0_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.680 4.000 866.280 ;
    END
  END slave0_wb_data_i[11]
  PIN slave0_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.160 4.000 873.760 ;
    END
  END slave0_wb_data_i[12]
  PIN slave0_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END slave0_wb_data_i[13]
  PIN slave0_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END slave0_wb_data_i[14]
  PIN slave0_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 895.600 4.000 896.200 ;
    END
  END slave0_wb_data_i[15]
  PIN slave0_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.080 4.000 903.680 ;
    END
  END slave0_wb_data_i[16]
  PIN slave0_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 910.560 4.000 911.160 ;
    END
  END slave0_wb_data_i[17]
  PIN slave0_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END slave0_wb_data_i[18]
  PIN slave0_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 925.520 4.000 926.120 ;
    END
  END slave0_wb_data_i[19]
  PIN slave0_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 783.400 4.000 784.000 ;
    END
  END slave0_wb_data_i[1]
  PIN slave0_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.000 4.000 933.600 ;
    END
  END slave0_wb_data_i[20]
  PIN slave0_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 940.480 4.000 941.080 ;
    END
  END slave0_wb_data_i[21]
  PIN slave0_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.960 4.000 948.560 ;
    END
  END slave0_wb_data_i[22]
  PIN slave0_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END slave0_wb_data_i[23]
  PIN slave0_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.880 4.000 961.480 ;
    END
  END slave0_wb_data_i[24]
  PIN slave0_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END slave0_wb_data_i[25]
  PIN slave0_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 970.400 4.000 971.000 ;
    END
  END slave0_wb_data_i[26]
  PIN slave0_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END slave0_wb_data_i[27]
  PIN slave0_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END slave0_wb_data_i[28]
  PIN slave0_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 985.360 4.000 985.960 ;
    END
  END slave0_wb_data_i[29]
  PIN slave0_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END slave0_wb_data_i[2]
  PIN slave0_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.800 4.000 991.400 ;
    END
  END slave0_wb_data_i[30]
  PIN slave0_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 995.560 4.000 996.160 ;
    END
  END slave0_wb_data_i[31]
  PIN slave0_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.120 4.000 803.720 ;
    END
  END slave0_wb_data_i[3]
  PIN slave0_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END slave0_wb_data_i[4]
  PIN slave0_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.800 4.000 821.400 ;
    END
  END slave0_wb_data_i[5]
  PIN slave0_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END slave0_wb_data_i[6]
  PIN slave0_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.760 4.000 836.360 ;
    END
  END slave0_wb_data_i[7]
  PIN slave0_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END slave0_wb_data_i[8]
  PIN slave0_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.720 4.000 851.320 ;
    END
  END slave0_wb_data_i[9]
  PIN slave0_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.920 4.000 776.520 ;
    END
  END slave0_wb_data_o[0]
  PIN slave0_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.920 4.000 861.520 ;
    END
  END slave0_wb_data_o[10]
  PIN slave0_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 868.400 4.000 869.000 ;
    END
  END slave0_wb_data_o[11]
  PIN slave0_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END slave0_wb_data_o[12]
  PIN slave0_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 883.360 4.000 883.960 ;
    END
  END slave0_wb_data_o[13]
  PIN slave0_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END slave0_wb_data_o[14]
  PIN slave0_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 898.320 4.000 898.920 ;
    END
  END slave0_wb_data_o[15]
  PIN slave0_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END slave0_wb_data_o[16]
  PIN slave0_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 913.280 4.000 913.880 ;
    END
  END slave0_wb_data_o[17]
  PIN slave0_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.760 4.000 921.360 ;
    END
  END slave0_wb_data_o[18]
  PIN slave0_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END slave0_wb_data_o[19]
  PIN slave0_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END slave0_wb_data_o[1]
  PIN slave0_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.720 4.000 936.320 ;
    END
  END slave0_wb_data_o[20]
  PIN slave0_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.200 4.000 943.800 ;
    END
  END slave0_wb_data_o[21]
  PIN slave0_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.680 4.000 951.280 ;
    END
  END slave0_wb_data_o[22]
  PIN slave0_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.160 4.000 958.760 ;
    END
  END slave0_wb_data_o[23]
  PIN slave0_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.920 4.000 963.520 ;
    END
  END slave0_wb_data_o[24]
  PIN slave0_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 968.360 4.000 968.960 ;
    END
  END slave0_wb_data_o[25]
  PIN slave0_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.120 4.000 973.720 ;
    END
  END slave0_wb_data_o[26]
  PIN slave0_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.880 4.000 978.480 ;
    END
  END slave0_wb_data_o[27]
  PIN slave0_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END slave0_wb_data_o[28]
  PIN slave0_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 988.080 4.000 988.680 ;
    END
  END slave0_wb_data_o[29]
  PIN slave0_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END slave0_wb_data_o[2]
  PIN slave0_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END slave0_wb_data_o[30]
  PIN slave0_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 998.280 4.000 998.880 ;
    END
  END slave0_wb_data_o[31]
  PIN slave0_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END slave0_wb_data_o[3]
  PIN slave0_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END slave0_wb_data_o[4]
  PIN slave0_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END slave0_wb_data_o[5]
  PIN slave0_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 830.320 4.000 830.920 ;
    END
  END slave0_wb_data_o[6]
  PIN slave0_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END slave0_wb_data_o[7]
  PIN slave0_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.280 4.000 845.880 ;
    END
  END slave0_wb_data_o[8]
  PIN slave0_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END slave0_wb_data_o[9]
  PIN slave0_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END slave0_wb_error_o
  PIN slave0_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.960 4.000 778.560 ;
    END
  END slave0_wb_sel_i[0]
  PIN slave0_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.160 4.000 788.760 ;
    END
  END slave0_wb_sel_i[1]
  PIN slave0_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 798.360 4.000 798.960 ;
    END
  END slave0_wb_sel_i[2]
  PIN slave0_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END slave0_wb_sel_i[3]
  PIN slave0_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END slave0_wb_stall_o
  PIN slave0_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END slave0_wb_stb_i
  PIN slave0_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 767.760 4.000 768.360 ;
    END
  END slave0_wb_we_i
  PIN slave1_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END slave1_wb_ack_o
  PIN slave1_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END slave1_wb_adr_i[0]
  PIN slave1_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END slave1_wb_adr_i[10]
  PIN slave1_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END slave1_wb_adr_i[11]
  PIN slave1_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END slave1_wb_adr_i[12]
  PIN slave1_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END slave1_wb_adr_i[13]
  PIN slave1_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END slave1_wb_adr_i[14]
  PIN slave1_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END slave1_wb_adr_i[15]
  PIN slave1_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END slave1_wb_adr_i[16]
  PIN slave1_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END slave1_wb_adr_i[17]
  PIN slave1_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END slave1_wb_adr_i[18]
  PIN slave1_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END slave1_wb_adr_i[19]
  PIN slave1_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END slave1_wb_adr_i[1]
  PIN slave1_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END slave1_wb_adr_i[20]
  PIN slave1_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END slave1_wb_adr_i[21]
  PIN slave1_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END slave1_wb_adr_i[22]
  PIN slave1_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END slave1_wb_adr_i[23]
  PIN slave1_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END slave1_wb_adr_i[2]
  PIN slave1_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END slave1_wb_adr_i[3]
  PIN slave1_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END slave1_wb_adr_i[4]
  PIN slave1_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END slave1_wb_adr_i[5]
  PIN slave1_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END slave1_wb_adr_i[6]
  PIN slave1_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END slave1_wb_adr_i[7]
  PIN slave1_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END slave1_wb_adr_i[8]
  PIN slave1_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END slave1_wb_adr_i[9]
  PIN slave1_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END slave1_wb_cyc_i
  PIN slave1_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END slave1_wb_data_i[0]
  PIN slave1_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END slave1_wb_data_i[10]
  PIN slave1_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END slave1_wb_data_i[11]
  PIN slave1_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END slave1_wb_data_i[12]
  PIN slave1_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END slave1_wb_data_i[13]
  PIN slave1_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END slave1_wb_data_i[14]
  PIN slave1_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END slave1_wb_data_i[15]
  PIN slave1_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END slave1_wb_data_i[16]
  PIN slave1_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END slave1_wb_data_i[17]
  PIN slave1_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END slave1_wb_data_i[18]
  PIN slave1_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END slave1_wb_data_i[19]
  PIN slave1_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END slave1_wb_data_i[1]
  PIN slave1_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END slave1_wb_data_i[20]
  PIN slave1_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END slave1_wb_data_i[21]
  PIN slave1_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END slave1_wb_data_i[22]
  PIN slave1_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END slave1_wb_data_i[23]
  PIN slave1_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END slave1_wb_data_i[24]
  PIN slave1_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END slave1_wb_data_i[25]
  PIN slave1_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END slave1_wb_data_i[26]
  PIN slave1_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END slave1_wb_data_i[27]
  PIN slave1_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END slave1_wb_data_i[28]
  PIN slave1_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END slave1_wb_data_i[29]
  PIN slave1_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END slave1_wb_data_i[2]
  PIN slave1_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END slave1_wb_data_i[30]
  PIN slave1_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END slave1_wb_data_i[31]
  PIN slave1_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END slave1_wb_data_i[3]
  PIN slave1_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END slave1_wb_data_i[4]
  PIN slave1_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END slave1_wb_data_i[5]
  PIN slave1_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END slave1_wb_data_i[6]
  PIN slave1_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END slave1_wb_data_i[7]
  PIN slave1_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END slave1_wb_data_i[8]
  PIN slave1_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END slave1_wb_data_i[9]
  PIN slave1_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END slave1_wb_data_o[0]
  PIN slave1_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END slave1_wb_data_o[10]
  PIN slave1_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END slave1_wb_data_o[11]
  PIN slave1_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END slave1_wb_data_o[12]
  PIN slave1_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END slave1_wb_data_o[13]
  PIN slave1_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END slave1_wb_data_o[14]
  PIN slave1_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END slave1_wb_data_o[15]
  PIN slave1_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END slave1_wb_data_o[16]
  PIN slave1_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END slave1_wb_data_o[17]
  PIN slave1_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END slave1_wb_data_o[18]
  PIN slave1_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END slave1_wb_data_o[19]
  PIN slave1_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END slave1_wb_data_o[1]
  PIN slave1_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END slave1_wb_data_o[20]
  PIN slave1_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END slave1_wb_data_o[21]
  PIN slave1_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END slave1_wb_data_o[22]
  PIN slave1_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END slave1_wb_data_o[23]
  PIN slave1_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END slave1_wb_data_o[24]
  PIN slave1_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END slave1_wb_data_o[25]
  PIN slave1_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END slave1_wb_data_o[26]
  PIN slave1_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END slave1_wb_data_o[27]
  PIN slave1_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END slave1_wb_data_o[28]
  PIN slave1_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END slave1_wb_data_o[29]
  PIN slave1_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END slave1_wb_data_o[2]
  PIN slave1_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END slave1_wb_data_o[30]
  PIN slave1_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END slave1_wb_data_o[31]
  PIN slave1_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END slave1_wb_data_o[3]
  PIN slave1_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END slave1_wb_data_o[4]
  PIN slave1_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END slave1_wb_data_o[5]
  PIN slave1_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END slave1_wb_data_o[6]
  PIN slave1_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END slave1_wb_data_o[7]
  PIN slave1_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END slave1_wb_data_o[8]
  PIN slave1_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END slave1_wb_data_o[9]
  PIN slave1_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END slave1_wb_error_o
  PIN slave1_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END slave1_wb_sel_i[0]
  PIN slave1_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END slave1_wb_sel_i[1]
  PIN slave1_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END slave1_wb_sel_i[2]
  PIN slave1_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END slave1_wb_sel_i[3]
  PIN slave1_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END slave1_wb_stall_o
  PIN slave1_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END slave1_wb_stb_i
  PIN slave1_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END slave1_wb_we_i
  PIN slave2_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 996.000 1.750 1000.000 ;
    END
  END slave2_wb_ack_o
  PIN slave2_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 996.000 22.910 1000.000 ;
    END
  END slave2_wb_adr_i[0]
  PIN slave2_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 996.000 144.350 1000.000 ;
    END
  END slave2_wb_adr_i[10]
  PIN slave2_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 996.000 154.930 1000.000 ;
    END
  END slave2_wb_adr_i[11]
  PIN slave2_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 996.000 165.970 1000.000 ;
    END
  END slave2_wb_adr_i[12]
  PIN slave2_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 996.000 176.550 1000.000 ;
    END
  END slave2_wb_adr_i[13]
  PIN slave2_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 996.000 187.130 1000.000 ;
    END
  END slave2_wb_adr_i[14]
  PIN slave2_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 996.000 198.170 1000.000 ;
    END
  END slave2_wb_adr_i[15]
  PIN slave2_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 996.000 208.750 1000.000 ;
    END
  END slave2_wb_adr_i[16]
  PIN slave2_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 996.000 219.330 1000.000 ;
    END
  END slave2_wb_adr_i[17]
  PIN slave2_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 996.000 229.910 1000.000 ;
    END
  END slave2_wb_adr_i[18]
  PIN slave2_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 996.000 240.950 1000.000 ;
    END
  END slave2_wb_adr_i[19]
  PIN slave2_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 996.000 37.170 1000.000 ;
    END
  END slave2_wb_adr_i[1]
  PIN slave2_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 996.000 251.530 1000.000 ;
    END
  END slave2_wb_adr_i[20]
  PIN slave2_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 996.000 262.110 1000.000 ;
    END
  END slave2_wb_adr_i[21]
  PIN slave2_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 996.000 273.150 1000.000 ;
    END
  END slave2_wb_adr_i[22]
  PIN slave2_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 996.000 283.730 1000.000 ;
    END
  END slave2_wb_adr_i[23]
  PIN slave2_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 996.000 51.430 1000.000 ;
    END
  END slave2_wb_adr_i[2]
  PIN slave2_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 996.000 65.690 1000.000 ;
    END
  END slave2_wb_adr_i[3]
  PIN slave2_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 996.000 79.950 1000.000 ;
    END
  END slave2_wb_adr_i[4]
  PIN slave2_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 996.000 90.990 1000.000 ;
    END
  END slave2_wb_adr_i[5]
  PIN slave2_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 996.000 101.570 1000.000 ;
    END
  END slave2_wb_adr_i[6]
  PIN slave2_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 996.000 112.150 1000.000 ;
    END
  END slave2_wb_adr_i[7]
  PIN slave2_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 996.000 123.190 1000.000 ;
    END
  END slave2_wb_adr_i[8]
  PIN slave2_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 996.000 133.770 1000.000 ;
    END
  END slave2_wb_adr_i[9]
  PIN slave2_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 996.000 4.970 1000.000 ;
    END
  END slave2_wb_cyc_i
  PIN slave2_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 996.000 26.590 1000.000 ;
    END
  END slave2_wb_data_i[0]
  PIN slave2_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 996.000 148.030 1000.000 ;
    END
  END slave2_wb_data_i[10]
  PIN slave2_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 996.000 158.610 1000.000 ;
    END
  END slave2_wb_data_i[11]
  PIN slave2_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 996.000 169.190 1000.000 ;
    END
  END slave2_wb_data_i[12]
  PIN slave2_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 996.000 180.230 1000.000 ;
    END
  END slave2_wb_data_i[13]
  PIN slave2_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 996.000 190.810 1000.000 ;
    END
  END slave2_wb_data_i[14]
  PIN slave2_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 996.000 201.390 1000.000 ;
    END
  END slave2_wb_data_i[15]
  PIN slave2_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 996.000 212.430 1000.000 ;
    END
  END slave2_wb_data_i[16]
  PIN slave2_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 996.000 223.010 1000.000 ;
    END
  END slave2_wb_data_i[17]
  PIN slave2_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 996.000 233.590 1000.000 ;
    END
  END slave2_wb_data_i[18]
  PIN slave2_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 996.000 244.630 1000.000 ;
    END
  END slave2_wb_data_i[19]
  PIN slave2_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 996.000 40.850 1000.000 ;
    END
  END slave2_wb_data_i[1]
  PIN slave2_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 996.000 255.210 1000.000 ;
    END
  END slave2_wb_data_i[20]
  PIN slave2_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 996.000 265.790 1000.000 ;
    END
  END slave2_wb_data_i[21]
  PIN slave2_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 996.000 276.370 1000.000 ;
    END
  END slave2_wb_data_i[22]
  PIN slave2_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 996.000 287.410 1000.000 ;
    END
  END slave2_wb_data_i[23]
  PIN slave2_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 996.000 294.310 1000.000 ;
    END
  END slave2_wb_data_i[24]
  PIN slave2_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 996.000 301.670 1000.000 ;
    END
  END slave2_wb_data_i[25]
  PIN slave2_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 996.000 308.570 1000.000 ;
    END
  END slave2_wb_data_i[26]
  PIN slave2_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 996.000 315.930 1000.000 ;
    END
  END slave2_wb_data_i[27]
  PIN slave2_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 996.000 322.830 1000.000 ;
    END
  END slave2_wb_data_i[28]
  PIN slave2_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 996.000 330.190 1000.000 ;
    END
  END slave2_wb_data_i[29]
  PIN slave2_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 996.000 55.110 1000.000 ;
    END
  END slave2_wb_data_i[2]
  PIN slave2_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 996.000 337.090 1000.000 ;
    END
  END slave2_wb_data_i[30]
  PIN slave2_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 996.000 344.450 1000.000 ;
    END
  END slave2_wb_data_i[31]
  PIN slave2_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 996.000 69.370 1000.000 ;
    END
  END slave2_wb_data_i[3]
  PIN slave2_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 996.000 83.630 1000.000 ;
    END
  END slave2_wb_data_i[4]
  PIN slave2_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 996.000 94.210 1000.000 ;
    END
  END slave2_wb_data_i[5]
  PIN slave2_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 996.000 105.250 1000.000 ;
    END
  END slave2_wb_data_i[6]
  PIN slave2_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 996.000 115.830 1000.000 ;
    END
  END slave2_wb_data_i[7]
  PIN slave2_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 996.000 126.410 1000.000 ;
    END
  END slave2_wb_data_i[8]
  PIN slave2_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 996.000 137.450 1000.000 ;
    END
  END slave2_wb_data_i[9]
  PIN slave2_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 996.000 30.270 1000.000 ;
    END
  END slave2_wb_data_o[0]
  PIN slave2_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 996.000 151.710 1000.000 ;
    END
  END slave2_wb_data_o[10]
  PIN slave2_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 996.000 162.290 1000.000 ;
    END
  END slave2_wb_data_o[11]
  PIN slave2_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 996.000 172.870 1000.000 ;
    END
  END slave2_wb_data_o[12]
  PIN slave2_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 996.000 183.910 1000.000 ;
    END
  END slave2_wb_data_o[13]
  PIN slave2_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 996.000 194.490 1000.000 ;
    END
  END slave2_wb_data_o[14]
  PIN slave2_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 996.000 205.070 1000.000 ;
    END
  END slave2_wb_data_o[15]
  PIN slave2_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 996.000 215.650 1000.000 ;
    END
  END slave2_wb_data_o[16]
  PIN slave2_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 996.000 226.690 1000.000 ;
    END
  END slave2_wb_data_o[17]
  PIN slave2_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 996.000 237.270 1000.000 ;
    END
  END slave2_wb_data_o[18]
  PIN slave2_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 996.000 247.850 1000.000 ;
    END
  END slave2_wb_data_o[19]
  PIN slave2_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 996.000 44.530 1000.000 ;
    END
  END slave2_wb_data_o[1]
  PIN slave2_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 996.000 258.890 1000.000 ;
    END
  END slave2_wb_data_o[20]
  PIN slave2_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 996.000 269.470 1000.000 ;
    END
  END slave2_wb_data_o[21]
  PIN slave2_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 996.000 280.050 1000.000 ;
    END
  END slave2_wb_data_o[22]
  PIN slave2_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 996.000 290.630 1000.000 ;
    END
  END slave2_wb_data_o[23]
  PIN slave2_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 996.000 297.990 1000.000 ;
    END
  END slave2_wb_data_o[24]
  PIN slave2_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 996.000 305.350 1000.000 ;
    END
  END slave2_wb_data_o[25]
  PIN slave2_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 996.000 312.250 1000.000 ;
    END
  END slave2_wb_data_o[26]
  PIN slave2_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 996.000 319.610 1000.000 ;
    END
  END slave2_wb_data_o[27]
  PIN slave2_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 996.000 326.510 1000.000 ;
    END
  END slave2_wb_data_o[28]
  PIN slave2_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 996.000 333.870 1000.000 ;
    END
  END slave2_wb_data_o[29]
  PIN slave2_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 996.000 58.790 1000.000 ;
    END
  END slave2_wb_data_o[2]
  PIN slave2_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 996.000 340.770 1000.000 ;
    END
  END slave2_wb_data_o[30]
  PIN slave2_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 996.000 348.130 1000.000 ;
    END
  END slave2_wb_data_o[31]
  PIN slave2_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 996.000 73.050 1000.000 ;
    END
  END slave2_wb_data_o[3]
  PIN slave2_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 996.000 87.310 1000.000 ;
    END
  END slave2_wb_data_o[4]
  PIN slave2_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 996.000 97.890 1000.000 ;
    END
  END slave2_wb_data_o[5]
  PIN slave2_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 996.000 108.470 1000.000 ;
    END
  END slave2_wb_data_o[6]
  PIN slave2_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 996.000 119.510 1000.000 ;
    END
  END slave2_wb_data_o[7]
  PIN slave2_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 996.000 130.090 1000.000 ;
    END
  END slave2_wb_data_o[8]
  PIN slave2_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 996.000 140.670 1000.000 ;
    END
  END slave2_wb_data_o[9]
  PIN slave2_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 996.000 8.650 1000.000 ;
    END
  END slave2_wb_error_o
  PIN slave2_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 996.000 33.490 1000.000 ;
    END
  END slave2_wb_sel_i[0]
  PIN slave2_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 996.000 47.750 1000.000 ;
    END
  END slave2_wb_sel_i[1]
  PIN slave2_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 996.000 62.470 1000.000 ;
    END
  END slave2_wb_sel_i[2]
  PIN slave2_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 996.000 76.730 1000.000 ;
    END
  END slave2_wb_sel_i[3]
  PIN slave2_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 996.000 12.330 1000.000 ;
    END
  END slave2_wb_stall_o
  PIN slave2_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 996.000 16.010 1000.000 ;
    END
  END slave2_wb_stb_i
  PIN slave2_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 996.000 19.230 1000.000 ;
    END
  END slave2_wb_we_i
  PIN slave3_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 4.800 350.000 5.400 ;
    END
  END slave3_wb_ack_o
  PIN slave3_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 66.000 350.000 66.600 ;
    END
  END slave3_wb_adr_i[0]
  PIN slave3_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 412.800 350.000 413.400 ;
    END
  END slave3_wb_adr_i[10]
  PIN slave3_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 443.400 350.000 444.000 ;
    END
  END slave3_wb_adr_i[11]
  PIN slave3_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 474.000 350.000 474.600 ;
    END
  END slave3_wb_adr_i[12]
  PIN slave3_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 504.600 350.000 505.200 ;
    END
  END slave3_wb_adr_i[13]
  PIN slave3_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 535.200 350.000 535.800 ;
    END
  END slave3_wb_adr_i[14]
  PIN slave3_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 565.800 350.000 566.400 ;
    END
  END slave3_wb_adr_i[15]
  PIN slave3_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 596.400 350.000 597.000 ;
    END
  END slave3_wb_adr_i[16]
  PIN slave3_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 627.000 350.000 627.600 ;
    END
  END slave3_wb_adr_i[17]
  PIN slave3_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 657.600 350.000 658.200 ;
    END
  END slave3_wb_adr_i[18]
  PIN slave3_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 688.200 350.000 688.800 ;
    END
  END slave3_wb_adr_i[19]
  PIN slave3_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 106.800 350.000 107.400 ;
    END
  END slave3_wb_adr_i[1]
  PIN slave3_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 718.800 350.000 719.400 ;
    END
  END slave3_wb_adr_i[20]
  PIN slave3_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 749.400 350.000 750.000 ;
    END
  END slave3_wb_adr_i[21]
  PIN slave3_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 780.000 350.000 780.600 ;
    END
  END slave3_wb_adr_i[22]
  PIN slave3_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 810.600 350.000 811.200 ;
    END
  END slave3_wb_adr_i[23]
  PIN slave3_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 147.600 350.000 148.200 ;
    END
  END slave3_wb_adr_i[2]
  PIN slave3_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 188.400 350.000 189.000 ;
    END
  END slave3_wb_adr_i[3]
  PIN slave3_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 229.200 350.000 229.800 ;
    END
  END slave3_wb_adr_i[4]
  PIN slave3_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 259.800 350.000 260.400 ;
    END
  END slave3_wb_adr_i[5]
  PIN slave3_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 290.400 350.000 291.000 ;
    END
  END slave3_wb_adr_i[6]
  PIN slave3_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 321.000 350.000 321.600 ;
    END
  END slave3_wb_adr_i[7]
  PIN slave3_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 351.600 350.000 352.200 ;
    END
  END slave3_wb_adr_i[8]
  PIN slave3_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 382.200 350.000 382.800 ;
    END
  END slave3_wb_adr_i[9]
  PIN slave3_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 15.000 350.000 15.600 ;
    END
  END slave3_wb_cyc_i
  PIN slave3_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 76.200 350.000 76.800 ;
    END
  END slave3_wb_data_i[0]
  PIN slave3_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 423.000 350.000 423.600 ;
    END
  END slave3_wb_data_i[10]
  PIN slave3_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 453.600 350.000 454.200 ;
    END
  END slave3_wb_data_i[11]
  PIN slave3_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 484.200 350.000 484.800 ;
    END
  END slave3_wb_data_i[12]
  PIN slave3_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 514.800 350.000 515.400 ;
    END
  END slave3_wb_data_i[13]
  PIN slave3_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 545.400 350.000 546.000 ;
    END
  END slave3_wb_data_i[14]
  PIN slave3_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 576.000 350.000 576.600 ;
    END
  END slave3_wb_data_i[15]
  PIN slave3_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 606.600 350.000 607.200 ;
    END
  END slave3_wb_data_i[16]
  PIN slave3_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 637.200 350.000 637.800 ;
    END
  END slave3_wb_data_i[17]
  PIN slave3_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 667.800 350.000 668.400 ;
    END
  END slave3_wb_data_i[18]
  PIN slave3_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 698.400 350.000 699.000 ;
    END
  END slave3_wb_data_i[19]
  PIN slave3_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 117.000 350.000 117.600 ;
    END
  END slave3_wb_data_i[1]
  PIN slave3_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 729.000 350.000 729.600 ;
    END
  END slave3_wb_data_i[20]
  PIN slave3_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 759.600 350.000 760.200 ;
    END
  END slave3_wb_data_i[21]
  PIN slave3_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 790.200 350.000 790.800 ;
    END
  END slave3_wb_data_i[22]
  PIN slave3_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 820.800 350.000 821.400 ;
    END
  END slave3_wb_data_i[23]
  PIN slave3_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 841.200 350.000 841.800 ;
    END
  END slave3_wb_data_i[24]
  PIN slave3_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 861.600 350.000 862.200 ;
    END
  END slave3_wb_data_i[25]
  PIN slave3_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 882.000 350.000 882.600 ;
    END
  END slave3_wb_data_i[26]
  PIN slave3_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 902.400 350.000 903.000 ;
    END
  END slave3_wb_data_i[27]
  PIN slave3_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 922.800 350.000 923.400 ;
    END
  END slave3_wb_data_i[28]
  PIN slave3_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 943.200 350.000 943.800 ;
    END
  END slave3_wb_data_i[29]
  PIN slave3_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 157.800 350.000 158.400 ;
    END
  END slave3_wb_data_i[2]
  PIN slave3_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 963.600 350.000 964.200 ;
    END
  END slave3_wb_data_i[30]
  PIN slave3_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 984.000 350.000 984.600 ;
    END
  END slave3_wb_data_i[31]
  PIN slave3_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 198.600 350.000 199.200 ;
    END
  END slave3_wb_data_i[3]
  PIN slave3_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 239.400 350.000 240.000 ;
    END
  END slave3_wb_data_i[4]
  PIN slave3_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 270.000 350.000 270.600 ;
    END
  END slave3_wb_data_i[5]
  PIN slave3_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 300.600 350.000 301.200 ;
    END
  END slave3_wb_data_i[6]
  PIN slave3_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 331.200 350.000 331.800 ;
    END
  END slave3_wb_data_i[7]
  PIN slave3_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 361.800 350.000 362.400 ;
    END
  END slave3_wb_data_i[8]
  PIN slave3_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 392.400 350.000 393.000 ;
    END
  END slave3_wb_data_i[9]
  PIN slave3_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 86.400 350.000 87.000 ;
    END
  END slave3_wb_data_o[0]
  PIN slave3_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 433.200 350.000 433.800 ;
    END
  END slave3_wb_data_o[10]
  PIN slave3_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 463.800 350.000 464.400 ;
    END
  END slave3_wb_data_o[11]
  PIN slave3_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 494.400 350.000 495.000 ;
    END
  END slave3_wb_data_o[12]
  PIN slave3_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 525.000 350.000 525.600 ;
    END
  END slave3_wb_data_o[13]
  PIN slave3_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 555.600 350.000 556.200 ;
    END
  END slave3_wb_data_o[14]
  PIN slave3_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 586.200 350.000 586.800 ;
    END
  END slave3_wb_data_o[15]
  PIN slave3_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 616.800 350.000 617.400 ;
    END
  END slave3_wb_data_o[16]
  PIN slave3_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 647.400 350.000 648.000 ;
    END
  END slave3_wb_data_o[17]
  PIN slave3_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 678.000 350.000 678.600 ;
    END
  END slave3_wb_data_o[18]
  PIN slave3_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 708.600 350.000 709.200 ;
    END
  END slave3_wb_data_o[19]
  PIN slave3_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 127.200 350.000 127.800 ;
    END
  END slave3_wb_data_o[1]
  PIN slave3_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 739.200 350.000 739.800 ;
    END
  END slave3_wb_data_o[20]
  PIN slave3_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 769.800 350.000 770.400 ;
    END
  END slave3_wb_data_o[21]
  PIN slave3_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 800.400 350.000 801.000 ;
    END
  END slave3_wb_data_o[22]
  PIN slave3_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 831.000 350.000 831.600 ;
    END
  END slave3_wb_data_o[23]
  PIN slave3_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 851.400 350.000 852.000 ;
    END
  END slave3_wb_data_o[24]
  PIN slave3_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 871.800 350.000 872.400 ;
    END
  END slave3_wb_data_o[25]
  PIN slave3_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 892.200 350.000 892.800 ;
    END
  END slave3_wb_data_o[26]
  PIN slave3_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 912.600 350.000 913.200 ;
    END
  END slave3_wb_data_o[27]
  PIN slave3_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 933.000 350.000 933.600 ;
    END
  END slave3_wb_data_o[28]
  PIN slave3_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 953.400 350.000 954.000 ;
    END
  END slave3_wb_data_o[29]
  PIN slave3_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 168.000 350.000 168.600 ;
    END
  END slave3_wb_data_o[2]
  PIN slave3_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 973.800 350.000 974.400 ;
    END
  END slave3_wb_data_o[30]
  PIN slave3_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 994.200 350.000 994.800 ;
    END
  END slave3_wb_data_o[31]
  PIN slave3_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 208.800 350.000 209.400 ;
    END
  END slave3_wb_data_o[3]
  PIN slave3_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 249.600 350.000 250.200 ;
    END
  END slave3_wb_data_o[4]
  PIN slave3_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 280.200 350.000 280.800 ;
    END
  END slave3_wb_data_o[5]
  PIN slave3_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 310.800 350.000 311.400 ;
    END
  END slave3_wb_data_o[6]
  PIN slave3_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 341.400 350.000 342.000 ;
    END
  END slave3_wb_data_o[7]
  PIN slave3_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 372.000 350.000 372.600 ;
    END
  END slave3_wb_data_o[8]
  PIN slave3_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 402.600 350.000 403.200 ;
    END
  END slave3_wb_data_o[9]
  PIN slave3_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 25.200 350.000 25.800 ;
    END
  END slave3_wb_error_o
  PIN slave3_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 96.600 350.000 97.200 ;
    END
  END slave3_wb_sel_i[0]
  PIN slave3_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 137.400 350.000 138.000 ;
    END
  END slave3_wb_sel_i[1]
  PIN slave3_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 178.200 350.000 178.800 ;
    END
  END slave3_wb_sel_i[2]
  PIN slave3_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 219.000 350.000 219.600 ;
    END
  END slave3_wb_sel_i[3]
  PIN slave3_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 35.400 350.000 36.000 ;
    END
  END slave3_wb_stall_o
  PIN slave3_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 45.600 350.000 46.200 ;
    END
  END slave3_wb_stb_i
  PIN slave3_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 55.800 350.000 56.400 ;
    END
  END slave3_wb_we_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 987.600 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 987.445 ;
      LAYER met1 ;
        RECT 1.450 9.560 348.610 987.600 ;
      LAYER met2 ;
        RECT 2.030 995.720 4.410 998.765 ;
        RECT 5.250 995.720 8.090 998.765 ;
        RECT 8.930 995.720 11.770 998.765 ;
        RECT 12.610 995.720 15.450 998.765 ;
        RECT 16.290 995.720 18.670 998.765 ;
        RECT 19.510 995.720 22.350 998.765 ;
        RECT 23.190 995.720 26.030 998.765 ;
        RECT 26.870 995.720 29.710 998.765 ;
        RECT 30.550 995.720 32.930 998.765 ;
        RECT 33.770 995.720 36.610 998.765 ;
        RECT 37.450 995.720 40.290 998.765 ;
        RECT 41.130 995.720 43.970 998.765 ;
        RECT 44.810 995.720 47.190 998.765 ;
        RECT 48.030 995.720 50.870 998.765 ;
        RECT 51.710 995.720 54.550 998.765 ;
        RECT 55.390 995.720 58.230 998.765 ;
        RECT 59.070 995.720 61.910 998.765 ;
        RECT 62.750 995.720 65.130 998.765 ;
        RECT 65.970 995.720 68.810 998.765 ;
        RECT 69.650 995.720 72.490 998.765 ;
        RECT 73.330 995.720 76.170 998.765 ;
        RECT 77.010 995.720 79.390 998.765 ;
        RECT 80.230 995.720 83.070 998.765 ;
        RECT 83.910 995.720 86.750 998.765 ;
        RECT 87.590 995.720 90.430 998.765 ;
        RECT 91.270 995.720 93.650 998.765 ;
        RECT 94.490 995.720 97.330 998.765 ;
        RECT 98.170 995.720 101.010 998.765 ;
        RECT 101.850 995.720 104.690 998.765 ;
        RECT 105.530 995.720 107.910 998.765 ;
        RECT 108.750 995.720 111.590 998.765 ;
        RECT 112.430 995.720 115.270 998.765 ;
        RECT 116.110 995.720 118.950 998.765 ;
        RECT 119.790 995.720 122.630 998.765 ;
        RECT 123.470 995.720 125.850 998.765 ;
        RECT 126.690 995.720 129.530 998.765 ;
        RECT 130.370 995.720 133.210 998.765 ;
        RECT 134.050 995.720 136.890 998.765 ;
        RECT 137.730 995.720 140.110 998.765 ;
        RECT 140.950 995.720 143.790 998.765 ;
        RECT 144.630 995.720 147.470 998.765 ;
        RECT 148.310 995.720 151.150 998.765 ;
        RECT 151.990 995.720 154.370 998.765 ;
        RECT 155.210 995.720 158.050 998.765 ;
        RECT 158.890 995.720 161.730 998.765 ;
        RECT 162.570 995.720 165.410 998.765 ;
        RECT 166.250 995.720 168.630 998.765 ;
        RECT 169.470 995.720 172.310 998.765 ;
        RECT 173.150 995.720 175.990 998.765 ;
        RECT 176.830 995.720 179.670 998.765 ;
        RECT 180.510 995.720 183.350 998.765 ;
        RECT 184.190 995.720 186.570 998.765 ;
        RECT 187.410 995.720 190.250 998.765 ;
        RECT 191.090 995.720 193.930 998.765 ;
        RECT 194.770 995.720 197.610 998.765 ;
        RECT 198.450 995.720 200.830 998.765 ;
        RECT 201.670 995.720 204.510 998.765 ;
        RECT 205.350 995.720 208.190 998.765 ;
        RECT 209.030 995.720 211.870 998.765 ;
        RECT 212.710 995.720 215.090 998.765 ;
        RECT 215.930 995.720 218.770 998.765 ;
        RECT 219.610 995.720 222.450 998.765 ;
        RECT 223.290 995.720 226.130 998.765 ;
        RECT 226.970 995.720 229.350 998.765 ;
        RECT 230.190 995.720 233.030 998.765 ;
        RECT 233.870 995.720 236.710 998.765 ;
        RECT 237.550 995.720 240.390 998.765 ;
        RECT 241.230 995.720 244.070 998.765 ;
        RECT 244.910 995.720 247.290 998.765 ;
        RECT 248.130 995.720 250.970 998.765 ;
        RECT 251.810 995.720 254.650 998.765 ;
        RECT 255.490 995.720 258.330 998.765 ;
        RECT 259.170 995.720 261.550 998.765 ;
        RECT 262.390 995.720 265.230 998.765 ;
        RECT 266.070 995.720 268.910 998.765 ;
        RECT 269.750 995.720 272.590 998.765 ;
        RECT 273.430 995.720 275.810 998.765 ;
        RECT 276.650 995.720 279.490 998.765 ;
        RECT 280.330 995.720 283.170 998.765 ;
        RECT 284.010 995.720 286.850 998.765 ;
        RECT 287.690 995.720 290.070 998.765 ;
        RECT 290.910 995.720 293.750 998.765 ;
        RECT 294.590 995.720 297.430 998.765 ;
        RECT 298.270 995.720 301.110 998.765 ;
        RECT 301.950 995.720 304.790 998.765 ;
        RECT 305.630 995.720 308.010 998.765 ;
        RECT 308.850 995.720 311.690 998.765 ;
        RECT 312.530 995.720 315.370 998.765 ;
        RECT 316.210 995.720 319.050 998.765 ;
        RECT 319.890 995.720 322.270 998.765 ;
        RECT 323.110 995.720 325.950 998.765 ;
        RECT 326.790 995.720 329.630 998.765 ;
        RECT 330.470 995.720 333.310 998.765 ;
        RECT 334.150 995.720 336.530 998.765 ;
        RECT 337.370 995.720 340.210 998.765 ;
        RECT 341.050 995.720 343.890 998.765 ;
        RECT 344.730 995.720 347.570 998.765 ;
        RECT 348.410 995.720 348.580 998.765 ;
        RECT 1.480 4.280 348.580 995.720 ;
        RECT 2.030 0.835 3.950 4.280 ;
        RECT 4.790 0.835 6.710 4.280 ;
        RECT 7.550 0.835 9.930 4.280 ;
        RECT 10.770 0.835 12.690 4.280 ;
        RECT 13.530 0.835 15.450 4.280 ;
        RECT 16.290 0.835 18.670 4.280 ;
        RECT 19.510 0.835 21.430 4.280 ;
        RECT 22.270 0.835 24.190 4.280 ;
        RECT 25.030 0.835 27.410 4.280 ;
        RECT 28.250 0.835 30.170 4.280 ;
        RECT 31.010 0.835 32.930 4.280 ;
        RECT 33.770 0.835 36.150 4.280 ;
        RECT 36.990 0.835 38.910 4.280 ;
        RECT 39.750 0.835 41.670 4.280 ;
        RECT 42.510 0.835 44.890 4.280 ;
        RECT 45.730 0.835 47.650 4.280 ;
        RECT 48.490 0.835 50.410 4.280 ;
        RECT 51.250 0.835 53.630 4.280 ;
        RECT 54.470 0.835 56.390 4.280 ;
        RECT 57.230 0.835 59.150 4.280 ;
        RECT 59.990 0.835 62.370 4.280 ;
        RECT 63.210 0.835 65.130 4.280 ;
        RECT 65.970 0.835 67.890 4.280 ;
        RECT 68.730 0.835 71.110 4.280 ;
        RECT 71.950 0.835 73.870 4.280 ;
        RECT 74.710 0.835 76.630 4.280 ;
        RECT 77.470 0.835 79.850 4.280 ;
        RECT 80.690 0.835 82.610 4.280 ;
        RECT 83.450 0.835 85.370 4.280 ;
        RECT 86.210 0.835 88.590 4.280 ;
        RECT 89.430 0.835 91.350 4.280 ;
        RECT 92.190 0.835 94.110 4.280 ;
        RECT 94.950 0.835 97.330 4.280 ;
        RECT 98.170 0.835 100.090 4.280 ;
        RECT 100.930 0.835 102.850 4.280 ;
        RECT 103.690 0.835 106.070 4.280 ;
        RECT 106.910 0.835 108.830 4.280 ;
        RECT 109.670 0.835 111.590 4.280 ;
        RECT 112.430 0.835 114.810 4.280 ;
        RECT 115.650 0.835 117.570 4.280 ;
        RECT 118.410 0.835 120.790 4.280 ;
        RECT 121.630 0.835 123.550 4.280 ;
        RECT 124.390 0.835 126.310 4.280 ;
        RECT 127.150 0.835 129.530 4.280 ;
        RECT 130.370 0.835 132.290 4.280 ;
        RECT 133.130 0.835 135.050 4.280 ;
        RECT 135.890 0.835 138.270 4.280 ;
        RECT 139.110 0.835 141.030 4.280 ;
        RECT 141.870 0.835 143.790 4.280 ;
        RECT 144.630 0.835 147.010 4.280 ;
        RECT 147.850 0.835 149.770 4.280 ;
        RECT 150.610 0.835 152.530 4.280 ;
        RECT 153.370 0.835 155.750 4.280 ;
        RECT 156.590 0.835 158.510 4.280 ;
        RECT 159.350 0.835 161.270 4.280 ;
        RECT 162.110 0.835 164.490 4.280 ;
        RECT 165.330 0.835 167.250 4.280 ;
        RECT 168.090 0.835 170.010 4.280 ;
        RECT 170.850 0.835 173.230 4.280 ;
        RECT 174.070 0.835 175.990 4.280 ;
        RECT 176.830 0.835 178.750 4.280 ;
        RECT 179.590 0.835 181.970 4.280 ;
        RECT 182.810 0.835 184.730 4.280 ;
        RECT 185.570 0.835 187.490 4.280 ;
        RECT 188.330 0.835 190.710 4.280 ;
        RECT 191.550 0.835 193.470 4.280 ;
        RECT 194.310 0.835 196.230 4.280 ;
        RECT 197.070 0.835 199.450 4.280 ;
        RECT 200.290 0.835 202.210 4.280 ;
        RECT 203.050 0.835 204.970 4.280 ;
        RECT 205.810 0.835 208.190 4.280 ;
        RECT 209.030 0.835 210.950 4.280 ;
        RECT 211.790 0.835 213.710 4.280 ;
        RECT 214.550 0.835 216.930 4.280 ;
        RECT 217.770 0.835 219.690 4.280 ;
        RECT 220.530 0.835 222.450 4.280 ;
        RECT 223.290 0.835 225.670 4.280 ;
        RECT 226.510 0.835 228.430 4.280 ;
        RECT 229.270 0.835 231.190 4.280 ;
        RECT 232.030 0.835 234.410 4.280 ;
        RECT 235.250 0.835 237.170 4.280 ;
        RECT 238.010 0.835 240.390 4.280 ;
        RECT 241.230 0.835 243.150 4.280 ;
        RECT 243.990 0.835 245.910 4.280 ;
        RECT 246.750 0.835 249.130 4.280 ;
        RECT 249.970 0.835 251.890 4.280 ;
        RECT 252.730 0.835 254.650 4.280 ;
        RECT 255.490 0.835 257.870 4.280 ;
        RECT 258.710 0.835 260.630 4.280 ;
        RECT 261.470 0.835 263.390 4.280 ;
        RECT 264.230 0.835 266.610 4.280 ;
        RECT 267.450 0.835 269.370 4.280 ;
        RECT 270.210 0.835 272.130 4.280 ;
        RECT 272.970 0.835 275.350 4.280 ;
        RECT 276.190 0.835 278.110 4.280 ;
        RECT 278.950 0.835 280.870 4.280 ;
        RECT 281.710 0.835 284.090 4.280 ;
        RECT 284.930 0.835 286.850 4.280 ;
        RECT 287.690 0.835 289.610 4.280 ;
        RECT 290.450 0.835 292.830 4.280 ;
        RECT 293.670 0.835 295.590 4.280 ;
        RECT 296.430 0.835 298.350 4.280 ;
        RECT 299.190 0.835 301.570 4.280 ;
        RECT 302.410 0.835 304.330 4.280 ;
        RECT 305.170 0.835 307.090 4.280 ;
        RECT 307.930 0.835 310.310 4.280 ;
        RECT 311.150 0.835 313.070 4.280 ;
        RECT 313.910 0.835 315.830 4.280 ;
        RECT 316.670 0.835 319.050 4.280 ;
        RECT 319.890 0.835 321.810 4.280 ;
        RECT 322.650 0.835 324.570 4.280 ;
        RECT 325.410 0.835 327.790 4.280 ;
        RECT 328.630 0.835 330.550 4.280 ;
        RECT 331.390 0.835 333.310 4.280 ;
        RECT 334.150 0.835 336.530 4.280 ;
        RECT 337.370 0.835 339.290 4.280 ;
        RECT 340.130 0.835 342.050 4.280 ;
        RECT 342.890 0.835 345.270 4.280 ;
        RECT 346.110 0.835 348.030 4.280 ;
      LAYER met3 ;
        RECT 4.400 997.880 346.000 998.745 ;
        RECT 1.905 996.560 346.000 997.880 ;
        RECT 4.400 995.200 346.000 996.560 ;
        RECT 4.400 995.160 345.600 995.200 ;
        RECT 1.905 993.840 345.600 995.160 ;
        RECT 4.400 993.800 345.600 993.840 ;
        RECT 4.400 992.440 346.000 993.800 ;
        RECT 1.905 991.800 346.000 992.440 ;
        RECT 4.400 990.400 346.000 991.800 ;
        RECT 1.905 989.080 346.000 990.400 ;
        RECT 4.400 987.680 346.000 989.080 ;
        RECT 1.905 986.360 346.000 987.680 ;
        RECT 4.400 985.000 346.000 986.360 ;
        RECT 4.400 984.960 345.600 985.000 ;
        RECT 1.905 984.320 345.600 984.960 ;
        RECT 4.400 983.600 345.600 984.320 ;
        RECT 4.400 982.920 346.000 983.600 ;
        RECT 1.905 981.600 346.000 982.920 ;
        RECT 4.400 980.200 346.000 981.600 ;
        RECT 1.905 978.880 346.000 980.200 ;
        RECT 4.400 977.480 346.000 978.880 ;
        RECT 1.905 976.840 346.000 977.480 ;
        RECT 4.400 975.440 346.000 976.840 ;
        RECT 1.905 974.800 346.000 975.440 ;
        RECT 1.905 974.120 345.600 974.800 ;
        RECT 4.400 973.400 345.600 974.120 ;
        RECT 4.400 972.720 346.000 973.400 ;
        RECT 1.905 971.400 346.000 972.720 ;
        RECT 4.400 970.000 346.000 971.400 ;
        RECT 1.905 969.360 346.000 970.000 ;
        RECT 4.400 967.960 346.000 969.360 ;
        RECT 1.905 966.640 346.000 967.960 ;
        RECT 4.400 965.240 346.000 966.640 ;
        RECT 1.905 964.600 346.000 965.240 ;
        RECT 1.905 963.920 345.600 964.600 ;
        RECT 4.400 963.200 345.600 963.920 ;
        RECT 4.400 962.520 346.000 963.200 ;
        RECT 1.905 961.880 346.000 962.520 ;
        RECT 4.400 960.480 346.000 961.880 ;
        RECT 1.905 959.160 346.000 960.480 ;
        RECT 4.400 957.760 346.000 959.160 ;
        RECT 1.905 956.440 346.000 957.760 ;
        RECT 4.400 955.040 346.000 956.440 ;
        RECT 1.905 954.400 346.000 955.040 ;
        RECT 4.400 953.000 345.600 954.400 ;
        RECT 1.905 951.680 346.000 953.000 ;
        RECT 4.400 950.280 346.000 951.680 ;
        RECT 1.905 948.960 346.000 950.280 ;
        RECT 4.400 947.560 346.000 948.960 ;
        RECT 1.905 946.920 346.000 947.560 ;
        RECT 4.400 945.520 346.000 946.920 ;
        RECT 1.905 944.200 346.000 945.520 ;
        RECT 4.400 942.800 345.600 944.200 ;
        RECT 1.905 941.480 346.000 942.800 ;
        RECT 4.400 940.080 346.000 941.480 ;
        RECT 1.905 939.440 346.000 940.080 ;
        RECT 4.400 938.040 346.000 939.440 ;
        RECT 1.905 936.720 346.000 938.040 ;
        RECT 4.400 935.320 346.000 936.720 ;
        RECT 1.905 934.000 346.000 935.320 ;
        RECT 4.400 932.600 345.600 934.000 ;
        RECT 1.905 931.960 346.000 932.600 ;
        RECT 4.400 930.560 346.000 931.960 ;
        RECT 1.905 929.240 346.000 930.560 ;
        RECT 4.400 927.840 346.000 929.240 ;
        RECT 1.905 926.520 346.000 927.840 ;
        RECT 4.400 925.120 346.000 926.520 ;
        RECT 1.905 923.800 346.000 925.120 ;
        RECT 4.400 922.400 345.600 923.800 ;
        RECT 1.905 921.760 346.000 922.400 ;
        RECT 4.400 920.360 346.000 921.760 ;
        RECT 1.905 919.040 346.000 920.360 ;
        RECT 4.400 917.640 346.000 919.040 ;
        RECT 1.905 916.320 346.000 917.640 ;
        RECT 4.400 914.920 346.000 916.320 ;
        RECT 1.905 914.280 346.000 914.920 ;
        RECT 4.400 913.600 346.000 914.280 ;
        RECT 4.400 912.880 345.600 913.600 ;
        RECT 1.905 912.200 345.600 912.880 ;
        RECT 1.905 911.560 346.000 912.200 ;
        RECT 4.400 910.160 346.000 911.560 ;
        RECT 1.905 908.840 346.000 910.160 ;
        RECT 4.400 907.440 346.000 908.840 ;
        RECT 1.905 906.800 346.000 907.440 ;
        RECT 4.400 905.400 346.000 906.800 ;
        RECT 1.905 904.080 346.000 905.400 ;
        RECT 4.400 903.400 346.000 904.080 ;
        RECT 4.400 902.680 345.600 903.400 ;
        RECT 1.905 902.000 345.600 902.680 ;
        RECT 1.905 901.360 346.000 902.000 ;
        RECT 4.400 899.960 346.000 901.360 ;
        RECT 1.905 899.320 346.000 899.960 ;
        RECT 4.400 897.920 346.000 899.320 ;
        RECT 1.905 896.600 346.000 897.920 ;
        RECT 4.400 895.200 346.000 896.600 ;
        RECT 1.905 893.880 346.000 895.200 ;
        RECT 4.400 893.200 346.000 893.880 ;
        RECT 4.400 892.480 345.600 893.200 ;
        RECT 1.905 891.840 345.600 892.480 ;
        RECT 4.400 891.800 345.600 891.840 ;
        RECT 4.400 890.440 346.000 891.800 ;
        RECT 1.905 889.120 346.000 890.440 ;
        RECT 4.400 887.720 346.000 889.120 ;
        RECT 1.905 886.400 346.000 887.720 ;
        RECT 4.400 885.000 346.000 886.400 ;
        RECT 1.905 884.360 346.000 885.000 ;
        RECT 4.400 883.000 346.000 884.360 ;
        RECT 4.400 882.960 345.600 883.000 ;
        RECT 1.905 881.640 345.600 882.960 ;
        RECT 4.400 881.600 345.600 881.640 ;
        RECT 4.400 880.240 346.000 881.600 ;
        RECT 1.905 878.920 346.000 880.240 ;
        RECT 4.400 877.520 346.000 878.920 ;
        RECT 1.905 876.880 346.000 877.520 ;
        RECT 4.400 875.480 346.000 876.880 ;
        RECT 1.905 874.160 346.000 875.480 ;
        RECT 4.400 872.800 346.000 874.160 ;
        RECT 4.400 872.760 345.600 872.800 ;
        RECT 1.905 871.440 345.600 872.760 ;
        RECT 4.400 871.400 345.600 871.440 ;
        RECT 4.400 870.040 346.000 871.400 ;
        RECT 1.905 869.400 346.000 870.040 ;
        RECT 4.400 868.000 346.000 869.400 ;
        RECT 1.905 866.680 346.000 868.000 ;
        RECT 4.400 865.280 346.000 866.680 ;
        RECT 1.905 863.960 346.000 865.280 ;
        RECT 4.400 862.600 346.000 863.960 ;
        RECT 4.400 862.560 345.600 862.600 ;
        RECT 1.905 861.920 345.600 862.560 ;
        RECT 4.400 861.200 345.600 861.920 ;
        RECT 4.400 860.520 346.000 861.200 ;
        RECT 1.905 859.200 346.000 860.520 ;
        RECT 4.400 857.800 346.000 859.200 ;
        RECT 1.905 856.480 346.000 857.800 ;
        RECT 4.400 855.080 346.000 856.480 ;
        RECT 1.905 854.440 346.000 855.080 ;
        RECT 4.400 853.040 346.000 854.440 ;
        RECT 1.905 852.400 346.000 853.040 ;
        RECT 1.905 851.720 345.600 852.400 ;
        RECT 4.400 851.000 345.600 851.720 ;
        RECT 4.400 850.320 346.000 851.000 ;
        RECT 1.905 849.000 346.000 850.320 ;
        RECT 4.400 847.600 346.000 849.000 ;
        RECT 1.905 846.280 346.000 847.600 ;
        RECT 4.400 844.880 346.000 846.280 ;
        RECT 1.905 844.240 346.000 844.880 ;
        RECT 4.400 842.840 346.000 844.240 ;
        RECT 1.905 842.200 346.000 842.840 ;
        RECT 1.905 841.520 345.600 842.200 ;
        RECT 4.400 840.800 345.600 841.520 ;
        RECT 4.400 840.120 346.000 840.800 ;
        RECT 1.905 838.800 346.000 840.120 ;
        RECT 4.400 837.400 346.000 838.800 ;
        RECT 1.905 836.760 346.000 837.400 ;
        RECT 4.400 835.360 346.000 836.760 ;
        RECT 1.905 834.040 346.000 835.360 ;
        RECT 4.400 832.640 346.000 834.040 ;
        RECT 1.905 832.000 346.000 832.640 ;
        RECT 1.905 831.320 345.600 832.000 ;
        RECT 4.400 830.600 345.600 831.320 ;
        RECT 4.400 829.920 346.000 830.600 ;
        RECT 1.905 829.280 346.000 829.920 ;
        RECT 4.400 827.880 346.000 829.280 ;
        RECT 1.905 826.560 346.000 827.880 ;
        RECT 4.400 825.160 346.000 826.560 ;
        RECT 1.905 823.840 346.000 825.160 ;
        RECT 4.400 822.440 346.000 823.840 ;
        RECT 1.905 821.800 346.000 822.440 ;
        RECT 4.400 820.400 345.600 821.800 ;
        RECT 1.905 819.080 346.000 820.400 ;
        RECT 4.400 817.680 346.000 819.080 ;
        RECT 1.905 816.360 346.000 817.680 ;
        RECT 4.400 814.960 346.000 816.360 ;
        RECT 1.905 814.320 346.000 814.960 ;
        RECT 4.400 812.920 346.000 814.320 ;
        RECT 1.905 811.600 346.000 812.920 ;
        RECT 4.400 810.200 345.600 811.600 ;
        RECT 1.905 808.880 346.000 810.200 ;
        RECT 4.400 807.480 346.000 808.880 ;
        RECT 1.905 806.840 346.000 807.480 ;
        RECT 4.400 805.440 346.000 806.840 ;
        RECT 1.905 804.120 346.000 805.440 ;
        RECT 4.400 802.720 346.000 804.120 ;
        RECT 1.905 801.400 346.000 802.720 ;
        RECT 4.400 800.000 345.600 801.400 ;
        RECT 1.905 799.360 346.000 800.000 ;
        RECT 4.400 797.960 346.000 799.360 ;
        RECT 1.905 796.640 346.000 797.960 ;
        RECT 4.400 795.240 346.000 796.640 ;
        RECT 1.905 793.920 346.000 795.240 ;
        RECT 4.400 792.520 346.000 793.920 ;
        RECT 1.905 791.880 346.000 792.520 ;
        RECT 4.400 791.200 346.000 791.880 ;
        RECT 4.400 790.480 345.600 791.200 ;
        RECT 1.905 789.800 345.600 790.480 ;
        RECT 1.905 789.160 346.000 789.800 ;
        RECT 4.400 787.760 346.000 789.160 ;
        RECT 1.905 786.440 346.000 787.760 ;
        RECT 4.400 785.040 346.000 786.440 ;
        RECT 1.905 784.400 346.000 785.040 ;
        RECT 4.400 783.000 346.000 784.400 ;
        RECT 1.905 781.680 346.000 783.000 ;
        RECT 4.400 781.000 346.000 781.680 ;
        RECT 4.400 780.280 345.600 781.000 ;
        RECT 1.905 779.600 345.600 780.280 ;
        RECT 1.905 778.960 346.000 779.600 ;
        RECT 4.400 777.560 346.000 778.960 ;
        RECT 1.905 776.920 346.000 777.560 ;
        RECT 4.400 775.520 346.000 776.920 ;
        RECT 1.905 774.200 346.000 775.520 ;
        RECT 4.400 772.800 346.000 774.200 ;
        RECT 1.905 771.480 346.000 772.800 ;
        RECT 4.400 770.800 346.000 771.480 ;
        RECT 4.400 770.080 345.600 770.800 ;
        RECT 1.905 769.400 345.600 770.080 ;
        RECT 1.905 768.760 346.000 769.400 ;
        RECT 4.400 767.360 346.000 768.760 ;
        RECT 1.905 766.720 346.000 767.360 ;
        RECT 4.400 765.320 346.000 766.720 ;
        RECT 1.905 764.000 346.000 765.320 ;
        RECT 4.400 762.600 346.000 764.000 ;
        RECT 1.905 761.280 346.000 762.600 ;
        RECT 4.400 760.600 346.000 761.280 ;
        RECT 4.400 759.880 345.600 760.600 ;
        RECT 1.905 759.240 345.600 759.880 ;
        RECT 4.400 759.200 345.600 759.240 ;
        RECT 4.400 757.840 346.000 759.200 ;
        RECT 1.905 756.520 346.000 757.840 ;
        RECT 4.400 755.120 346.000 756.520 ;
        RECT 1.905 753.800 346.000 755.120 ;
        RECT 4.400 752.400 346.000 753.800 ;
        RECT 1.905 751.760 346.000 752.400 ;
        RECT 4.400 750.400 346.000 751.760 ;
        RECT 4.400 750.360 345.600 750.400 ;
        RECT 1.905 749.040 345.600 750.360 ;
        RECT 4.400 749.000 345.600 749.040 ;
        RECT 4.400 747.640 346.000 749.000 ;
        RECT 1.905 746.320 346.000 747.640 ;
        RECT 4.400 744.920 346.000 746.320 ;
        RECT 1.905 744.280 346.000 744.920 ;
        RECT 4.400 742.880 346.000 744.280 ;
        RECT 1.905 741.560 346.000 742.880 ;
        RECT 4.400 740.200 346.000 741.560 ;
        RECT 4.400 740.160 345.600 740.200 ;
        RECT 1.905 738.840 345.600 740.160 ;
        RECT 4.400 738.800 345.600 738.840 ;
        RECT 4.400 737.440 346.000 738.800 ;
        RECT 1.905 736.800 346.000 737.440 ;
        RECT 4.400 735.400 346.000 736.800 ;
        RECT 1.905 734.080 346.000 735.400 ;
        RECT 4.400 732.680 346.000 734.080 ;
        RECT 1.905 731.360 346.000 732.680 ;
        RECT 4.400 730.000 346.000 731.360 ;
        RECT 4.400 729.960 345.600 730.000 ;
        RECT 1.905 729.320 345.600 729.960 ;
        RECT 4.400 728.600 345.600 729.320 ;
        RECT 4.400 727.920 346.000 728.600 ;
        RECT 1.905 726.600 346.000 727.920 ;
        RECT 4.400 725.200 346.000 726.600 ;
        RECT 1.905 723.880 346.000 725.200 ;
        RECT 4.400 722.480 346.000 723.880 ;
        RECT 1.905 721.840 346.000 722.480 ;
        RECT 4.400 720.440 346.000 721.840 ;
        RECT 1.905 719.800 346.000 720.440 ;
        RECT 1.905 719.120 345.600 719.800 ;
        RECT 4.400 718.400 345.600 719.120 ;
        RECT 4.400 717.720 346.000 718.400 ;
        RECT 1.905 716.400 346.000 717.720 ;
        RECT 4.400 715.000 346.000 716.400 ;
        RECT 1.905 714.360 346.000 715.000 ;
        RECT 4.400 712.960 346.000 714.360 ;
        RECT 1.905 711.640 346.000 712.960 ;
        RECT 4.400 710.240 346.000 711.640 ;
        RECT 1.905 709.600 346.000 710.240 ;
        RECT 1.905 708.920 345.600 709.600 ;
        RECT 4.400 708.200 345.600 708.920 ;
        RECT 4.400 707.520 346.000 708.200 ;
        RECT 1.905 706.880 346.000 707.520 ;
        RECT 4.400 705.480 346.000 706.880 ;
        RECT 1.905 704.160 346.000 705.480 ;
        RECT 4.400 702.760 346.000 704.160 ;
        RECT 1.905 701.440 346.000 702.760 ;
        RECT 4.400 700.040 346.000 701.440 ;
        RECT 1.905 699.400 346.000 700.040 ;
        RECT 4.400 698.000 345.600 699.400 ;
        RECT 1.905 696.680 346.000 698.000 ;
        RECT 4.400 695.280 346.000 696.680 ;
        RECT 1.905 693.960 346.000 695.280 ;
        RECT 4.400 692.560 346.000 693.960 ;
        RECT 1.905 691.240 346.000 692.560 ;
        RECT 4.400 689.840 346.000 691.240 ;
        RECT 1.905 689.200 346.000 689.840 ;
        RECT 4.400 687.800 345.600 689.200 ;
        RECT 1.905 686.480 346.000 687.800 ;
        RECT 4.400 685.080 346.000 686.480 ;
        RECT 1.905 683.760 346.000 685.080 ;
        RECT 4.400 682.360 346.000 683.760 ;
        RECT 1.905 681.720 346.000 682.360 ;
        RECT 4.400 680.320 346.000 681.720 ;
        RECT 1.905 679.000 346.000 680.320 ;
        RECT 4.400 677.600 345.600 679.000 ;
        RECT 1.905 676.280 346.000 677.600 ;
        RECT 4.400 674.880 346.000 676.280 ;
        RECT 1.905 674.240 346.000 674.880 ;
        RECT 4.400 672.840 346.000 674.240 ;
        RECT 1.905 671.520 346.000 672.840 ;
        RECT 4.400 670.120 346.000 671.520 ;
        RECT 1.905 668.800 346.000 670.120 ;
        RECT 4.400 667.400 345.600 668.800 ;
        RECT 1.905 666.760 346.000 667.400 ;
        RECT 4.400 665.360 346.000 666.760 ;
        RECT 1.905 664.040 346.000 665.360 ;
        RECT 4.400 662.640 346.000 664.040 ;
        RECT 1.905 661.320 346.000 662.640 ;
        RECT 4.400 659.920 346.000 661.320 ;
        RECT 1.905 659.280 346.000 659.920 ;
        RECT 4.400 658.600 346.000 659.280 ;
        RECT 4.400 657.880 345.600 658.600 ;
        RECT 1.905 657.200 345.600 657.880 ;
        RECT 1.905 656.560 346.000 657.200 ;
        RECT 4.400 655.160 346.000 656.560 ;
        RECT 1.905 653.840 346.000 655.160 ;
        RECT 4.400 652.440 346.000 653.840 ;
        RECT 1.905 651.800 346.000 652.440 ;
        RECT 4.400 650.400 346.000 651.800 ;
        RECT 1.905 649.080 346.000 650.400 ;
        RECT 4.400 648.400 346.000 649.080 ;
        RECT 4.400 647.680 345.600 648.400 ;
        RECT 1.905 647.000 345.600 647.680 ;
        RECT 1.905 646.360 346.000 647.000 ;
        RECT 4.400 644.960 346.000 646.360 ;
        RECT 1.905 644.320 346.000 644.960 ;
        RECT 4.400 642.920 346.000 644.320 ;
        RECT 1.905 641.600 346.000 642.920 ;
        RECT 4.400 640.200 346.000 641.600 ;
        RECT 1.905 638.880 346.000 640.200 ;
        RECT 4.400 638.200 346.000 638.880 ;
        RECT 4.400 637.480 345.600 638.200 ;
        RECT 1.905 636.840 345.600 637.480 ;
        RECT 4.400 636.800 345.600 636.840 ;
        RECT 4.400 635.440 346.000 636.800 ;
        RECT 1.905 634.120 346.000 635.440 ;
        RECT 4.400 632.720 346.000 634.120 ;
        RECT 1.905 631.400 346.000 632.720 ;
        RECT 4.400 630.000 346.000 631.400 ;
        RECT 1.905 629.360 346.000 630.000 ;
        RECT 4.400 628.000 346.000 629.360 ;
        RECT 4.400 627.960 345.600 628.000 ;
        RECT 1.905 626.640 345.600 627.960 ;
        RECT 4.400 626.600 345.600 626.640 ;
        RECT 4.400 625.240 346.000 626.600 ;
        RECT 1.905 623.920 346.000 625.240 ;
        RECT 4.400 622.520 346.000 623.920 ;
        RECT 1.905 621.880 346.000 622.520 ;
        RECT 4.400 620.480 346.000 621.880 ;
        RECT 1.905 619.160 346.000 620.480 ;
        RECT 4.400 617.800 346.000 619.160 ;
        RECT 4.400 617.760 345.600 617.800 ;
        RECT 1.905 616.440 345.600 617.760 ;
        RECT 4.400 616.400 345.600 616.440 ;
        RECT 4.400 615.040 346.000 616.400 ;
        RECT 1.905 613.720 346.000 615.040 ;
        RECT 4.400 612.320 346.000 613.720 ;
        RECT 1.905 611.680 346.000 612.320 ;
        RECT 4.400 610.280 346.000 611.680 ;
        RECT 1.905 608.960 346.000 610.280 ;
        RECT 4.400 607.600 346.000 608.960 ;
        RECT 4.400 607.560 345.600 607.600 ;
        RECT 1.905 606.240 345.600 607.560 ;
        RECT 4.400 606.200 345.600 606.240 ;
        RECT 4.400 604.840 346.000 606.200 ;
        RECT 1.905 604.200 346.000 604.840 ;
        RECT 4.400 602.800 346.000 604.200 ;
        RECT 1.905 601.480 346.000 602.800 ;
        RECT 4.400 600.080 346.000 601.480 ;
        RECT 1.905 598.760 346.000 600.080 ;
        RECT 4.400 597.400 346.000 598.760 ;
        RECT 4.400 597.360 345.600 597.400 ;
        RECT 1.905 596.720 345.600 597.360 ;
        RECT 4.400 596.000 345.600 596.720 ;
        RECT 4.400 595.320 346.000 596.000 ;
        RECT 1.905 594.000 346.000 595.320 ;
        RECT 4.400 592.600 346.000 594.000 ;
        RECT 1.905 591.280 346.000 592.600 ;
        RECT 4.400 589.880 346.000 591.280 ;
        RECT 1.905 589.240 346.000 589.880 ;
        RECT 4.400 587.840 346.000 589.240 ;
        RECT 1.905 587.200 346.000 587.840 ;
        RECT 1.905 586.520 345.600 587.200 ;
        RECT 4.400 585.800 345.600 586.520 ;
        RECT 4.400 585.120 346.000 585.800 ;
        RECT 1.905 583.800 346.000 585.120 ;
        RECT 4.400 582.400 346.000 583.800 ;
        RECT 1.905 581.760 346.000 582.400 ;
        RECT 4.400 580.360 346.000 581.760 ;
        RECT 1.905 579.040 346.000 580.360 ;
        RECT 4.400 577.640 346.000 579.040 ;
        RECT 1.905 577.000 346.000 577.640 ;
        RECT 1.905 576.320 345.600 577.000 ;
        RECT 4.400 575.600 345.600 576.320 ;
        RECT 4.400 574.920 346.000 575.600 ;
        RECT 1.905 574.280 346.000 574.920 ;
        RECT 4.400 572.880 346.000 574.280 ;
        RECT 1.905 571.560 346.000 572.880 ;
        RECT 4.400 570.160 346.000 571.560 ;
        RECT 1.905 568.840 346.000 570.160 ;
        RECT 4.400 567.440 346.000 568.840 ;
        RECT 1.905 566.800 346.000 567.440 ;
        RECT 4.400 565.400 345.600 566.800 ;
        RECT 1.905 564.080 346.000 565.400 ;
        RECT 4.400 562.680 346.000 564.080 ;
        RECT 1.905 561.360 346.000 562.680 ;
        RECT 4.400 559.960 346.000 561.360 ;
        RECT 1.905 559.320 346.000 559.960 ;
        RECT 4.400 557.920 346.000 559.320 ;
        RECT 1.905 556.600 346.000 557.920 ;
        RECT 4.400 555.200 345.600 556.600 ;
        RECT 1.905 553.880 346.000 555.200 ;
        RECT 4.400 552.480 346.000 553.880 ;
        RECT 1.905 551.840 346.000 552.480 ;
        RECT 4.400 550.440 346.000 551.840 ;
        RECT 1.905 549.120 346.000 550.440 ;
        RECT 4.400 547.720 346.000 549.120 ;
        RECT 1.905 546.400 346.000 547.720 ;
        RECT 4.400 545.000 345.600 546.400 ;
        RECT 1.905 544.360 346.000 545.000 ;
        RECT 4.400 542.960 346.000 544.360 ;
        RECT 1.905 541.640 346.000 542.960 ;
        RECT 4.400 540.240 346.000 541.640 ;
        RECT 1.905 538.920 346.000 540.240 ;
        RECT 4.400 537.520 346.000 538.920 ;
        RECT 1.905 536.200 346.000 537.520 ;
        RECT 4.400 534.800 345.600 536.200 ;
        RECT 1.905 534.160 346.000 534.800 ;
        RECT 4.400 532.760 346.000 534.160 ;
        RECT 1.905 531.440 346.000 532.760 ;
        RECT 4.400 530.040 346.000 531.440 ;
        RECT 1.905 528.720 346.000 530.040 ;
        RECT 4.400 527.320 346.000 528.720 ;
        RECT 1.905 526.680 346.000 527.320 ;
        RECT 4.400 526.000 346.000 526.680 ;
        RECT 4.400 525.280 345.600 526.000 ;
        RECT 1.905 524.600 345.600 525.280 ;
        RECT 1.905 523.960 346.000 524.600 ;
        RECT 4.400 522.560 346.000 523.960 ;
        RECT 1.905 521.240 346.000 522.560 ;
        RECT 4.400 519.840 346.000 521.240 ;
        RECT 1.905 519.200 346.000 519.840 ;
        RECT 4.400 517.800 346.000 519.200 ;
        RECT 1.905 516.480 346.000 517.800 ;
        RECT 4.400 515.800 346.000 516.480 ;
        RECT 4.400 515.080 345.600 515.800 ;
        RECT 1.905 514.400 345.600 515.080 ;
        RECT 1.905 513.760 346.000 514.400 ;
        RECT 4.400 512.360 346.000 513.760 ;
        RECT 1.905 511.720 346.000 512.360 ;
        RECT 4.400 510.320 346.000 511.720 ;
        RECT 1.905 509.000 346.000 510.320 ;
        RECT 4.400 507.600 346.000 509.000 ;
        RECT 1.905 506.280 346.000 507.600 ;
        RECT 4.400 505.600 346.000 506.280 ;
        RECT 4.400 504.880 345.600 505.600 ;
        RECT 1.905 504.240 345.600 504.880 ;
        RECT 4.400 504.200 345.600 504.240 ;
        RECT 4.400 502.840 346.000 504.200 ;
        RECT 1.905 501.520 346.000 502.840 ;
        RECT 4.400 500.120 346.000 501.520 ;
        RECT 1.905 498.800 346.000 500.120 ;
        RECT 4.400 497.400 346.000 498.800 ;
        RECT 1.905 496.760 346.000 497.400 ;
        RECT 4.400 495.400 346.000 496.760 ;
        RECT 4.400 495.360 345.600 495.400 ;
        RECT 1.905 494.040 345.600 495.360 ;
        RECT 4.400 494.000 345.600 494.040 ;
        RECT 4.400 492.640 346.000 494.000 ;
        RECT 1.905 491.320 346.000 492.640 ;
        RECT 4.400 489.920 346.000 491.320 ;
        RECT 1.905 489.280 346.000 489.920 ;
        RECT 4.400 487.880 346.000 489.280 ;
        RECT 1.905 486.560 346.000 487.880 ;
        RECT 4.400 485.200 346.000 486.560 ;
        RECT 4.400 485.160 345.600 485.200 ;
        RECT 1.905 483.840 345.600 485.160 ;
        RECT 4.400 483.800 345.600 483.840 ;
        RECT 4.400 482.440 346.000 483.800 ;
        RECT 1.905 481.800 346.000 482.440 ;
        RECT 4.400 480.400 346.000 481.800 ;
        RECT 1.905 479.080 346.000 480.400 ;
        RECT 4.400 477.680 346.000 479.080 ;
        RECT 1.905 476.360 346.000 477.680 ;
        RECT 4.400 475.000 346.000 476.360 ;
        RECT 4.400 474.960 345.600 475.000 ;
        RECT 1.905 474.320 345.600 474.960 ;
        RECT 4.400 473.600 345.600 474.320 ;
        RECT 4.400 472.920 346.000 473.600 ;
        RECT 1.905 471.600 346.000 472.920 ;
        RECT 4.400 470.200 346.000 471.600 ;
        RECT 1.905 468.880 346.000 470.200 ;
        RECT 4.400 467.480 346.000 468.880 ;
        RECT 1.905 466.840 346.000 467.480 ;
        RECT 4.400 465.440 346.000 466.840 ;
        RECT 1.905 464.800 346.000 465.440 ;
        RECT 1.905 464.120 345.600 464.800 ;
        RECT 4.400 463.400 345.600 464.120 ;
        RECT 4.400 462.720 346.000 463.400 ;
        RECT 1.905 461.400 346.000 462.720 ;
        RECT 4.400 460.000 346.000 461.400 ;
        RECT 1.905 458.680 346.000 460.000 ;
        RECT 4.400 457.280 346.000 458.680 ;
        RECT 1.905 456.640 346.000 457.280 ;
        RECT 4.400 455.240 346.000 456.640 ;
        RECT 1.905 454.600 346.000 455.240 ;
        RECT 1.905 453.920 345.600 454.600 ;
        RECT 4.400 453.200 345.600 453.920 ;
        RECT 4.400 452.520 346.000 453.200 ;
        RECT 1.905 451.200 346.000 452.520 ;
        RECT 4.400 449.800 346.000 451.200 ;
        RECT 1.905 449.160 346.000 449.800 ;
        RECT 4.400 447.760 346.000 449.160 ;
        RECT 1.905 446.440 346.000 447.760 ;
        RECT 4.400 445.040 346.000 446.440 ;
        RECT 1.905 444.400 346.000 445.040 ;
        RECT 1.905 443.720 345.600 444.400 ;
        RECT 4.400 443.000 345.600 443.720 ;
        RECT 4.400 442.320 346.000 443.000 ;
        RECT 1.905 441.680 346.000 442.320 ;
        RECT 4.400 440.280 346.000 441.680 ;
        RECT 1.905 438.960 346.000 440.280 ;
        RECT 4.400 437.560 346.000 438.960 ;
        RECT 1.905 436.240 346.000 437.560 ;
        RECT 4.400 434.840 346.000 436.240 ;
        RECT 1.905 434.200 346.000 434.840 ;
        RECT 4.400 432.800 345.600 434.200 ;
        RECT 1.905 431.480 346.000 432.800 ;
        RECT 4.400 430.080 346.000 431.480 ;
        RECT 1.905 428.760 346.000 430.080 ;
        RECT 4.400 427.360 346.000 428.760 ;
        RECT 1.905 426.720 346.000 427.360 ;
        RECT 4.400 425.320 346.000 426.720 ;
        RECT 1.905 424.000 346.000 425.320 ;
        RECT 4.400 422.600 345.600 424.000 ;
        RECT 1.905 421.280 346.000 422.600 ;
        RECT 4.400 419.880 346.000 421.280 ;
        RECT 1.905 419.240 346.000 419.880 ;
        RECT 4.400 417.840 346.000 419.240 ;
        RECT 1.905 416.520 346.000 417.840 ;
        RECT 4.400 415.120 346.000 416.520 ;
        RECT 1.905 413.800 346.000 415.120 ;
        RECT 4.400 412.400 345.600 413.800 ;
        RECT 1.905 411.760 346.000 412.400 ;
        RECT 4.400 410.360 346.000 411.760 ;
        RECT 1.905 409.040 346.000 410.360 ;
        RECT 4.400 407.640 346.000 409.040 ;
        RECT 1.905 406.320 346.000 407.640 ;
        RECT 4.400 404.920 346.000 406.320 ;
        RECT 1.905 404.280 346.000 404.920 ;
        RECT 4.400 403.600 346.000 404.280 ;
        RECT 4.400 402.880 345.600 403.600 ;
        RECT 1.905 402.200 345.600 402.880 ;
        RECT 1.905 401.560 346.000 402.200 ;
        RECT 4.400 400.160 346.000 401.560 ;
        RECT 1.905 398.840 346.000 400.160 ;
        RECT 4.400 397.440 346.000 398.840 ;
        RECT 1.905 396.800 346.000 397.440 ;
        RECT 4.400 395.400 346.000 396.800 ;
        RECT 1.905 394.080 346.000 395.400 ;
        RECT 4.400 393.400 346.000 394.080 ;
        RECT 4.400 392.680 345.600 393.400 ;
        RECT 1.905 392.000 345.600 392.680 ;
        RECT 1.905 391.360 346.000 392.000 ;
        RECT 4.400 389.960 346.000 391.360 ;
        RECT 1.905 389.320 346.000 389.960 ;
        RECT 4.400 387.920 346.000 389.320 ;
        RECT 1.905 386.600 346.000 387.920 ;
        RECT 4.400 385.200 346.000 386.600 ;
        RECT 1.905 383.880 346.000 385.200 ;
        RECT 4.400 383.200 346.000 383.880 ;
        RECT 4.400 382.480 345.600 383.200 ;
        RECT 1.905 381.800 345.600 382.480 ;
        RECT 1.905 381.160 346.000 381.800 ;
        RECT 4.400 379.760 346.000 381.160 ;
        RECT 1.905 379.120 346.000 379.760 ;
        RECT 4.400 377.720 346.000 379.120 ;
        RECT 1.905 376.400 346.000 377.720 ;
        RECT 4.400 375.000 346.000 376.400 ;
        RECT 1.905 373.680 346.000 375.000 ;
        RECT 4.400 373.000 346.000 373.680 ;
        RECT 4.400 372.280 345.600 373.000 ;
        RECT 1.905 371.640 345.600 372.280 ;
        RECT 4.400 371.600 345.600 371.640 ;
        RECT 4.400 370.240 346.000 371.600 ;
        RECT 1.905 368.920 346.000 370.240 ;
        RECT 4.400 367.520 346.000 368.920 ;
        RECT 1.905 366.200 346.000 367.520 ;
        RECT 4.400 364.800 346.000 366.200 ;
        RECT 1.905 364.160 346.000 364.800 ;
        RECT 4.400 362.800 346.000 364.160 ;
        RECT 4.400 362.760 345.600 362.800 ;
        RECT 1.905 361.440 345.600 362.760 ;
        RECT 4.400 361.400 345.600 361.440 ;
        RECT 4.400 360.040 346.000 361.400 ;
        RECT 1.905 358.720 346.000 360.040 ;
        RECT 4.400 357.320 346.000 358.720 ;
        RECT 1.905 356.680 346.000 357.320 ;
        RECT 4.400 355.280 346.000 356.680 ;
        RECT 1.905 353.960 346.000 355.280 ;
        RECT 4.400 352.600 346.000 353.960 ;
        RECT 4.400 352.560 345.600 352.600 ;
        RECT 1.905 351.240 345.600 352.560 ;
        RECT 4.400 351.200 345.600 351.240 ;
        RECT 4.400 349.840 346.000 351.200 ;
        RECT 1.905 349.200 346.000 349.840 ;
        RECT 4.400 347.800 346.000 349.200 ;
        RECT 1.905 346.480 346.000 347.800 ;
        RECT 4.400 345.080 346.000 346.480 ;
        RECT 1.905 343.760 346.000 345.080 ;
        RECT 4.400 342.400 346.000 343.760 ;
        RECT 4.400 342.360 345.600 342.400 ;
        RECT 1.905 341.720 345.600 342.360 ;
        RECT 4.400 341.000 345.600 341.720 ;
        RECT 4.400 340.320 346.000 341.000 ;
        RECT 1.905 339.000 346.000 340.320 ;
        RECT 4.400 337.600 346.000 339.000 ;
        RECT 1.905 336.280 346.000 337.600 ;
        RECT 4.400 334.880 346.000 336.280 ;
        RECT 1.905 334.240 346.000 334.880 ;
        RECT 4.400 332.840 346.000 334.240 ;
        RECT 1.905 332.200 346.000 332.840 ;
        RECT 1.905 331.520 345.600 332.200 ;
        RECT 4.400 330.800 345.600 331.520 ;
        RECT 4.400 330.120 346.000 330.800 ;
        RECT 1.905 328.800 346.000 330.120 ;
        RECT 4.400 327.400 346.000 328.800 ;
        RECT 1.905 326.760 346.000 327.400 ;
        RECT 4.400 325.360 346.000 326.760 ;
        RECT 1.905 324.040 346.000 325.360 ;
        RECT 4.400 322.640 346.000 324.040 ;
        RECT 1.905 322.000 346.000 322.640 ;
        RECT 1.905 321.320 345.600 322.000 ;
        RECT 4.400 320.600 345.600 321.320 ;
        RECT 4.400 319.920 346.000 320.600 ;
        RECT 1.905 319.280 346.000 319.920 ;
        RECT 4.400 317.880 346.000 319.280 ;
        RECT 1.905 316.560 346.000 317.880 ;
        RECT 4.400 315.160 346.000 316.560 ;
        RECT 1.905 313.840 346.000 315.160 ;
        RECT 4.400 312.440 346.000 313.840 ;
        RECT 1.905 311.800 346.000 312.440 ;
        RECT 4.400 310.400 345.600 311.800 ;
        RECT 1.905 309.080 346.000 310.400 ;
        RECT 4.400 307.680 346.000 309.080 ;
        RECT 1.905 306.360 346.000 307.680 ;
        RECT 4.400 304.960 346.000 306.360 ;
        RECT 1.905 303.640 346.000 304.960 ;
        RECT 4.400 302.240 346.000 303.640 ;
        RECT 1.905 301.600 346.000 302.240 ;
        RECT 4.400 300.200 345.600 301.600 ;
        RECT 1.905 298.880 346.000 300.200 ;
        RECT 4.400 297.480 346.000 298.880 ;
        RECT 1.905 296.160 346.000 297.480 ;
        RECT 4.400 294.760 346.000 296.160 ;
        RECT 1.905 294.120 346.000 294.760 ;
        RECT 4.400 292.720 346.000 294.120 ;
        RECT 1.905 291.400 346.000 292.720 ;
        RECT 4.400 290.000 345.600 291.400 ;
        RECT 1.905 288.680 346.000 290.000 ;
        RECT 4.400 287.280 346.000 288.680 ;
        RECT 1.905 286.640 346.000 287.280 ;
        RECT 4.400 285.240 346.000 286.640 ;
        RECT 1.905 283.920 346.000 285.240 ;
        RECT 4.400 282.520 346.000 283.920 ;
        RECT 1.905 281.200 346.000 282.520 ;
        RECT 4.400 279.800 345.600 281.200 ;
        RECT 1.905 279.160 346.000 279.800 ;
        RECT 4.400 277.760 346.000 279.160 ;
        RECT 1.905 276.440 346.000 277.760 ;
        RECT 4.400 275.040 346.000 276.440 ;
        RECT 1.905 273.720 346.000 275.040 ;
        RECT 4.400 272.320 346.000 273.720 ;
        RECT 1.905 271.680 346.000 272.320 ;
        RECT 4.400 271.000 346.000 271.680 ;
        RECT 4.400 270.280 345.600 271.000 ;
        RECT 1.905 269.600 345.600 270.280 ;
        RECT 1.905 268.960 346.000 269.600 ;
        RECT 4.400 267.560 346.000 268.960 ;
        RECT 1.905 266.240 346.000 267.560 ;
        RECT 4.400 264.840 346.000 266.240 ;
        RECT 1.905 264.200 346.000 264.840 ;
        RECT 4.400 262.800 346.000 264.200 ;
        RECT 1.905 261.480 346.000 262.800 ;
        RECT 4.400 260.800 346.000 261.480 ;
        RECT 4.400 260.080 345.600 260.800 ;
        RECT 1.905 259.400 345.600 260.080 ;
        RECT 1.905 258.760 346.000 259.400 ;
        RECT 4.400 257.360 346.000 258.760 ;
        RECT 1.905 256.720 346.000 257.360 ;
        RECT 4.400 255.320 346.000 256.720 ;
        RECT 1.905 254.000 346.000 255.320 ;
        RECT 4.400 252.600 346.000 254.000 ;
        RECT 1.905 251.280 346.000 252.600 ;
        RECT 4.400 250.600 346.000 251.280 ;
        RECT 4.400 249.880 345.600 250.600 ;
        RECT 1.905 249.240 345.600 249.880 ;
        RECT 4.400 249.200 345.600 249.240 ;
        RECT 4.400 247.840 346.000 249.200 ;
        RECT 1.905 246.520 346.000 247.840 ;
        RECT 4.400 245.120 346.000 246.520 ;
        RECT 1.905 243.800 346.000 245.120 ;
        RECT 4.400 242.400 346.000 243.800 ;
        RECT 1.905 241.760 346.000 242.400 ;
        RECT 4.400 240.400 346.000 241.760 ;
        RECT 4.400 240.360 345.600 240.400 ;
        RECT 1.905 239.040 345.600 240.360 ;
        RECT 4.400 239.000 345.600 239.040 ;
        RECT 4.400 237.640 346.000 239.000 ;
        RECT 1.905 236.320 346.000 237.640 ;
        RECT 4.400 234.920 346.000 236.320 ;
        RECT 1.905 234.280 346.000 234.920 ;
        RECT 4.400 232.880 346.000 234.280 ;
        RECT 1.905 231.560 346.000 232.880 ;
        RECT 4.400 230.200 346.000 231.560 ;
        RECT 4.400 230.160 345.600 230.200 ;
        RECT 1.905 228.840 345.600 230.160 ;
        RECT 4.400 228.800 345.600 228.840 ;
        RECT 4.400 227.440 346.000 228.800 ;
        RECT 1.905 226.120 346.000 227.440 ;
        RECT 4.400 224.720 346.000 226.120 ;
        RECT 1.905 224.080 346.000 224.720 ;
        RECT 4.400 222.680 346.000 224.080 ;
        RECT 1.905 221.360 346.000 222.680 ;
        RECT 4.400 220.000 346.000 221.360 ;
        RECT 4.400 219.960 345.600 220.000 ;
        RECT 1.905 218.640 345.600 219.960 ;
        RECT 4.400 218.600 345.600 218.640 ;
        RECT 4.400 217.240 346.000 218.600 ;
        RECT 1.905 216.600 346.000 217.240 ;
        RECT 4.400 215.200 346.000 216.600 ;
        RECT 1.905 213.880 346.000 215.200 ;
        RECT 4.400 212.480 346.000 213.880 ;
        RECT 1.905 211.160 346.000 212.480 ;
        RECT 4.400 209.800 346.000 211.160 ;
        RECT 4.400 209.760 345.600 209.800 ;
        RECT 1.905 209.120 345.600 209.760 ;
        RECT 4.400 208.400 345.600 209.120 ;
        RECT 4.400 207.720 346.000 208.400 ;
        RECT 1.905 206.400 346.000 207.720 ;
        RECT 4.400 205.000 346.000 206.400 ;
        RECT 1.905 203.680 346.000 205.000 ;
        RECT 4.400 202.280 346.000 203.680 ;
        RECT 1.905 201.640 346.000 202.280 ;
        RECT 4.400 200.240 346.000 201.640 ;
        RECT 1.905 199.600 346.000 200.240 ;
        RECT 1.905 198.920 345.600 199.600 ;
        RECT 4.400 198.200 345.600 198.920 ;
        RECT 4.400 197.520 346.000 198.200 ;
        RECT 1.905 196.200 346.000 197.520 ;
        RECT 4.400 194.800 346.000 196.200 ;
        RECT 1.905 194.160 346.000 194.800 ;
        RECT 4.400 192.760 346.000 194.160 ;
        RECT 1.905 191.440 346.000 192.760 ;
        RECT 4.400 190.040 346.000 191.440 ;
        RECT 1.905 189.400 346.000 190.040 ;
        RECT 1.905 188.720 345.600 189.400 ;
        RECT 4.400 188.000 345.600 188.720 ;
        RECT 4.400 187.320 346.000 188.000 ;
        RECT 1.905 186.680 346.000 187.320 ;
        RECT 4.400 185.280 346.000 186.680 ;
        RECT 1.905 183.960 346.000 185.280 ;
        RECT 4.400 182.560 346.000 183.960 ;
        RECT 1.905 181.240 346.000 182.560 ;
        RECT 4.400 179.840 346.000 181.240 ;
        RECT 1.905 179.200 346.000 179.840 ;
        RECT 4.400 177.800 345.600 179.200 ;
        RECT 1.905 176.480 346.000 177.800 ;
        RECT 4.400 175.080 346.000 176.480 ;
        RECT 1.905 173.760 346.000 175.080 ;
        RECT 4.400 172.360 346.000 173.760 ;
        RECT 1.905 171.720 346.000 172.360 ;
        RECT 4.400 170.320 346.000 171.720 ;
        RECT 1.905 169.000 346.000 170.320 ;
        RECT 4.400 167.600 345.600 169.000 ;
        RECT 1.905 166.280 346.000 167.600 ;
        RECT 4.400 164.880 346.000 166.280 ;
        RECT 1.905 164.240 346.000 164.880 ;
        RECT 4.400 162.840 346.000 164.240 ;
        RECT 1.905 161.520 346.000 162.840 ;
        RECT 4.400 160.120 346.000 161.520 ;
        RECT 1.905 158.800 346.000 160.120 ;
        RECT 4.400 157.400 345.600 158.800 ;
        RECT 1.905 156.760 346.000 157.400 ;
        RECT 4.400 155.360 346.000 156.760 ;
        RECT 1.905 154.040 346.000 155.360 ;
        RECT 4.400 152.640 346.000 154.040 ;
        RECT 1.905 151.320 346.000 152.640 ;
        RECT 4.400 149.920 346.000 151.320 ;
        RECT 1.905 148.600 346.000 149.920 ;
        RECT 4.400 147.200 345.600 148.600 ;
        RECT 1.905 146.560 346.000 147.200 ;
        RECT 4.400 145.160 346.000 146.560 ;
        RECT 1.905 143.840 346.000 145.160 ;
        RECT 4.400 142.440 346.000 143.840 ;
        RECT 1.905 141.120 346.000 142.440 ;
        RECT 4.400 139.720 346.000 141.120 ;
        RECT 1.905 139.080 346.000 139.720 ;
        RECT 4.400 138.400 346.000 139.080 ;
        RECT 4.400 137.680 345.600 138.400 ;
        RECT 1.905 137.000 345.600 137.680 ;
        RECT 1.905 136.360 346.000 137.000 ;
        RECT 4.400 134.960 346.000 136.360 ;
        RECT 1.905 133.640 346.000 134.960 ;
        RECT 4.400 132.240 346.000 133.640 ;
        RECT 1.905 131.600 346.000 132.240 ;
        RECT 4.400 130.200 346.000 131.600 ;
        RECT 1.905 128.880 346.000 130.200 ;
        RECT 4.400 128.200 346.000 128.880 ;
        RECT 4.400 127.480 345.600 128.200 ;
        RECT 1.905 126.800 345.600 127.480 ;
        RECT 1.905 126.160 346.000 126.800 ;
        RECT 4.400 124.760 346.000 126.160 ;
        RECT 1.905 124.120 346.000 124.760 ;
        RECT 4.400 122.720 346.000 124.120 ;
        RECT 1.905 121.400 346.000 122.720 ;
        RECT 4.400 120.000 346.000 121.400 ;
        RECT 1.905 118.680 346.000 120.000 ;
        RECT 4.400 118.000 346.000 118.680 ;
        RECT 4.400 117.280 345.600 118.000 ;
        RECT 1.905 116.640 345.600 117.280 ;
        RECT 4.400 116.600 345.600 116.640 ;
        RECT 4.400 115.240 346.000 116.600 ;
        RECT 1.905 113.920 346.000 115.240 ;
        RECT 4.400 112.520 346.000 113.920 ;
        RECT 1.905 111.200 346.000 112.520 ;
        RECT 4.400 109.800 346.000 111.200 ;
        RECT 1.905 109.160 346.000 109.800 ;
        RECT 4.400 107.800 346.000 109.160 ;
        RECT 4.400 107.760 345.600 107.800 ;
        RECT 1.905 106.440 345.600 107.760 ;
        RECT 4.400 106.400 345.600 106.440 ;
        RECT 4.400 105.040 346.000 106.400 ;
        RECT 1.905 103.720 346.000 105.040 ;
        RECT 4.400 102.320 346.000 103.720 ;
        RECT 1.905 101.680 346.000 102.320 ;
        RECT 4.400 100.280 346.000 101.680 ;
        RECT 1.905 98.960 346.000 100.280 ;
        RECT 4.400 97.600 346.000 98.960 ;
        RECT 4.400 97.560 345.600 97.600 ;
        RECT 1.905 96.240 345.600 97.560 ;
        RECT 4.400 96.200 345.600 96.240 ;
        RECT 4.400 94.840 346.000 96.200 ;
        RECT 1.905 94.200 346.000 94.840 ;
        RECT 4.400 92.800 346.000 94.200 ;
        RECT 1.905 91.480 346.000 92.800 ;
        RECT 4.400 90.080 346.000 91.480 ;
        RECT 1.905 88.760 346.000 90.080 ;
        RECT 4.400 87.400 346.000 88.760 ;
        RECT 4.400 87.360 345.600 87.400 ;
        RECT 1.905 86.720 345.600 87.360 ;
        RECT 4.400 86.000 345.600 86.720 ;
        RECT 4.400 85.320 346.000 86.000 ;
        RECT 1.905 84.000 346.000 85.320 ;
        RECT 4.400 82.600 346.000 84.000 ;
        RECT 1.905 81.280 346.000 82.600 ;
        RECT 4.400 79.880 346.000 81.280 ;
        RECT 1.905 79.240 346.000 79.880 ;
        RECT 4.400 77.840 346.000 79.240 ;
        RECT 1.905 77.200 346.000 77.840 ;
        RECT 1.905 76.520 345.600 77.200 ;
        RECT 4.400 75.800 345.600 76.520 ;
        RECT 4.400 75.120 346.000 75.800 ;
        RECT 1.905 73.800 346.000 75.120 ;
        RECT 4.400 72.400 346.000 73.800 ;
        RECT 1.905 71.080 346.000 72.400 ;
        RECT 4.400 69.680 346.000 71.080 ;
        RECT 1.905 69.040 346.000 69.680 ;
        RECT 4.400 67.640 346.000 69.040 ;
        RECT 1.905 67.000 346.000 67.640 ;
        RECT 1.905 66.320 345.600 67.000 ;
        RECT 4.400 65.600 345.600 66.320 ;
        RECT 4.400 64.920 346.000 65.600 ;
        RECT 1.905 63.600 346.000 64.920 ;
        RECT 4.400 62.200 346.000 63.600 ;
        RECT 1.905 61.560 346.000 62.200 ;
        RECT 4.400 60.160 346.000 61.560 ;
        RECT 1.905 58.840 346.000 60.160 ;
        RECT 4.400 57.440 346.000 58.840 ;
        RECT 1.905 56.800 346.000 57.440 ;
        RECT 1.905 56.120 345.600 56.800 ;
        RECT 4.400 55.400 345.600 56.120 ;
        RECT 4.400 54.720 346.000 55.400 ;
        RECT 1.905 54.080 346.000 54.720 ;
        RECT 4.400 52.680 346.000 54.080 ;
        RECT 1.905 51.360 346.000 52.680 ;
        RECT 4.400 49.960 346.000 51.360 ;
        RECT 1.905 48.640 346.000 49.960 ;
        RECT 4.400 47.240 346.000 48.640 ;
        RECT 1.905 46.600 346.000 47.240 ;
        RECT 4.400 45.200 345.600 46.600 ;
        RECT 1.905 43.880 346.000 45.200 ;
        RECT 4.400 42.480 346.000 43.880 ;
        RECT 1.905 41.160 346.000 42.480 ;
        RECT 4.400 39.760 346.000 41.160 ;
        RECT 1.905 39.120 346.000 39.760 ;
        RECT 4.400 37.720 346.000 39.120 ;
        RECT 1.905 36.400 346.000 37.720 ;
        RECT 4.400 35.000 345.600 36.400 ;
        RECT 1.905 33.680 346.000 35.000 ;
        RECT 4.400 32.280 346.000 33.680 ;
        RECT 1.905 31.640 346.000 32.280 ;
        RECT 4.400 30.240 346.000 31.640 ;
        RECT 1.905 28.920 346.000 30.240 ;
        RECT 4.400 27.520 346.000 28.920 ;
        RECT 1.905 26.200 346.000 27.520 ;
        RECT 4.400 24.800 345.600 26.200 ;
        RECT 1.905 24.160 346.000 24.800 ;
        RECT 4.400 22.760 346.000 24.160 ;
        RECT 1.905 21.440 346.000 22.760 ;
        RECT 4.400 20.040 346.000 21.440 ;
        RECT 1.905 18.720 346.000 20.040 ;
        RECT 4.400 17.320 346.000 18.720 ;
        RECT 1.905 16.680 346.000 17.320 ;
        RECT 4.400 16.000 346.000 16.680 ;
        RECT 4.400 15.280 345.600 16.000 ;
        RECT 1.905 14.600 345.600 15.280 ;
        RECT 1.905 13.960 346.000 14.600 ;
        RECT 4.400 12.560 346.000 13.960 ;
        RECT 1.905 11.240 346.000 12.560 ;
        RECT 4.400 9.840 346.000 11.240 ;
        RECT 1.905 9.200 346.000 9.840 ;
        RECT 4.400 7.800 346.000 9.200 ;
        RECT 1.905 6.480 346.000 7.800 ;
        RECT 4.400 5.800 346.000 6.480 ;
        RECT 4.400 5.080 345.600 5.800 ;
        RECT 1.905 4.400 345.600 5.080 ;
        RECT 1.905 3.760 346.000 4.400 ;
        RECT 4.400 2.360 346.000 3.760 ;
        RECT 1.905 1.720 346.000 2.360 ;
        RECT 4.400 0.855 346.000 1.720 ;
      LAYER met4 ;
        RECT 3.070 18.535 20.640 985.825 ;
        RECT 23.040 18.535 97.440 985.825 ;
        RECT 99.840 18.535 174.240 985.825 ;
        RECT 176.640 18.535 226.945 985.825 ;
  END
END WishboneInterconnect
END LIBRARY

