magic
tech sky130A
magscale 1 2
timestamp 1685098217
<< obsli1 >>
rect 1104 2159 98808 157777
<< obsm1 >>
rect 14 892 99990 158704
<< metal2 >>
rect 2778 159200 2834 160000
rect 5262 159200 5318 160000
rect 7746 159200 7802 160000
rect 10230 159200 10286 160000
rect 12714 159200 12770 160000
rect 15198 159200 15254 160000
rect 17682 159200 17738 160000
rect 20166 159200 20222 160000
rect 22650 159200 22706 160000
rect 25134 159200 25190 160000
rect 27618 159200 27674 160000
rect 30102 159200 30158 160000
rect 32586 159200 32642 160000
rect 35070 159200 35126 160000
rect 37554 159200 37610 160000
rect 40038 159200 40094 160000
rect 42522 159200 42578 160000
rect 45006 159200 45062 160000
rect 47490 159200 47546 160000
rect 49974 159200 50030 160000
rect 52458 159200 52514 160000
rect 54942 159200 54998 160000
rect 57426 159200 57482 160000
rect 59910 159200 59966 160000
rect 62394 159200 62450 160000
rect 64878 159200 64934 160000
rect 67362 159200 67418 160000
rect 69846 159200 69902 160000
rect 72330 159200 72386 160000
rect 74814 159200 74870 160000
rect 77298 159200 77354 160000
rect 79782 159200 79838 160000
rect 82266 159200 82322 160000
rect 84750 159200 84806 160000
rect 87234 159200 87290 160000
rect 89718 159200 89774 160000
rect 92202 159200 92258 160000
rect 94686 159200 94742 160000
rect 97170 159200 97226 160000
rect 1858 0 1914 800
rect 3606 0 3662 800
rect 5354 0 5410 800
rect 7102 0 7158 800
rect 8850 0 8906 800
rect 10598 0 10654 800
rect 12346 0 12402 800
rect 14094 0 14150 800
rect 15842 0 15898 800
rect 17590 0 17646 800
rect 19338 0 19394 800
rect 21086 0 21142 800
rect 22834 0 22890 800
rect 24582 0 24638 800
rect 26330 0 26386 800
rect 28078 0 28134 800
rect 29826 0 29882 800
rect 31574 0 31630 800
rect 33322 0 33378 800
rect 35070 0 35126 800
rect 36818 0 36874 800
rect 38566 0 38622 800
rect 40314 0 40370 800
rect 42062 0 42118 800
rect 43810 0 43866 800
rect 45558 0 45614 800
rect 47306 0 47362 800
rect 49054 0 49110 800
rect 50802 0 50858 800
rect 52550 0 52606 800
rect 54298 0 54354 800
rect 56046 0 56102 800
rect 57794 0 57850 800
rect 59542 0 59598 800
rect 61290 0 61346 800
rect 63038 0 63094 800
rect 64786 0 64842 800
rect 66534 0 66590 800
rect 68282 0 68338 800
rect 70030 0 70086 800
rect 71778 0 71834 800
rect 73526 0 73582 800
rect 75274 0 75330 800
rect 77022 0 77078 800
rect 78770 0 78826 800
rect 80518 0 80574 800
rect 82266 0 82322 800
rect 84014 0 84070 800
rect 85762 0 85818 800
rect 87510 0 87566 800
rect 89258 0 89314 800
rect 91006 0 91062 800
rect 92754 0 92810 800
rect 94502 0 94558 800
rect 96250 0 96306 800
rect 97998 0 98054 800
<< obsm2 >>
rect 18 159144 2722 159338
rect 2890 159144 5206 159338
rect 5374 159144 7690 159338
rect 7858 159144 10174 159338
rect 10342 159144 12658 159338
rect 12826 159144 15142 159338
rect 15310 159144 17626 159338
rect 17794 159144 20110 159338
rect 20278 159144 22594 159338
rect 22762 159144 25078 159338
rect 25246 159144 27562 159338
rect 27730 159144 30046 159338
rect 30214 159144 32530 159338
rect 32698 159144 35014 159338
rect 35182 159144 37498 159338
rect 37666 159144 39982 159338
rect 40150 159144 42466 159338
rect 42634 159144 44950 159338
rect 45118 159144 47434 159338
rect 47602 159144 49918 159338
rect 50086 159144 52402 159338
rect 52570 159144 54886 159338
rect 55054 159144 57370 159338
rect 57538 159144 59854 159338
rect 60022 159144 62338 159338
rect 62506 159144 64822 159338
rect 64990 159144 67306 159338
rect 67474 159144 69790 159338
rect 69958 159144 72274 159338
rect 72442 159144 74758 159338
rect 74926 159144 77242 159338
rect 77410 159144 79726 159338
rect 79894 159144 82210 159338
rect 82378 159144 84694 159338
rect 84862 159144 87178 159338
rect 87346 159144 89662 159338
rect 89830 159144 92146 159338
rect 92314 159144 94630 159338
rect 94798 159144 97114 159338
rect 97282 159144 99986 159338
rect 18 856 99986 159144
rect 18 734 1802 856
rect 1970 734 3550 856
rect 3718 734 5298 856
rect 5466 734 7046 856
rect 7214 734 8794 856
rect 8962 734 10542 856
rect 10710 734 12290 856
rect 12458 734 14038 856
rect 14206 734 15786 856
rect 15954 734 17534 856
rect 17702 734 19282 856
rect 19450 734 21030 856
rect 21198 734 22778 856
rect 22946 734 24526 856
rect 24694 734 26274 856
rect 26442 734 28022 856
rect 28190 734 29770 856
rect 29938 734 31518 856
rect 31686 734 33266 856
rect 33434 734 35014 856
rect 35182 734 36762 856
rect 36930 734 38510 856
rect 38678 734 40258 856
rect 40426 734 42006 856
rect 42174 734 43754 856
rect 43922 734 45502 856
rect 45670 734 47250 856
rect 47418 734 48998 856
rect 49166 734 50746 856
rect 50914 734 52494 856
rect 52662 734 54242 856
rect 54410 734 55990 856
rect 56158 734 57738 856
rect 57906 734 59486 856
rect 59654 734 61234 856
rect 61402 734 62982 856
rect 63150 734 64730 856
rect 64898 734 66478 856
rect 66646 734 68226 856
rect 68394 734 69974 856
rect 70142 734 71722 856
rect 71890 734 73470 856
rect 73638 734 75218 856
rect 75386 734 76966 856
rect 77134 734 78714 856
rect 78882 734 80462 856
rect 80630 734 82210 856
rect 82378 734 83958 856
rect 84126 734 85706 856
rect 85874 734 87454 856
rect 87622 734 89202 856
rect 89370 734 90950 856
rect 91118 734 92698 856
rect 92866 734 94446 856
rect 94614 734 96194 856
rect 96362 734 97942 856
rect 98110 734 99986 856
<< metal3 >>
rect 0 158176 800 158296
rect 0 157360 800 157480
rect 0 156544 800 156664
rect 0 155728 800 155848
rect 0 154912 800 155032
rect 0 154096 800 154216
rect 0 153280 800 153400
rect 0 152464 800 152584
rect 0 151648 800 151768
rect 0 150832 800 150952
rect 0 150016 800 150136
rect 0 149200 800 149320
rect 0 148384 800 148504
rect 99200 148248 100000 148368
rect 0 147568 800 147688
rect 99200 147568 100000 147688
rect 0 146752 800 146872
rect 99200 146888 100000 147008
rect 99200 146208 100000 146328
rect 0 145936 800 146056
rect 99200 145528 100000 145648
rect 0 145120 800 145240
rect 99200 144848 100000 144968
rect 0 144304 800 144424
rect 99200 144168 100000 144288
rect 0 143488 800 143608
rect 99200 143488 100000 143608
rect 0 142672 800 142792
rect 99200 142808 100000 142928
rect 99200 142128 100000 142248
rect 0 141856 800 141976
rect 99200 141448 100000 141568
rect 0 141040 800 141160
rect 99200 140768 100000 140888
rect 0 140224 800 140344
rect 99200 140088 100000 140208
rect 0 139408 800 139528
rect 99200 139408 100000 139528
rect 0 138592 800 138712
rect 99200 138728 100000 138848
rect 99200 138048 100000 138168
rect 0 137776 800 137896
rect 99200 137368 100000 137488
rect 0 136960 800 137080
rect 99200 136688 100000 136808
rect 0 136144 800 136264
rect 99200 136008 100000 136128
rect 0 135328 800 135448
rect 99200 135328 100000 135448
rect 0 134512 800 134632
rect 99200 134648 100000 134768
rect 99200 133968 100000 134088
rect 0 133696 800 133816
rect 99200 133288 100000 133408
rect 0 132880 800 133000
rect 99200 132608 100000 132728
rect 0 132064 800 132184
rect 99200 131928 100000 132048
rect 0 131248 800 131368
rect 99200 131248 100000 131368
rect 0 130432 800 130552
rect 99200 130568 100000 130688
rect 99200 129888 100000 130008
rect 0 129616 800 129736
rect 99200 129208 100000 129328
rect 0 128800 800 128920
rect 99200 128528 100000 128648
rect 0 127984 800 128104
rect 99200 127848 100000 127968
rect 0 127168 800 127288
rect 99200 127168 100000 127288
rect 0 126352 800 126472
rect 99200 126488 100000 126608
rect 99200 125808 100000 125928
rect 0 125536 800 125656
rect 99200 125128 100000 125248
rect 0 124720 800 124840
rect 99200 124448 100000 124568
rect 0 123904 800 124024
rect 99200 123768 100000 123888
rect 0 123088 800 123208
rect 99200 123088 100000 123208
rect 0 122272 800 122392
rect 99200 122408 100000 122528
rect 99200 121728 100000 121848
rect 0 121456 800 121576
rect 99200 121048 100000 121168
rect 0 120640 800 120760
rect 99200 120368 100000 120488
rect 0 119824 800 119944
rect 99200 119688 100000 119808
rect 0 119008 800 119128
rect 99200 119008 100000 119128
rect 0 118192 800 118312
rect 99200 118328 100000 118448
rect 99200 117648 100000 117768
rect 0 117376 800 117496
rect 99200 116968 100000 117088
rect 0 116560 800 116680
rect 99200 116288 100000 116408
rect 0 115744 800 115864
rect 99200 115608 100000 115728
rect 0 114928 800 115048
rect 99200 114928 100000 115048
rect 0 114112 800 114232
rect 99200 114248 100000 114368
rect 99200 113568 100000 113688
rect 0 113296 800 113416
rect 99200 112888 100000 113008
rect 0 112480 800 112600
rect 99200 112208 100000 112328
rect 0 111664 800 111784
rect 99200 111528 100000 111648
rect 0 110848 800 110968
rect 99200 110848 100000 110968
rect 0 110032 800 110152
rect 99200 110168 100000 110288
rect 99200 109488 100000 109608
rect 0 109216 800 109336
rect 99200 108808 100000 108928
rect 0 108400 800 108520
rect 99200 108128 100000 108248
rect 0 107584 800 107704
rect 99200 107448 100000 107568
rect 0 106768 800 106888
rect 99200 106768 100000 106888
rect 0 105952 800 106072
rect 99200 106088 100000 106208
rect 99200 105408 100000 105528
rect 0 105136 800 105256
rect 99200 104728 100000 104848
rect 0 104320 800 104440
rect 99200 104048 100000 104168
rect 0 103504 800 103624
rect 99200 103368 100000 103488
rect 0 102688 800 102808
rect 99200 102688 100000 102808
rect 0 101872 800 101992
rect 99200 102008 100000 102128
rect 99200 101328 100000 101448
rect 0 101056 800 101176
rect 99200 100648 100000 100768
rect 0 100240 800 100360
rect 99200 99968 100000 100088
rect 0 99424 800 99544
rect 99200 99288 100000 99408
rect 0 98608 800 98728
rect 99200 98608 100000 98728
rect 0 97792 800 97912
rect 99200 97928 100000 98048
rect 99200 97248 100000 97368
rect 0 96976 800 97096
rect 99200 96568 100000 96688
rect 0 96160 800 96280
rect 99200 95888 100000 96008
rect 0 95344 800 95464
rect 99200 95208 100000 95328
rect 0 94528 800 94648
rect 99200 94528 100000 94648
rect 0 93712 800 93832
rect 99200 93848 100000 93968
rect 99200 93168 100000 93288
rect 0 92896 800 93016
rect 99200 92488 100000 92608
rect 0 92080 800 92200
rect 99200 91808 100000 91928
rect 0 91264 800 91384
rect 99200 91128 100000 91248
rect 0 90448 800 90568
rect 99200 90448 100000 90568
rect 0 89632 800 89752
rect 99200 89768 100000 89888
rect 99200 89088 100000 89208
rect 0 88816 800 88936
rect 99200 88408 100000 88528
rect 0 88000 800 88120
rect 99200 87728 100000 87848
rect 0 87184 800 87304
rect 99200 87048 100000 87168
rect 0 86368 800 86488
rect 99200 86368 100000 86488
rect 0 85552 800 85672
rect 99200 85688 100000 85808
rect 99200 85008 100000 85128
rect 0 84736 800 84856
rect 99200 84328 100000 84448
rect 0 83920 800 84040
rect 99200 83648 100000 83768
rect 0 83104 800 83224
rect 99200 82968 100000 83088
rect 0 82288 800 82408
rect 99200 82288 100000 82408
rect 0 81472 800 81592
rect 99200 81608 100000 81728
rect 99200 80928 100000 81048
rect 0 80656 800 80776
rect 99200 80248 100000 80368
rect 0 79840 800 79960
rect 99200 79568 100000 79688
rect 0 79024 800 79144
rect 99200 78888 100000 79008
rect 0 78208 800 78328
rect 99200 78208 100000 78328
rect 0 77392 800 77512
rect 99200 77528 100000 77648
rect 99200 76848 100000 76968
rect 0 76576 800 76696
rect 99200 76168 100000 76288
rect 0 75760 800 75880
rect 99200 75488 100000 75608
rect 0 74944 800 75064
rect 99200 74808 100000 74928
rect 0 74128 800 74248
rect 99200 74128 100000 74248
rect 0 73312 800 73432
rect 99200 73448 100000 73568
rect 99200 72768 100000 72888
rect 0 72496 800 72616
rect 99200 72088 100000 72208
rect 0 71680 800 71800
rect 99200 71408 100000 71528
rect 0 70864 800 70984
rect 99200 70728 100000 70848
rect 0 70048 800 70168
rect 99200 70048 100000 70168
rect 0 69232 800 69352
rect 99200 69368 100000 69488
rect 99200 68688 100000 68808
rect 0 68416 800 68536
rect 99200 68008 100000 68128
rect 0 67600 800 67720
rect 99200 67328 100000 67448
rect 0 66784 800 66904
rect 99200 66648 100000 66768
rect 0 65968 800 66088
rect 99200 65968 100000 66088
rect 0 65152 800 65272
rect 99200 65288 100000 65408
rect 99200 64608 100000 64728
rect 0 64336 800 64456
rect 99200 63928 100000 64048
rect 0 63520 800 63640
rect 99200 63248 100000 63368
rect 0 62704 800 62824
rect 99200 62568 100000 62688
rect 0 61888 800 62008
rect 99200 61888 100000 62008
rect 0 61072 800 61192
rect 99200 61208 100000 61328
rect 99200 60528 100000 60648
rect 0 60256 800 60376
rect 99200 59848 100000 59968
rect 0 59440 800 59560
rect 99200 59168 100000 59288
rect 0 58624 800 58744
rect 99200 58488 100000 58608
rect 0 57808 800 57928
rect 99200 57808 100000 57928
rect 0 56992 800 57112
rect 99200 57128 100000 57248
rect 99200 56448 100000 56568
rect 0 56176 800 56296
rect 99200 55768 100000 55888
rect 0 55360 800 55480
rect 99200 55088 100000 55208
rect 0 54544 800 54664
rect 99200 54408 100000 54528
rect 0 53728 800 53848
rect 99200 53728 100000 53848
rect 0 52912 800 53032
rect 99200 53048 100000 53168
rect 99200 52368 100000 52488
rect 0 52096 800 52216
rect 99200 51688 100000 51808
rect 0 51280 800 51400
rect 99200 51008 100000 51128
rect 0 50464 800 50584
rect 99200 50328 100000 50448
rect 0 49648 800 49768
rect 99200 49648 100000 49768
rect 0 48832 800 48952
rect 99200 48968 100000 49088
rect 99200 48288 100000 48408
rect 0 48016 800 48136
rect 99200 47608 100000 47728
rect 0 47200 800 47320
rect 99200 46928 100000 47048
rect 0 46384 800 46504
rect 99200 46248 100000 46368
rect 0 45568 800 45688
rect 99200 45568 100000 45688
rect 0 44752 800 44872
rect 99200 44888 100000 45008
rect 99200 44208 100000 44328
rect 0 43936 800 44056
rect 99200 43528 100000 43648
rect 0 43120 800 43240
rect 99200 42848 100000 42968
rect 0 42304 800 42424
rect 99200 42168 100000 42288
rect 0 41488 800 41608
rect 99200 41488 100000 41608
rect 0 40672 800 40792
rect 99200 40808 100000 40928
rect 99200 40128 100000 40248
rect 0 39856 800 39976
rect 99200 39448 100000 39568
rect 0 39040 800 39160
rect 99200 38768 100000 38888
rect 0 38224 800 38344
rect 99200 38088 100000 38208
rect 0 37408 800 37528
rect 99200 37408 100000 37528
rect 0 36592 800 36712
rect 99200 36728 100000 36848
rect 99200 36048 100000 36168
rect 0 35776 800 35896
rect 99200 35368 100000 35488
rect 0 34960 800 35080
rect 99200 34688 100000 34808
rect 0 34144 800 34264
rect 99200 34008 100000 34128
rect 0 33328 800 33448
rect 99200 33328 100000 33448
rect 0 32512 800 32632
rect 99200 32648 100000 32768
rect 99200 31968 100000 32088
rect 0 31696 800 31816
rect 99200 31288 100000 31408
rect 0 30880 800 31000
rect 99200 30608 100000 30728
rect 0 30064 800 30184
rect 99200 29928 100000 30048
rect 0 29248 800 29368
rect 99200 29248 100000 29368
rect 0 28432 800 28552
rect 99200 28568 100000 28688
rect 99200 27888 100000 28008
rect 0 27616 800 27736
rect 99200 27208 100000 27328
rect 0 26800 800 26920
rect 99200 26528 100000 26648
rect 0 25984 800 26104
rect 99200 25848 100000 25968
rect 0 25168 800 25288
rect 99200 25168 100000 25288
rect 0 24352 800 24472
rect 99200 24488 100000 24608
rect 99200 23808 100000 23928
rect 0 23536 800 23656
rect 99200 23128 100000 23248
rect 0 22720 800 22840
rect 99200 22448 100000 22568
rect 0 21904 800 22024
rect 99200 21768 100000 21888
rect 0 21088 800 21208
rect 99200 21088 100000 21208
rect 0 20272 800 20392
rect 99200 20408 100000 20528
rect 99200 19728 100000 19848
rect 0 19456 800 19576
rect 99200 19048 100000 19168
rect 0 18640 800 18760
rect 99200 18368 100000 18488
rect 0 17824 800 17944
rect 99200 17688 100000 17808
rect 0 17008 800 17128
rect 99200 17008 100000 17128
rect 0 16192 800 16312
rect 99200 16328 100000 16448
rect 99200 15648 100000 15768
rect 0 15376 800 15496
rect 99200 14968 100000 15088
rect 0 14560 800 14680
rect 99200 14288 100000 14408
rect 0 13744 800 13864
rect 99200 13608 100000 13728
rect 0 12928 800 13048
rect 99200 12928 100000 13048
rect 0 12112 800 12232
rect 99200 12248 100000 12368
rect 99200 11568 100000 11688
rect 0 11296 800 11416
rect 0 10480 800 10600
rect 0 9664 800 9784
rect 0 8848 800 8968
rect 0 8032 800 8152
rect 0 7216 800 7336
rect 0 6400 800 6520
rect 0 5584 800 5704
rect 0 4768 800 4888
rect 0 3952 800 4072
rect 0 3136 800 3256
rect 0 2320 800 2440
rect 0 1504 800 1624
<< obsm3 >>
rect 880 158096 99991 158269
rect 13 157560 99991 158096
rect 880 157280 99991 157560
rect 13 156744 99991 157280
rect 880 156464 99991 156744
rect 13 155928 99991 156464
rect 880 155648 99991 155928
rect 13 155112 99991 155648
rect 880 154832 99991 155112
rect 13 154296 99991 154832
rect 880 154016 99991 154296
rect 13 153480 99991 154016
rect 880 153200 99991 153480
rect 13 152664 99991 153200
rect 880 152384 99991 152664
rect 13 151848 99991 152384
rect 880 151568 99991 151848
rect 13 151032 99991 151568
rect 880 150752 99991 151032
rect 13 150216 99991 150752
rect 880 149936 99991 150216
rect 13 149400 99991 149936
rect 880 149120 99991 149400
rect 13 148584 99991 149120
rect 880 148448 99991 148584
rect 880 148304 99120 148448
rect 13 148168 99120 148304
rect 13 147768 99991 148168
rect 880 147488 99120 147768
rect 13 147088 99991 147488
rect 13 146952 99120 147088
rect 880 146808 99120 146952
rect 880 146672 99991 146808
rect 13 146408 99991 146672
rect 13 146136 99120 146408
rect 880 146128 99120 146136
rect 880 145856 99991 146128
rect 13 145728 99991 145856
rect 13 145448 99120 145728
rect 13 145320 99991 145448
rect 880 145048 99991 145320
rect 880 145040 99120 145048
rect 13 144768 99120 145040
rect 13 144504 99991 144768
rect 880 144368 99991 144504
rect 880 144224 99120 144368
rect 13 144088 99120 144224
rect 13 143688 99991 144088
rect 880 143408 99120 143688
rect 13 143008 99991 143408
rect 13 142872 99120 143008
rect 880 142728 99120 142872
rect 880 142592 99991 142728
rect 13 142328 99991 142592
rect 13 142056 99120 142328
rect 880 142048 99120 142056
rect 880 141776 99991 142048
rect 13 141648 99991 141776
rect 13 141368 99120 141648
rect 13 141240 99991 141368
rect 880 140968 99991 141240
rect 880 140960 99120 140968
rect 13 140688 99120 140960
rect 13 140424 99991 140688
rect 880 140288 99991 140424
rect 880 140144 99120 140288
rect 13 140008 99120 140144
rect 13 139608 99991 140008
rect 880 139328 99120 139608
rect 13 138928 99991 139328
rect 13 138792 99120 138928
rect 880 138648 99120 138792
rect 880 138512 99991 138648
rect 13 138248 99991 138512
rect 13 137976 99120 138248
rect 880 137968 99120 137976
rect 880 137696 99991 137968
rect 13 137568 99991 137696
rect 13 137288 99120 137568
rect 13 137160 99991 137288
rect 880 136888 99991 137160
rect 880 136880 99120 136888
rect 13 136608 99120 136880
rect 13 136344 99991 136608
rect 880 136208 99991 136344
rect 880 136064 99120 136208
rect 13 135928 99120 136064
rect 13 135528 99991 135928
rect 880 135248 99120 135528
rect 13 134848 99991 135248
rect 13 134712 99120 134848
rect 880 134568 99120 134712
rect 880 134432 99991 134568
rect 13 134168 99991 134432
rect 13 133896 99120 134168
rect 880 133888 99120 133896
rect 880 133616 99991 133888
rect 13 133488 99991 133616
rect 13 133208 99120 133488
rect 13 133080 99991 133208
rect 880 132808 99991 133080
rect 880 132800 99120 132808
rect 13 132528 99120 132800
rect 13 132264 99991 132528
rect 880 132128 99991 132264
rect 880 131984 99120 132128
rect 13 131848 99120 131984
rect 13 131448 99991 131848
rect 880 131168 99120 131448
rect 13 130768 99991 131168
rect 13 130632 99120 130768
rect 880 130488 99120 130632
rect 880 130352 99991 130488
rect 13 130088 99991 130352
rect 13 129816 99120 130088
rect 880 129808 99120 129816
rect 880 129536 99991 129808
rect 13 129408 99991 129536
rect 13 129128 99120 129408
rect 13 129000 99991 129128
rect 880 128728 99991 129000
rect 880 128720 99120 128728
rect 13 128448 99120 128720
rect 13 128184 99991 128448
rect 880 128048 99991 128184
rect 880 127904 99120 128048
rect 13 127768 99120 127904
rect 13 127368 99991 127768
rect 880 127088 99120 127368
rect 13 126688 99991 127088
rect 13 126552 99120 126688
rect 880 126408 99120 126552
rect 880 126272 99991 126408
rect 13 126008 99991 126272
rect 13 125736 99120 126008
rect 880 125728 99120 125736
rect 880 125456 99991 125728
rect 13 125328 99991 125456
rect 13 125048 99120 125328
rect 13 124920 99991 125048
rect 880 124648 99991 124920
rect 880 124640 99120 124648
rect 13 124368 99120 124640
rect 13 124104 99991 124368
rect 880 123968 99991 124104
rect 880 123824 99120 123968
rect 13 123688 99120 123824
rect 13 123288 99991 123688
rect 880 123008 99120 123288
rect 13 122608 99991 123008
rect 13 122472 99120 122608
rect 880 122328 99120 122472
rect 880 122192 99991 122328
rect 13 121928 99991 122192
rect 13 121656 99120 121928
rect 880 121648 99120 121656
rect 880 121376 99991 121648
rect 13 121248 99991 121376
rect 13 120968 99120 121248
rect 13 120840 99991 120968
rect 880 120568 99991 120840
rect 880 120560 99120 120568
rect 13 120288 99120 120560
rect 13 120024 99991 120288
rect 880 119888 99991 120024
rect 880 119744 99120 119888
rect 13 119608 99120 119744
rect 13 119208 99991 119608
rect 880 118928 99120 119208
rect 13 118528 99991 118928
rect 13 118392 99120 118528
rect 880 118248 99120 118392
rect 880 118112 99991 118248
rect 13 117848 99991 118112
rect 13 117576 99120 117848
rect 880 117568 99120 117576
rect 880 117296 99991 117568
rect 13 117168 99991 117296
rect 13 116888 99120 117168
rect 13 116760 99991 116888
rect 880 116488 99991 116760
rect 880 116480 99120 116488
rect 13 116208 99120 116480
rect 13 115944 99991 116208
rect 880 115808 99991 115944
rect 880 115664 99120 115808
rect 13 115528 99120 115664
rect 13 115128 99991 115528
rect 880 114848 99120 115128
rect 13 114448 99991 114848
rect 13 114312 99120 114448
rect 880 114168 99120 114312
rect 880 114032 99991 114168
rect 13 113768 99991 114032
rect 13 113496 99120 113768
rect 880 113488 99120 113496
rect 880 113216 99991 113488
rect 13 113088 99991 113216
rect 13 112808 99120 113088
rect 13 112680 99991 112808
rect 880 112408 99991 112680
rect 880 112400 99120 112408
rect 13 112128 99120 112400
rect 13 111864 99991 112128
rect 880 111728 99991 111864
rect 880 111584 99120 111728
rect 13 111448 99120 111584
rect 13 111048 99991 111448
rect 880 110768 99120 111048
rect 13 110368 99991 110768
rect 13 110232 99120 110368
rect 880 110088 99120 110232
rect 880 109952 99991 110088
rect 13 109688 99991 109952
rect 13 109416 99120 109688
rect 880 109408 99120 109416
rect 880 109136 99991 109408
rect 13 109008 99991 109136
rect 13 108728 99120 109008
rect 13 108600 99991 108728
rect 880 108328 99991 108600
rect 880 108320 99120 108328
rect 13 108048 99120 108320
rect 13 107784 99991 108048
rect 880 107648 99991 107784
rect 880 107504 99120 107648
rect 13 107368 99120 107504
rect 13 106968 99991 107368
rect 880 106688 99120 106968
rect 13 106288 99991 106688
rect 13 106152 99120 106288
rect 880 106008 99120 106152
rect 880 105872 99991 106008
rect 13 105608 99991 105872
rect 13 105336 99120 105608
rect 880 105328 99120 105336
rect 880 105056 99991 105328
rect 13 104928 99991 105056
rect 13 104648 99120 104928
rect 13 104520 99991 104648
rect 880 104248 99991 104520
rect 880 104240 99120 104248
rect 13 103968 99120 104240
rect 13 103704 99991 103968
rect 880 103568 99991 103704
rect 880 103424 99120 103568
rect 13 103288 99120 103424
rect 13 102888 99991 103288
rect 880 102608 99120 102888
rect 13 102208 99991 102608
rect 13 102072 99120 102208
rect 880 101928 99120 102072
rect 880 101792 99991 101928
rect 13 101528 99991 101792
rect 13 101256 99120 101528
rect 880 101248 99120 101256
rect 880 100976 99991 101248
rect 13 100848 99991 100976
rect 13 100568 99120 100848
rect 13 100440 99991 100568
rect 880 100168 99991 100440
rect 880 100160 99120 100168
rect 13 99888 99120 100160
rect 13 99624 99991 99888
rect 880 99488 99991 99624
rect 880 99344 99120 99488
rect 13 99208 99120 99344
rect 13 98808 99991 99208
rect 880 98528 99120 98808
rect 13 98128 99991 98528
rect 13 97992 99120 98128
rect 880 97848 99120 97992
rect 880 97712 99991 97848
rect 13 97448 99991 97712
rect 13 97176 99120 97448
rect 880 97168 99120 97176
rect 880 96896 99991 97168
rect 13 96768 99991 96896
rect 13 96488 99120 96768
rect 13 96360 99991 96488
rect 880 96088 99991 96360
rect 880 96080 99120 96088
rect 13 95808 99120 96080
rect 13 95544 99991 95808
rect 880 95408 99991 95544
rect 880 95264 99120 95408
rect 13 95128 99120 95264
rect 13 94728 99991 95128
rect 880 94448 99120 94728
rect 13 94048 99991 94448
rect 13 93912 99120 94048
rect 880 93768 99120 93912
rect 880 93632 99991 93768
rect 13 93368 99991 93632
rect 13 93096 99120 93368
rect 880 93088 99120 93096
rect 880 92816 99991 93088
rect 13 92688 99991 92816
rect 13 92408 99120 92688
rect 13 92280 99991 92408
rect 880 92008 99991 92280
rect 880 92000 99120 92008
rect 13 91728 99120 92000
rect 13 91464 99991 91728
rect 880 91328 99991 91464
rect 880 91184 99120 91328
rect 13 91048 99120 91184
rect 13 90648 99991 91048
rect 880 90368 99120 90648
rect 13 89968 99991 90368
rect 13 89832 99120 89968
rect 880 89688 99120 89832
rect 880 89552 99991 89688
rect 13 89288 99991 89552
rect 13 89016 99120 89288
rect 880 89008 99120 89016
rect 880 88736 99991 89008
rect 13 88608 99991 88736
rect 13 88328 99120 88608
rect 13 88200 99991 88328
rect 880 87928 99991 88200
rect 880 87920 99120 87928
rect 13 87648 99120 87920
rect 13 87384 99991 87648
rect 880 87248 99991 87384
rect 880 87104 99120 87248
rect 13 86968 99120 87104
rect 13 86568 99991 86968
rect 880 86288 99120 86568
rect 13 85888 99991 86288
rect 13 85752 99120 85888
rect 880 85608 99120 85752
rect 880 85472 99991 85608
rect 13 85208 99991 85472
rect 13 84936 99120 85208
rect 880 84928 99120 84936
rect 880 84656 99991 84928
rect 13 84528 99991 84656
rect 13 84248 99120 84528
rect 13 84120 99991 84248
rect 880 83848 99991 84120
rect 880 83840 99120 83848
rect 13 83568 99120 83840
rect 13 83304 99991 83568
rect 880 83168 99991 83304
rect 880 83024 99120 83168
rect 13 82888 99120 83024
rect 13 82488 99991 82888
rect 880 82208 99120 82488
rect 13 81808 99991 82208
rect 13 81672 99120 81808
rect 880 81528 99120 81672
rect 880 81392 99991 81528
rect 13 81128 99991 81392
rect 13 80856 99120 81128
rect 880 80848 99120 80856
rect 880 80576 99991 80848
rect 13 80448 99991 80576
rect 13 80168 99120 80448
rect 13 80040 99991 80168
rect 880 79768 99991 80040
rect 880 79760 99120 79768
rect 13 79488 99120 79760
rect 13 79224 99991 79488
rect 880 79088 99991 79224
rect 880 78944 99120 79088
rect 13 78808 99120 78944
rect 13 78408 99991 78808
rect 880 78128 99120 78408
rect 13 77728 99991 78128
rect 13 77592 99120 77728
rect 880 77448 99120 77592
rect 880 77312 99991 77448
rect 13 77048 99991 77312
rect 13 76776 99120 77048
rect 880 76768 99120 76776
rect 880 76496 99991 76768
rect 13 76368 99991 76496
rect 13 76088 99120 76368
rect 13 75960 99991 76088
rect 880 75688 99991 75960
rect 880 75680 99120 75688
rect 13 75408 99120 75680
rect 13 75144 99991 75408
rect 880 75008 99991 75144
rect 880 74864 99120 75008
rect 13 74728 99120 74864
rect 13 74328 99991 74728
rect 880 74048 99120 74328
rect 13 73648 99991 74048
rect 13 73512 99120 73648
rect 880 73368 99120 73512
rect 880 73232 99991 73368
rect 13 72968 99991 73232
rect 13 72696 99120 72968
rect 880 72688 99120 72696
rect 880 72416 99991 72688
rect 13 72288 99991 72416
rect 13 72008 99120 72288
rect 13 71880 99991 72008
rect 880 71608 99991 71880
rect 880 71600 99120 71608
rect 13 71328 99120 71600
rect 13 71064 99991 71328
rect 880 70928 99991 71064
rect 880 70784 99120 70928
rect 13 70648 99120 70784
rect 13 70248 99991 70648
rect 880 69968 99120 70248
rect 13 69568 99991 69968
rect 13 69432 99120 69568
rect 880 69288 99120 69432
rect 880 69152 99991 69288
rect 13 68888 99991 69152
rect 13 68616 99120 68888
rect 880 68608 99120 68616
rect 880 68336 99991 68608
rect 13 68208 99991 68336
rect 13 67928 99120 68208
rect 13 67800 99991 67928
rect 880 67528 99991 67800
rect 880 67520 99120 67528
rect 13 67248 99120 67520
rect 13 66984 99991 67248
rect 880 66848 99991 66984
rect 880 66704 99120 66848
rect 13 66568 99120 66704
rect 13 66168 99991 66568
rect 880 65888 99120 66168
rect 13 65488 99991 65888
rect 13 65352 99120 65488
rect 880 65208 99120 65352
rect 880 65072 99991 65208
rect 13 64808 99991 65072
rect 13 64536 99120 64808
rect 880 64528 99120 64536
rect 880 64256 99991 64528
rect 13 64128 99991 64256
rect 13 63848 99120 64128
rect 13 63720 99991 63848
rect 880 63448 99991 63720
rect 880 63440 99120 63448
rect 13 63168 99120 63440
rect 13 62904 99991 63168
rect 880 62768 99991 62904
rect 880 62624 99120 62768
rect 13 62488 99120 62624
rect 13 62088 99991 62488
rect 880 61808 99120 62088
rect 13 61408 99991 61808
rect 13 61272 99120 61408
rect 880 61128 99120 61272
rect 880 60992 99991 61128
rect 13 60728 99991 60992
rect 13 60456 99120 60728
rect 880 60448 99120 60456
rect 880 60176 99991 60448
rect 13 60048 99991 60176
rect 13 59768 99120 60048
rect 13 59640 99991 59768
rect 880 59368 99991 59640
rect 880 59360 99120 59368
rect 13 59088 99120 59360
rect 13 58824 99991 59088
rect 880 58688 99991 58824
rect 880 58544 99120 58688
rect 13 58408 99120 58544
rect 13 58008 99991 58408
rect 880 57728 99120 58008
rect 13 57328 99991 57728
rect 13 57192 99120 57328
rect 880 57048 99120 57192
rect 880 56912 99991 57048
rect 13 56648 99991 56912
rect 13 56376 99120 56648
rect 880 56368 99120 56376
rect 880 56096 99991 56368
rect 13 55968 99991 56096
rect 13 55688 99120 55968
rect 13 55560 99991 55688
rect 880 55288 99991 55560
rect 880 55280 99120 55288
rect 13 55008 99120 55280
rect 13 54744 99991 55008
rect 880 54608 99991 54744
rect 880 54464 99120 54608
rect 13 54328 99120 54464
rect 13 53928 99991 54328
rect 880 53648 99120 53928
rect 13 53248 99991 53648
rect 13 53112 99120 53248
rect 880 52968 99120 53112
rect 880 52832 99991 52968
rect 13 52568 99991 52832
rect 13 52296 99120 52568
rect 880 52288 99120 52296
rect 880 52016 99991 52288
rect 13 51888 99991 52016
rect 13 51608 99120 51888
rect 13 51480 99991 51608
rect 880 51208 99991 51480
rect 880 51200 99120 51208
rect 13 50928 99120 51200
rect 13 50664 99991 50928
rect 880 50528 99991 50664
rect 880 50384 99120 50528
rect 13 50248 99120 50384
rect 13 49848 99991 50248
rect 880 49568 99120 49848
rect 13 49168 99991 49568
rect 13 49032 99120 49168
rect 880 48888 99120 49032
rect 880 48752 99991 48888
rect 13 48488 99991 48752
rect 13 48216 99120 48488
rect 880 48208 99120 48216
rect 880 47936 99991 48208
rect 13 47808 99991 47936
rect 13 47528 99120 47808
rect 13 47400 99991 47528
rect 880 47128 99991 47400
rect 880 47120 99120 47128
rect 13 46848 99120 47120
rect 13 46584 99991 46848
rect 880 46448 99991 46584
rect 880 46304 99120 46448
rect 13 46168 99120 46304
rect 13 45768 99991 46168
rect 880 45488 99120 45768
rect 13 45088 99991 45488
rect 13 44952 99120 45088
rect 880 44808 99120 44952
rect 880 44672 99991 44808
rect 13 44408 99991 44672
rect 13 44136 99120 44408
rect 880 44128 99120 44136
rect 880 43856 99991 44128
rect 13 43728 99991 43856
rect 13 43448 99120 43728
rect 13 43320 99991 43448
rect 880 43048 99991 43320
rect 880 43040 99120 43048
rect 13 42768 99120 43040
rect 13 42504 99991 42768
rect 880 42368 99991 42504
rect 880 42224 99120 42368
rect 13 42088 99120 42224
rect 13 41688 99991 42088
rect 880 41408 99120 41688
rect 13 41008 99991 41408
rect 13 40872 99120 41008
rect 880 40728 99120 40872
rect 880 40592 99991 40728
rect 13 40328 99991 40592
rect 13 40056 99120 40328
rect 880 40048 99120 40056
rect 880 39776 99991 40048
rect 13 39648 99991 39776
rect 13 39368 99120 39648
rect 13 39240 99991 39368
rect 880 38968 99991 39240
rect 880 38960 99120 38968
rect 13 38688 99120 38960
rect 13 38424 99991 38688
rect 880 38288 99991 38424
rect 880 38144 99120 38288
rect 13 38008 99120 38144
rect 13 37608 99991 38008
rect 880 37328 99120 37608
rect 13 36928 99991 37328
rect 13 36792 99120 36928
rect 880 36648 99120 36792
rect 880 36512 99991 36648
rect 13 36248 99991 36512
rect 13 35976 99120 36248
rect 880 35968 99120 35976
rect 880 35696 99991 35968
rect 13 35568 99991 35696
rect 13 35288 99120 35568
rect 13 35160 99991 35288
rect 880 34888 99991 35160
rect 880 34880 99120 34888
rect 13 34608 99120 34880
rect 13 34344 99991 34608
rect 880 34208 99991 34344
rect 880 34064 99120 34208
rect 13 33928 99120 34064
rect 13 33528 99991 33928
rect 880 33248 99120 33528
rect 13 32848 99991 33248
rect 13 32712 99120 32848
rect 880 32568 99120 32712
rect 880 32432 99991 32568
rect 13 32168 99991 32432
rect 13 31896 99120 32168
rect 880 31888 99120 31896
rect 880 31616 99991 31888
rect 13 31488 99991 31616
rect 13 31208 99120 31488
rect 13 31080 99991 31208
rect 880 30808 99991 31080
rect 880 30800 99120 30808
rect 13 30528 99120 30800
rect 13 30264 99991 30528
rect 880 30128 99991 30264
rect 880 29984 99120 30128
rect 13 29848 99120 29984
rect 13 29448 99991 29848
rect 880 29168 99120 29448
rect 13 28768 99991 29168
rect 13 28632 99120 28768
rect 880 28488 99120 28632
rect 880 28352 99991 28488
rect 13 28088 99991 28352
rect 13 27816 99120 28088
rect 880 27808 99120 27816
rect 880 27536 99991 27808
rect 13 27408 99991 27536
rect 13 27128 99120 27408
rect 13 27000 99991 27128
rect 880 26728 99991 27000
rect 880 26720 99120 26728
rect 13 26448 99120 26720
rect 13 26184 99991 26448
rect 880 26048 99991 26184
rect 880 25904 99120 26048
rect 13 25768 99120 25904
rect 13 25368 99991 25768
rect 880 25088 99120 25368
rect 13 24688 99991 25088
rect 13 24552 99120 24688
rect 880 24408 99120 24552
rect 880 24272 99991 24408
rect 13 24008 99991 24272
rect 13 23736 99120 24008
rect 880 23728 99120 23736
rect 880 23456 99991 23728
rect 13 23328 99991 23456
rect 13 23048 99120 23328
rect 13 22920 99991 23048
rect 880 22648 99991 22920
rect 880 22640 99120 22648
rect 13 22368 99120 22640
rect 13 22104 99991 22368
rect 880 21968 99991 22104
rect 880 21824 99120 21968
rect 13 21688 99120 21824
rect 13 21288 99991 21688
rect 880 21008 99120 21288
rect 13 20608 99991 21008
rect 13 20472 99120 20608
rect 880 20328 99120 20472
rect 880 20192 99991 20328
rect 13 19928 99991 20192
rect 13 19656 99120 19928
rect 880 19648 99120 19656
rect 880 19376 99991 19648
rect 13 19248 99991 19376
rect 13 18968 99120 19248
rect 13 18840 99991 18968
rect 880 18568 99991 18840
rect 880 18560 99120 18568
rect 13 18288 99120 18560
rect 13 18024 99991 18288
rect 880 17888 99991 18024
rect 880 17744 99120 17888
rect 13 17608 99120 17744
rect 13 17208 99991 17608
rect 880 16928 99120 17208
rect 13 16528 99991 16928
rect 13 16392 99120 16528
rect 880 16248 99120 16392
rect 880 16112 99991 16248
rect 13 15848 99991 16112
rect 13 15576 99120 15848
rect 880 15568 99120 15576
rect 880 15296 99991 15568
rect 13 15168 99991 15296
rect 13 14888 99120 15168
rect 13 14760 99991 14888
rect 880 14488 99991 14760
rect 880 14480 99120 14488
rect 13 14208 99120 14480
rect 13 13944 99991 14208
rect 880 13808 99991 13944
rect 880 13664 99120 13808
rect 13 13528 99120 13664
rect 13 13128 99991 13528
rect 880 12848 99120 13128
rect 13 12448 99991 12848
rect 13 12312 99120 12448
rect 880 12168 99120 12312
rect 880 12032 99991 12168
rect 13 11768 99991 12032
rect 13 11496 99120 11768
rect 880 11488 99120 11496
rect 880 11216 99991 11488
rect 13 10680 99991 11216
rect 880 10400 99991 10680
rect 13 9864 99991 10400
rect 880 9584 99991 9864
rect 13 9048 99991 9584
rect 880 8768 99991 9048
rect 13 8232 99991 8768
rect 880 7952 99991 8232
rect 13 7416 99991 7952
rect 880 7136 99991 7416
rect 13 6600 99991 7136
rect 880 6320 99991 6600
rect 13 5784 99991 6320
rect 880 5504 99991 5784
rect 13 4968 99991 5504
rect 880 4688 99991 4968
rect 13 4152 99991 4688
rect 880 3872 99991 4152
rect 13 3336 99991 3872
rect 880 3056 99991 3336
rect 13 2520 99991 3056
rect 880 2240 99991 2520
rect 13 1704 99991 2240
rect 880 1531 99991 1704
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
<< obsm4 >>
rect 427 2347 4128 156365
rect 4608 2347 19488 156365
rect 19968 2347 34848 156365
rect 35328 2347 50208 156365
rect 50688 2347 65568 156365
rect 66048 2347 80928 156365
rect 81408 2347 96288 156365
rect 96768 2347 99117 156365
<< labels >>
rlabel metal3 s 0 11296 800 11416 6 addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 12112 800 12232 6 addr0[1]
port 2 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 addr0[2]
port 3 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 addr0[3]
port 4 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 addr0[4]
port 5 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 addr0[5]
port 6 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 addr0[6]
port 7 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 addr0[7]
port 8 nsew signal output
rlabel metal3 s 0 17824 800 17944 6 addr0[8]
port 9 nsew signal output
rlabel metal3 s 0 99424 800 99544 6 addr1[0]
port 10 nsew signal output
rlabel metal3 s 0 100240 800 100360 6 addr1[1]
port 11 nsew signal output
rlabel metal3 s 0 101056 800 101176 6 addr1[2]
port 12 nsew signal output
rlabel metal3 s 0 101872 800 101992 6 addr1[3]
port 13 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 addr1[4]
port 14 nsew signal output
rlabel metal3 s 0 103504 800 103624 6 addr1[5]
port 15 nsew signal output
rlabel metal3 s 0 104320 800 104440 6 addr1[6]
port 16 nsew signal output
rlabel metal3 s 0 105136 800 105256 6 addr1[7]
port 17 nsew signal output
rlabel metal3 s 0 105952 800 106072 6 addr1[8]
port 18 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 clk0
port 19 nsew signal output
rlabel metal3 s 0 96976 800 97096 6 clk1
port 20 nsew signal output
rlabel metal2 s 2778 159200 2834 160000 6 coreIndex[0]
port 21 nsew signal input
rlabel metal2 s 5262 159200 5318 160000 6 coreIndex[1]
port 22 nsew signal input
rlabel metal2 s 7746 159200 7802 160000 6 coreIndex[2]
port 23 nsew signal input
rlabel metal2 s 10230 159200 10286 160000 6 coreIndex[3]
port 24 nsew signal input
rlabel metal2 s 12714 159200 12770 160000 6 coreIndex[4]
port 25 nsew signal input
rlabel metal2 s 15198 159200 15254 160000 6 coreIndex[5]
port 26 nsew signal input
rlabel metal2 s 17682 159200 17738 160000 6 coreIndex[6]
port 27 nsew signal input
rlabel metal2 s 20166 159200 20222 160000 6 coreIndex[7]
port 28 nsew signal input
rlabel metal3 s 99200 12928 100000 13048 6 core_wb_ack_i
port 29 nsew signal input
rlabel metal3 s 99200 17008 100000 17128 6 core_wb_adr_o[0]
port 30 nsew signal output
rlabel metal3 s 99200 40128 100000 40248 6 core_wb_adr_o[10]
port 31 nsew signal output
rlabel metal3 s 99200 42168 100000 42288 6 core_wb_adr_o[11]
port 32 nsew signal output
rlabel metal3 s 99200 44208 100000 44328 6 core_wb_adr_o[12]
port 33 nsew signal output
rlabel metal3 s 99200 46248 100000 46368 6 core_wb_adr_o[13]
port 34 nsew signal output
rlabel metal3 s 99200 48288 100000 48408 6 core_wb_adr_o[14]
port 35 nsew signal output
rlabel metal3 s 99200 50328 100000 50448 6 core_wb_adr_o[15]
port 36 nsew signal output
rlabel metal3 s 99200 52368 100000 52488 6 core_wb_adr_o[16]
port 37 nsew signal output
rlabel metal3 s 99200 54408 100000 54528 6 core_wb_adr_o[17]
port 38 nsew signal output
rlabel metal3 s 99200 56448 100000 56568 6 core_wb_adr_o[18]
port 39 nsew signal output
rlabel metal3 s 99200 58488 100000 58608 6 core_wb_adr_o[19]
port 40 nsew signal output
rlabel metal3 s 99200 19728 100000 19848 6 core_wb_adr_o[1]
port 41 nsew signal output
rlabel metal3 s 99200 60528 100000 60648 6 core_wb_adr_o[20]
port 42 nsew signal output
rlabel metal3 s 99200 62568 100000 62688 6 core_wb_adr_o[21]
port 43 nsew signal output
rlabel metal3 s 99200 64608 100000 64728 6 core_wb_adr_o[22]
port 44 nsew signal output
rlabel metal3 s 99200 66648 100000 66768 6 core_wb_adr_o[23]
port 45 nsew signal output
rlabel metal3 s 99200 68688 100000 68808 6 core_wb_adr_o[24]
port 46 nsew signal output
rlabel metal3 s 99200 70728 100000 70848 6 core_wb_adr_o[25]
port 47 nsew signal output
rlabel metal3 s 99200 72768 100000 72888 6 core_wb_adr_o[26]
port 48 nsew signal output
rlabel metal3 s 99200 74808 100000 74928 6 core_wb_adr_o[27]
port 49 nsew signal output
rlabel metal3 s 99200 22448 100000 22568 6 core_wb_adr_o[2]
port 50 nsew signal output
rlabel metal3 s 99200 25168 100000 25288 6 core_wb_adr_o[3]
port 51 nsew signal output
rlabel metal3 s 99200 27888 100000 28008 6 core_wb_adr_o[4]
port 52 nsew signal output
rlabel metal3 s 99200 29928 100000 30048 6 core_wb_adr_o[5]
port 53 nsew signal output
rlabel metal3 s 99200 31968 100000 32088 6 core_wb_adr_o[6]
port 54 nsew signal output
rlabel metal3 s 99200 34008 100000 34128 6 core_wb_adr_o[7]
port 55 nsew signal output
rlabel metal3 s 99200 36048 100000 36168 6 core_wb_adr_o[8]
port 56 nsew signal output
rlabel metal3 s 99200 38088 100000 38208 6 core_wb_adr_o[9]
port 57 nsew signal output
rlabel metal3 s 99200 13608 100000 13728 6 core_wb_cyc_o
port 58 nsew signal output
rlabel metal3 s 99200 17688 100000 17808 6 core_wb_data_i[0]
port 59 nsew signal input
rlabel metal3 s 99200 40808 100000 40928 6 core_wb_data_i[10]
port 60 nsew signal input
rlabel metal3 s 99200 42848 100000 42968 6 core_wb_data_i[11]
port 61 nsew signal input
rlabel metal3 s 99200 44888 100000 45008 6 core_wb_data_i[12]
port 62 nsew signal input
rlabel metal3 s 99200 46928 100000 47048 6 core_wb_data_i[13]
port 63 nsew signal input
rlabel metal3 s 99200 48968 100000 49088 6 core_wb_data_i[14]
port 64 nsew signal input
rlabel metal3 s 99200 51008 100000 51128 6 core_wb_data_i[15]
port 65 nsew signal input
rlabel metal3 s 99200 53048 100000 53168 6 core_wb_data_i[16]
port 66 nsew signal input
rlabel metal3 s 99200 55088 100000 55208 6 core_wb_data_i[17]
port 67 nsew signal input
rlabel metal3 s 99200 57128 100000 57248 6 core_wb_data_i[18]
port 68 nsew signal input
rlabel metal3 s 99200 59168 100000 59288 6 core_wb_data_i[19]
port 69 nsew signal input
rlabel metal3 s 99200 20408 100000 20528 6 core_wb_data_i[1]
port 70 nsew signal input
rlabel metal3 s 99200 61208 100000 61328 6 core_wb_data_i[20]
port 71 nsew signal input
rlabel metal3 s 99200 63248 100000 63368 6 core_wb_data_i[21]
port 72 nsew signal input
rlabel metal3 s 99200 65288 100000 65408 6 core_wb_data_i[22]
port 73 nsew signal input
rlabel metal3 s 99200 67328 100000 67448 6 core_wb_data_i[23]
port 74 nsew signal input
rlabel metal3 s 99200 69368 100000 69488 6 core_wb_data_i[24]
port 75 nsew signal input
rlabel metal3 s 99200 71408 100000 71528 6 core_wb_data_i[25]
port 76 nsew signal input
rlabel metal3 s 99200 73448 100000 73568 6 core_wb_data_i[26]
port 77 nsew signal input
rlabel metal3 s 99200 75488 100000 75608 6 core_wb_data_i[27]
port 78 nsew signal input
rlabel metal3 s 99200 76848 100000 76968 6 core_wb_data_i[28]
port 79 nsew signal input
rlabel metal3 s 99200 78208 100000 78328 6 core_wb_data_i[29]
port 80 nsew signal input
rlabel metal3 s 99200 23128 100000 23248 6 core_wb_data_i[2]
port 81 nsew signal input
rlabel metal3 s 99200 79568 100000 79688 6 core_wb_data_i[30]
port 82 nsew signal input
rlabel metal3 s 99200 80928 100000 81048 6 core_wb_data_i[31]
port 83 nsew signal input
rlabel metal3 s 99200 25848 100000 25968 6 core_wb_data_i[3]
port 84 nsew signal input
rlabel metal3 s 99200 28568 100000 28688 6 core_wb_data_i[4]
port 85 nsew signal input
rlabel metal3 s 99200 30608 100000 30728 6 core_wb_data_i[5]
port 86 nsew signal input
rlabel metal3 s 99200 32648 100000 32768 6 core_wb_data_i[6]
port 87 nsew signal input
rlabel metal3 s 99200 34688 100000 34808 6 core_wb_data_i[7]
port 88 nsew signal input
rlabel metal3 s 99200 36728 100000 36848 6 core_wb_data_i[8]
port 89 nsew signal input
rlabel metal3 s 99200 38768 100000 38888 6 core_wb_data_i[9]
port 90 nsew signal input
rlabel metal3 s 99200 18368 100000 18488 6 core_wb_data_o[0]
port 91 nsew signal output
rlabel metal3 s 99200 41488 100000 41608 6 core_wb_data_o[10]
port 92 nsew signal output
rlabel metal3 s 99200 43528 100000 43648 6 core_wb_data_o[11]
port 93 nsew signal output
rlabel metal3 s 99200 45568 100000 45688 6 core_wb_data_o[12]
port 94 nsew signal output
rlabel metal3 s 99200 47608 100000 47728 6 core_wb_data_o[13]
port 95 nsew signal output
rlabel metal3 s 99200 49648 100000 49768 6 core_wb_data_o[14]
port 96 nsew signal output
rlabel metal3 s 99200 51688 100000 51808 6 core_wb_data_o[15]
port 97 nsew signal output
rlabel metal3 s 99200 53728 100000 53848 6 core_wb_data_o[16]
port 98 nsew signal output
rlabel metal3 s 99200 55768 100000 55888 6 core_wb_data_o[17]
port 99 nsew signal output
rlabel metal3 s 99200 57808 100000 57928 6 core_wb_data_o[18]
port 100 nsew signal output
rlabel metal3 s 99200 59848 100000 59968 6 core_wb_data_o[19]
port 101 nsew signal output
rlabel metal3 s 99200 21088 100000 21208 6 core_wb_data_o[1]
port 102 nsew signal output
rlabel metal3 s 99200 61888 100000 62008 6 core_wb_data_o[20]
port 103 nsew signal output
rlabel metal3 s 99200 63928 100000 64048 6 core_wb_data_o[21]
port 104 nsew signal output
rlabel metal3 s 99200 65968 100000 66088 6 core_wb_data_o[22]
port 105 nsew signal output
rlabel metal3 s 99200 68008 100000 68128 6 core_wb_data_o[23]
port 106 nsew signal output
rlabel metal3 s 99200 70048 100000 70168 6 core_wb_data_o[24]
port 107 nsew signal output
rlabel metal3 s 99200 72088 100000 72208 6 core_wb_data_o[25]
port 108 nsew signal output
rlabel metal3 s 99200 74128 100000 74248 6 core_wb_data_o[26]
port 109 nsew signal output
rlabel metal3 s 99200 76168 100000 76288 6 core_wb_data_o[27]
port 110 nsew signal output
rlabel metal3 s 99200 77528 100000 77648 6 core_wb_data_o[28]
port 111 nsew signal output
rlabel metal3 s 99200 78888 100000 79008 6 core_wb_data_o[29]
port 112 nsew signal output
rlabel metal3 s 99200 23808 100000 23928 6 core_wb_data_o[2]
port 113 nsew signal output
rlabel metal3 s 99200 80248 100000 80368 6 core_wb_data_o[30]
port 114 nsew signal output
rlabel metal3 s 99200 81608 100000 81728 6 core_wb_data_o[31]
port 115 nsew signal output
rlabel metal3 s 99200 26528 100000 26648 6 core_wb_data_o[3]
port 116 nsew signal output
rlabel metal3 s 99200 29248 100000 29368 6 core_wb_data_o[4]
port 117 nsew signal output
rlabel metal3 s 99200 31288 100000 31408 6 core_wb_data_o[5]
port 118 nsew signal output
rlabel metal3 s 99200 33328 100000 33448 6 core_wb_data_o[6]
port 119 nsew signal output
rlabel metal3 s 99200 35368 100000 35488 6 core_wb_data_o[7]
port 120 nsew signal output
rlabel metal3 s 99200 37408 100000 37528 6 core_wb_data_o[8]
port 121 nsew signal output
rlabel metal3 s 99200 39448 100000 39568 6 core_wb_data_o[9]
port 122 nsew signal output
rlabel metal3 s 99200 14288 100000 14408 6 core_wb_error_i
port 123 nsew signal input
rlabel metal3 s 99200 19048 100000 19168 6 core_wb_sel_o[0]
port 124 nsew signal output
rlabel metal3 s 99200 21768 100000 21888 6 core_wb_sel_o[1]
port 125 nsew signal output
rlabel metal3 s 99200 24488 100000 24608 6 core_wb_sel_o[2]
port 126 nsew signal output
rlabel metal3 s 99200 27208 100000 27328 6 core_wb_sel_o[3]
port 127 nsew signal output
rlabel metal3 s 99200 14968 100000 15088 6 core_wb_stall_i
port 128 nsew signal input
rlabel metal3 s 99200 15648 100000 15768 6 core_wb_stb_o
port 129 nsew signal output
rlabel metal3 s 99200 16328 100000 16448 6 core_wb_we_o
port 130 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 csb0[0]
port 131 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 csb0[1]
port 132 nsew signal output
rlabel metal3 s 0 97792 800 97912 6 csb1[0]
port 133 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 csb1[1]
port 134 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 din0[0]
port 135 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 din0[10]
port 136 nsew signal output
rlabel metal3 s 0 27616 800 27736 6 din0[11]
port 137 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 din0[12]
port 138 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 din0[13]
port 139 nsew signal output
rlabel metal3 s 0 30064 800 30184 6 din0[14]
port 140 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 din0[15]
port 141 nsew signal output
rlabel metal3 s 0 31696 800 31816 6 din0[16]
port 142 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 din0[17]
port 143 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 din0[18]
port 144 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 din0[19]
port 145 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 din0[1]
port 146 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 din0[20]
port 147 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 din0[21]
port 148 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 din0[22]
port 149 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 din0[23]
port 150 nsew signal output
rlabel metal3 s 0 38224 800 38344 6 din0[24]
port 151 nsew signal output
rlabel metal3 s 0 39040 800 39160 6 din0[25]
port 152 nsew signal output
rlabel metal3 s 0 39856 800 39976 6 din0[26]
port 153 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 din0[27]
port 154 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 din0[28]
port 155 nsew signal output
rlabel metal3 s 0 42304 800 42424 6 din0[29]
port 156 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 din0[2]
port 157 nsew signal output
rlabel metal3 s 0 43120 800 43240 6 din0[30]
port 158 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 din0[31]
port 159 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 din0[3]
port 160 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 din0[4]
port 161 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 din0[5]
port 162 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 din0[6]
port 163 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 din0[7]
port 164 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 din0[8]
port 165 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 din0[9]
port 166 nsew signal output
rlabel metal3 s 0 44752 800 44872 6 dout0[0]
port 167 nsew signal input
rlabel metal3 s 0 52912 800 53032 6 dout0[10]
port 168 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 dout0[11]
port 169 nsew signal input
rlabel metal3 s 0 54544 800 54664 6 dout0[12]
port 170 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 dout0[13]
port 171 nsew signal input
rlabel metal3 s 0 56176 800 56296 6 dout0[14]
port 172 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 dout0[15]
port 173 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 dout0[16]
port 174 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 dout0[17]
port 175 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 dout0[18]
port 176 nsew signal input
rlabel metal3 s 0 60256 800 60376 6 dout0[19]
port 177 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 dout0[1]
port 178 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 dout0[20]
port 179 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 dout0[21]
port 180 nsew signal input
rlabel metal3 s 0 62704 800 62824 6 dout0[22]
port 181 nsew signal input
rlabel metal3 s 0 63520 800 63640 6 dout0[23]
port 182 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 dout0[24]
port 183 nsew signal input
rlabel metal3 s 0 65152 800 65272 6 dout0[25]
port 184 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 dout0[26]
port 185 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 dout0[27]
port 186 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 dout0[28]
port 187 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 dout0[29]
port 188 nsew signal input
rlabel metal3 s 0 46384 800 46504 6 dout0[2]
port 189 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 dout0[30]
port 190 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 dout0[31]
port 191 nsew signal input
rlabel metal3 s 0 70864 800 70984 6 dout0[32]
port 192 nsew signal input
rlabel metal3 s 0 71680 800 71800 6 dout0[33]
port 193 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 dout0[34]
port 194 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 dout0[35]
port 195 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 dout0[36]
port 196 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 dout0[37]
port 197 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 dout0[38]
port 198 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 dout0[39]
port 199 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 dout0[3]
port 200 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 dout0[40]
port 201 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 dout0[41]
port 202 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 dout0[42]
port 203 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 dout0[43]
port 204 nsew signal input
rlabel metal3 s 0 80656 800 80776 6 dout0[44]
port 205 nsew signal input
rlabel metal3 s 0 81472 800 81592 6 dout0[45]
port 206 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 dout0[46]
port 207 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 dout0[47]
port 208 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 dout0[48]
port 209 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 dout0[49]
port 210 nsew signal input
rlabel metal3 s 0 48016 800 48136 6 dout0[4]
port 211 nsew signal input
rlabel metal3 s 0 85552 800 85672 6 dout0[50]
port 212 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 dout0[51]
port 213 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 dout0[52]
port 214 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 dout0[53]
port 215 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 dout0[54]
port 216 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 dout0[55]
port 217 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 dout0[56]
port 218 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 dout0[57]
port 219 nsew signal input
rlabel metal3 s 0 92080 800 92200 6 dout0[58]
port 220 nsew signal input
rlabel metal3 s 0 92896 800 93016 6 dout0[59]
port 221 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 dout0[5]
port 222 nsew signal input
rlabel metal3 s 0 93712 800 93832 6 dout0[60]
port 223 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 dout0[61]
port 224 nsew signal input
rlabel metal3 s 0 95344 800 95464 6 dout0[62]
port 225 nsew signal input
rlabel metal3 s 0 96160 800 96280 6 dout0[63]
port 226 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 dout0[6]
port 227 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 dout0[7]
port 228 nsew signal input
rlabel metal3 s 0 51280 800 51400 6 dout0[8]
port 229 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 dout0[9]
port 230 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 dout1[0]
port 231 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 dout1[10]
port 232 nsew signal input
rlabel metal3 s 0 115744 800 115864 6 dout1[11]
port 233 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 dout1[12]
port 234 nsew signal input
rlabel metal3 s 0 117376 800 117496 6 dout1[13]
port 235 nsew signal input
rlabel metal3 s 0 118192 800 118312 6 dout1[14]
port 236 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 dout1[15]
port 237 nsew signal input
rlabel metal3 s 0 119824 800 119944 6 dout1[16]
port 238 nsew signal input
rlabel metal3 s 0 120640 800 120760 6 dout1[17]
port 239 nsew signal input
rlabel metal3 s 0 121456 800 121576 6 dout1[18]
port 240 nsew signal input
rlabel metal3 s 0 122272 800 122392 6 dout1[19]
port 241 nsew signal input
rlabel metal3 s 0 107584 800 107704 6 dout1[1]
port 242 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 dout1[20]
port 243 nsew signal input
rlabel metal3 s 0 123904 800 124024 6 dout1[21]
port 244 nsew signal input
rlabel metal3 s 0 124720 800 124840 6 dout1[22]
port 245 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 dout1[23]
port 246 nsew signal input
rlabel metal3 s 0 126352 800 126472 6 dout1[24]
port 247 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 dout1[25]
port 248 nsew signal input
rlabel metal3 s 0 127984 800 128104 6 dout1[26]
port 249 nsew signal input
rlabel metal3 s 0 128800 800 128920 6 dout1[27]
port 250 nsew signal input
rlabel metal3 s 0 129616 800 129736 6 dout1[28]
port 251 nsew signal input
rlabel metal3 s 0 130432 800 130552 6 dout1[29]
port 252 nsew signal input
rlabel metal3 s 0 108400 800 108520 6 dout1[2]
port 253 nsew signal input
rlabel metal3 s 0 131248 800 131368 6 dout1[30]
port 254 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 dout1[31]
port 255 nsew signal input
rlabel metal3 s 0 132880 800 133000 6 dout1[32]
port 256 nsew signal input
rlabel metal3 s 0 133696 800 133816 6 dout1[33]
port 257 nsew signal input
rlabel metal3 s 0 134512 800 134632 6 dout1[34]
port 258 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 dout1[35]
port 259 nsew signal input
rlabel metal3 s 0 136144 800 136264 6 dout1[36]
port 260 nsew signal input
rlabel metal3 s 0 136960 800 137080 6 dout1[37]
port 261 nsew signal input
rlabel metal3 s 0 137776 800 137896 6 dout1[38]
port 262 nsew signal input
rlabel metal3 s 0 138592 800 138712 6 dout1[39]
port 263 nsew signal input
rlabel metal3 s 0 109216 800 109336 6 dout1[3]
port 264 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 dout1[40]
port 265 nsew signal input
rlabel metal3 s 0 140224 800 140344 6 dout1[41]
port 266 nsew signal input
rlabel metal3 s 0 141040 800 141160 6 dout1[42]
port 267 nsew signal input
rlabel metal3 s 0 141856 800 141976 6 dout1[43]
port 268 nsew signal input
rlabel metal3 s 0 142672 800 142792 6 dout1[44]
port 269 nsew signal input
rlabel metal3 s 0 143488 800 143608 6 dout1[45]
port 270 nsew signal input
rlabel metal3 s 0 144304 800 144424 6 dout1[46]
port 271 nsew signal input
rlabel metal3 s 0 145120 800 145240 6 dout1[47]
port 272 nsew signal input
rlabel metal3 s 0 145936 800 146056 6 dout1[48]
port 273 nsew signal input
rlabel metal3 s 0 146752 800 146872 6 dout1[49]
port 274 nsew signal input
rlabel metal3 s 0 110032 800 110152 6 dout1[4]
port 275 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 dout1[50]
port 276 nsew signal input
rlabel metal3 s 0 148384 800 148504 6 dout1[51]
port 277 nsew signal input
rlabel metal3 s 0 149200 800 149320 6 dout1[52]
port 278 nsew signal input
rlabel metal3 s 0 150016 800 150136 6 dout1[53]
port 279 nsew signal input
rlabel metal3 s 0 150832 800 150952 6 dout1[54]
port 280 nsew signal input
rlabel metal3 s 0 151648 800 151768 6 dout1[55]
port 281 nsew signal input
rlabel metal3 s 0 152464 800 152584 6 dout1[56]
port 282 nsew signal input
rlabel metal3 s 0 153280 800 153400 6 dout1[57]
port 283 nsew signal input
rlabel metal3 s 0 154096 800 154216 6 dout1[58]
port 284 nsew signal input
rlabel metal3 s 0 154912 800 155032 6 dout1[59]
port 285 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 dout1[5]
port 286 nsew signal input
rlabel metal3 s 0 155728 800 155848 6 dout1[60]
port 287 nsew signal input
rlabel metal3 s 0 156544 800 156664 6 dout1[61]
port 288 nsew signal input
rlabel metal3 s 0 157360 800 157480 6 dout1[62]
port 289 nsew signal input
rlabel metal3 s 0 158176 800 158296 6 dout1[63]
port 290 nsew signal input
rlabel metal3 s 0 111664 800 111784 6 dout1[6]
port 291 nsew signal input
rlabel metal3 s 0 112480 800 112600 6 dout1[7]
port 292 nsew signal input
rlabel metal3 s 0 113296 800 113416 6 dout1[8]
port 293 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 dout1[9]
port 294 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 irq[0]
port 295 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 irq[10]
port 296 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 irq[11]
port 297 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 irq[12]
port 298 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 irq[13]
port 299 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 irq[14]
port 300 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 irq[15]
port 301 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 irq[1]
port 302 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 irq[2]
port 303 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 irq[3]
port 304 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 irq[4]
port 305 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 irq[5]
port 306 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 irq[6]
port 307 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 irq[7]
port 308 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 irq[8]
port 309 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 irq[9]
port 310 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 jtag_tck
port 311 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 jtag_tdi
port 312 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 jtag_tdo
port 313 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 jtag_tms
port 314 nsew signal input
rlabel metal3 s 99200 82288 100000 82408 6 localMemory_wb_ack_o
port 315 nsew signal output
rlabel metal3 s 99200 86368 100000 86488 6 localMemory_wb_adr_i[0]
port 316 nsew signal input
rlabel metal3 s 99200 109488 100000 109608 6 localMemory_wb_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 99200 111528 100000 111648 6 localMemory_wb_adr_i[11]
port 318 nsew signal input
rlabel metal3 s 99200 113568 100000 113688 6 localMemory_wb_adr_i[12]
port 319 nsew signal input
rlabel metal3 s 99200 115608 100000 115728 6 localMemory_wb_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 99200 117648 100000 117768 6 localMemory_wb_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 99200 119688 100000 119808 6 localMemory_wb_adr_i[15]
port 322 nsew signal input
rlabel metal3 s 99200 121728 100000 121848 6 localMemory_wb_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 99200 123768 100000 123888 6 localMemory_wb_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 99200 125808 100000 125928 6 localMemory_wb_adr_i[18]
port 325 nsew signal input
rlabel metal3 s 99200 127848 100000 127968 6 localMemory_wb_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 99200 89088 100000 89208 6 localMemory_wb_adr_i[1]
port 327 nsew signal input
rlabel metal3 s 99200 129888 100000 130008 6 localMemory_wb_adr_i[20]
port 328 nsew signal input
rlabel metal3 s 99200 131928 100000 132048 6 localMemory_wb_adr_i[21]
port 329 nsew signal input
rlabel metal3 s 99200 133968 100000 134088 6 localMemory_wb_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 99200 136008 100000 136128 6 localMemory_wb_adr_i[23]
port 331 nsew signal input
rlabel metal3 s 99200 91808 100000 91928 6 localMemory_wb_adr_i[2]
port 332 nsew signal input
rlabel metal3 s 99200 94528 100000 94648 6 localMemory_wb_adr_i[3]
port 333 nsew signal input
rlabel metal3 s 99200 97248 100000 97368 6 localMemory_wb_adr_i[4]
port 334 nsew signal input
rlabel metal3 s 99200 99288 100000 99408 6 localMemory_wb_adr_i[5]
port 335 nsew signal input
rlabel metal3 s 99200 101328 100000 101448 6 localMemory_wb_adr_i[6]
port 336 nsew signal input
rlabel metal3 s 99200 103368 100000 103488 6 localMemory_wb_adr_i[7]
port 337 nsew signal input
rlabel metal3 s 99200 105408 100000 105528 6 localMemory_wb_adr_i[8]
port 338 nsew signal input
rlabel metal3 s 99200 107448 100000 107568 6 localMemory_wb_adr_i[9]
port 339 nsew signal input
rlabel metal3 s 99200 82968 100000 83088 6 localMemory_wb_cyc_i
port 340 nsew signal input
rlabel metal3 s 99200 87048 100000 87168 6 localMemory_wb_data_i[0]
port 341 nsew signal input
rlabel metal3 s 99200 110168 100000 110288 6 localMemory_wb_data_i[10]
port 342 nsew signal input
rlabel metal3 s 99200 112208 100000 112328 6 localMemory_wb_data_i[11]
port 343 nsew signal input
rlabel metal3 s 99200 114248 100000 114368 6 localMemory_wb_data_i[12]
port 344 nsew signal input
rlabel metal3 s 99200 116288 100000 116408 6 localMemory_wb_data_i[13]
port 345 nsew signal input
rlabel metal3 s 99200 118328 100000 118448 6 localMemory_wb_data_i[14]
port 346 nsew signal input
rlabel metal3 s 99200 120368 100000 120488 6 localMemory_wb_data_i[15]
port 347 nsew signal input
rlabel metal3 s 99200 122408 100000 122528 6 localMemory_wb_data_i[16]
port 348 nsew signal input
rlabel metal3 s 99200 124448 100000 124568 6 localMemory_wb_data_i[17]
port 349 nsew signal input
rlabel metal3 s 99200 126488 100000 126608 6 localMemory_wb_data_i[18]
port 350 nsew signal input
rlabel metal3 s 99200 128528 100000 128648 6 localMemory_wb_data_i[19]
port 351 nsew signal input
rlabel metal3 s 99200 89768 100000 89888 6 localMemory_wb_data_i[1]
port 352 nsew signal input
rlabel metal3 s 99200 130568 100000 130688 6 localMemory_wb_data_i[20]
port 353 nsew signal input
rlabel metal3 s 99200 132608 100000 132728 6 localMemory_wb_data_i[21]
port 354 nsew signal input
rlabel metal3 s 99200 134648 100000 134768 6 localMemory_wb_data_i[22]
port 355 nsew signal input
rlabel metal3 s 99200 136688 100000 136808 6 localMemory_wb_data_i[23]
port 356 nsew signal input
rlabel metal3 s 99200 138048 100000 138168 6 localMemory_wb_data_i[24]
port 357 nsew signal input
rlabel metal3 s 99200 139408 100000 139528 6 localMemory_wb_data_i[25]
port 358 nsew signal input
rlabel metal3 s 99200 140768 100000 140888 6 localMemory_wb_data_i[26]
port 359 nsew signal input
rlabel metal3 s 99200 142128 100000 142248 6 localMemory_wb_data_i[27]
port 360 nsew signal input
rlabel metal3 s 99200 143488 100000 143608 6 localMemory_wb_data_i[28]
port 361 nsew signal input
rlabel metal3 s 99200 144848 100000 144968 6 localMemory_wb_data_i[29]
port 362 nsew signal input
rlabel metal3 s 99200 92488 100000 92608 6 localMemory_wb_data_i[2]
port 363 nsew signal input
rlabel metal3 s 99200 146208 100000 146328 6 localMemory_wb_data_i[30]
port 364 nsew signal input
rlabel metal3 s 99200 147568 100000 147688 6 localMemory_wb_data_i[31]
port 365 nsew signal input
rlabel metal3 s 99200 95208 100000 95328 6 localMemory_wb_data_i[3]
port 366 nsew signal input
rlabel metal3 s 99200 97928 100000 98048 6 localMemory_wb_data_i[4]
port 367 nsew signal input
rlabel metal3 s 99200 99968 100000 100088 6 localMemory_wb_data_i[5]
port 368 nsew signal input
rlabel metal3 s 99200 102008 100000 102128 6 localMemory_wb_data_i[6]
port 369 nsew signal input
rlabel metal3 s 99200 104048 100000 104168 6 localMemory_wb_data_i[7]
port 370 nsew signal input
rlabel metal3 s 99200 106088 100000 106208 6 localMemory_wb_data_i[8]
port 371 nsew signal input
rlabel metal3 s 99200 108128 100000 108248 6 localMemory_wb_data_i[9]
port 372 nsew signal input
rlabel metal3 s 99200 87728 100000 87848 6 localMemory_wb_data_o[0]
port 373 nsew signal output
rlabel metal3 s 99200 110848 100000 110968 6 localMemory_wb_data_o[10]
port 374 nsew signal output
rlabel metal3 s 99200 112888 100000 113008 6 localMemory_wb_data_o[11]
port 375 nsew signal output
rlabel metal3 s 99200 114928 100000 115048 6 localMemory_wb_data_o[12]
port 376 nsew signal output
rlabel metal3 s 99200 116968 100000 117088 6 localMemory_wb_data_o[13]
port 377 nsew signal output
rlabel metal3 s 99200 119008 100000 119128 6 localMemory_wb_data_o[14]
port 378 nsew signal output
rlabel metal3 s 99200 121048 100000 121168 6 localMemory_wb_data_o[15]
port 379 nsew signal output
rlabel metal3 s 99200 123088 100000 123208 6 localMemory_wb_data_o[16]
port 380 nsew signal output
rlabel metal3 s 99200 125128 100000 125248 6 localMemory_wb_data_o[17]
port 381 nsew signal output
rlabel metal3 s 99200 127168 100000 127288 6 localMemory_wb_data_o[18]
port 382 nsew signal output
rlabel metal3 s 99200 129208 100000 129328 6 localMemory_wb_data_o[19]
port 383 nsew signal output
rlabel metal3 s 99200 90448 100000 90568 6 localMemory_wb_data_o[1]
port 384 nsew signal output
rlabel metal3 s 99200 131248 100000 131368 6 localMemory_wb_data_o[20]
port 385 nsew signal output
rlabel metal3 s 99200 133288 100000 133408 6 localMemory_wb_data_o[21]
port 386 nsew signal output
rlabel metal3 s 99200 135328 100000 135448 6 localMemory_wb_data_o[22]
port 387 nsew signal output
rlabel metal3 s 99200 137368 100000 137488 6 localMemory_wb_data_o[23]
port 388 nsew signal output
rlabel metal3 s 99200 138728 100000 138848 6 localMemory_wb_data_o[24]
port 389 nsew signal output
rlabel metal3 s 99200 140088 100000 140208 6 localMemory_wb_data_o[25]
port 390 nsew signal output
rlabel metal3 s 99200 141448 100000 141568 6 localMemory_wb_data_o[26]
port 391 nsew signal output
rlabel metal3 s 99200 142808 100000 142928 6 localMemory_wb_data_o[27]
port 392 nsew signal output
rlabel metal3 s 99200 144168 100000 144288 6 localMemory_wb_data_o[28]
port 393 nsew signal output
rlabel metal3 s 99200 145528 100000 145648 6 localMemory_wb_data_o[29]
port 394 nsew signal output
rlabel metal3 s 99200 93168 100000 93288 6 localMemory_wb_data_o[2]
port 395 nsew signal output
rlabel metal3 s 99200 146888 100000 147008 6 localMemory_wb_data_o[30]
port 396 nsew signal output
rlabel metal3 s 99200 148248 100000 148368 6 localMemory_wb_data_o[31]
port 397 nsew signal output
rlabel metal3 s 99200 95888 100000 96008 6 localMemory_wb_data_o[3]
port 398 nsew signal output
rlabel metal3 s 99200 98608 100000 98728 6 localMemory_wb_data_o[4]
port 399 nsew signal output
rlabel metal3 s 99200 100648 100000 100768 6 localMemory_wb_data_o[5]
port 400 nsew signal output
rlabel metal3 s 99200 102688 100000 102808 6 localMemory_wb_data_o[6]
port 401 nsew signal output
rlabel metal3 s 99200 104728 100000 104848 6 localMemory_wb_data_o[7]
port 402 nsew signal output
rlabel metal3 s 99200 106768 100000 106888 6 localMemory_wb_data_o[8]
port 403 nsew signal output
rlabel metal3 s 99200 108808 100000 108928 6 localMemory_wb_data_o[9]
port 404 nsew signal output
rlabel metal3 s 99200 83648 100000 83768 6 localMemory_wb_error_o
port 405 nsew signal output
rlabel metal3 s 99200 88408 100000 88528 6 localMemory_wb_sel_i[0]
port 406 nsew signal input
rlabel metal3 s 99200 91128 100000 91248 6 localMemory_wb_sel_i[1]
port 407 nsew signal input
rlabel metal3 s 99200 93848 100000 93968 6 localMemory_wb_sel_i[2]
port 408 nsew signal input
rlabel metal3 s 99200 96568 100000 96688 6 localMemory_wb_sel_i[3]
port 409 nsew signal input
rlabel metal3 s 99200 84328 100000 84448 6 localMemory_wb_stall_o
port 410 nsew signal output
rlabel metal3 s 99200 85008 100000 85128 6 localMemory_wb_stb_i
port 411 nsew signal input
rlabel metal3 s 99200 85688 100000 85808 6 localMemory_wb_we_i
port 412 nsew signal input
rlabel metal2 s 22650 159200 22706 160000 6 manufacturerID[0]
port 413 nsew signal input
rlabel metal2 s 47490 159200 47546 160000 6 manufacturerID[10]
port 414 nsew signal input
rlabel metal2 s 25134 159200 25190 160000 6 manufacturerID[1]
port 415 nsew signal input
rlabel metal2 s 27618 159200 27674 160000 6 manufacturerID[2]
port 416 nsew signal input
rlabel metal2 s 30102 159200 30158 160000 6 manufacturerID[3]
port 417 nsew signal input
rlabel metal2 s 32586 159200 32642 160000 6 manufacturerID[4]
port 418 nsew signal input
rlabel metal2 s 35070 159200 35126 160000 6 manufacturerID[5]
port 419 nsew signal input
rlabel metal2 s 37554 159200 37610 160000 6 manufacturerID[6]
port 420 nsew signal input
rlabel metal2 s 40038 159200 40094 160000 6 manufacturerID[7]
port 421 nsew signal input
rlabel metal2 s 42522 159200 42578 160000 6 manufacturerID[8]
port 422 nsew signal input
rlabel metal2 s 45006 159200 45062 160000 6 manufacturerID[9]
port 423 nsew signal input
rlabel metal2 s 49974 159200 50030 160000 6 partID[0]
port 424 nsew signal input
rlabel metal2 s 74814 159200 74870 160000 6 partID[10]
port 425 nsew signal input
rlabel metal2 s 77298 159200 77354 160000 6 partID[11]
port 426 nsew signal input
rlabel metal2 s 79782 159200 79838 160000 6 partID[12]
port 427 nsew signal input
rlabel metal2 s 82266 159200 82322 160000 6 partID[13]
port 428 nsew signal input
rlabel metal2 s 84750 159200 84806 160000 6 partID[14]
port 429 nsew signal input
rlabel metal2 s 87234 159200 87290 160000 6 partID[15]
port 430 nsew signal input
rlabel metal2 s 52458 159200 52514 160000 6 partID[1]
port 431 nsew signal input
rlabel metal2 s 54942 159200 54998 160000 6 partID[2]
port 432 nsew signal input
rlabel metal2 s 57426 159200 57482 160000 6 partID[3]
port 433 nsew signal input
rlabel metal2 s 59910 159200 59966 160000 6 partID[4]
port 434 nsew signal input
rlabel metal2 s 62394 159200 62450 160000 6 partID[5]
port 435 nsew signal input
rlabel metal2 s 64878 159200 64934 160000 6 partID[6]
port 436 nsew signal input
rlabel metal2 s 67362 159200 67418 160000 6 partID[7]
port 437 nsew signal input
rlabel metal2 s 69846 159200 69902 160000 6 partID[8]
port 438 nsew signal input
rlabel metal2 s 72330 159200 72386 160000 6 partID[9]
port 439 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 probe_env[0]
port 440 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 probe_env[1]
port 441 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 probe_jtagInstruction[0]
port 442 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 probe_jtagInstruction[1]
port 443 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 probe_jtagInstruction[2]
port 444 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 probe_jtagInstruction[3]
port 445 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 probe_jtagInstruction[4]
port 446 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 probe_programCounter[0]
port 447 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 probe_programCounter[10]
port 448 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 probe_programCounter[11]
port 449 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 probe_programCounter[12]
port 450 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 probe_programCounter[13]
port 451 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 probe_programCounter[14]
port 452 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 probe_programCounter[15]
port 453 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 probe_programCounter[16]
port 454 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 probe_programCounter[17]
port 455 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 probe_programCounter[18]
port 456 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 probe_programCounter[19]
port 457 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 probe_programCounter[1]
port 458 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 probe_programCounter[20]
port 459 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 probe_programCounter[21]
port 460 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 probe_programCounter[22]
port 461 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 probe_programCounter[23]
port 462 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 probe_programCounter[24]
port 463 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 probe_programCounter[25]
port 464 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 probe_programCounter[26]
port 465 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 probe_programCounter[27]
port 466 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 probe_programCounter[28]
port 467 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 probe_programCounter[29]
port 468 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 probe_programCounter[2]
port 469 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 probe_programCounter[30]
port 470 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 probe_programCounter[31]
port 471 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 probe_programCounter[3]
port 472 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 probe_programCounter[4]
port 473 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 probe_programCounter[5]
port 474 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 probe_programCounter[6]
port 475 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 probe_programCounter[7]
port 476 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 probe_programCounter[8]
port 477 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 probe_programCounter[9]
port 478 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 probe_state
port 479 nsew signal output
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 480 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 480 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 480 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 480 nsew power bidirectional
rlabel metal2 s 89718 159200 89774 160000 6 versionID[0]
port 481 nsew signal input
rlabel metal2 s 92202 159200 92258 160000 6 versionID[1]
port 482 nsew signal input
rlabel metal2 s 94686 159200 94742 160000 6 versionID[2]
port 483 nsew signal input
rlabel metal2 s 97170 159200 97226 160000 6 versionID[3]
port 484 nsew signal input
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 485 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 485 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 485 nsew ground bidirectional
rlabel metal3 s 99200 11568 100000 11688 6 wb_clk_i
port 486 nsew signal input
rlabel metal3 s 99200 12248 100000 12368 6 wb_rst_i
port 487 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 web0
port 488 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 wmask0[0]
port 489 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 wmask0[1]
port 490 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 wmask0[2]
port 491 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 wmask0[3]
port 492 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 44219316
string GDS_FILE /mnt/f/WSL/ASIC/ExperiarSoC/openlane/ExperiarCore/runs/23_05_26_11_29/results/signoff/ExperiarCore.magic.gds
string GDS_START 1622128
<< end >>

