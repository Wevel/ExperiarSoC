VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Peripherals
  CLASS BLOCK ;
  FOREIGN Peripherals ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 850.000 ;
  PIN flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END flash_csb
  PIN flash_io0_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END flash_io0_read
  PIN flash_io0_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END flash_io0_we
  PIN flash_io0_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END flash_io0_write
  PIN flash_io1_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END flash_io1_read
  PIN flash_io1_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END flash_io1_we
  PIN flash_io1_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END flash_io1_write
  PIN flash_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END flash_sck
  PIN internal_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END internal_uart_rx
  PIN internal_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END internal_uart_tx
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 846.000 4.050 850.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 846.000 82.710 850.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 846.000 90.530 850.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 846.000 98.350 850.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 846.000 106.630 850.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 846.000 114.450 850.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 846.000 122.270 850.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 846.000 130.090 850.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 846.000 137.910 850.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 846.000 145.730 850.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 846.000 154.010 850.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 846.000 11.870 850.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 846.000 161.830 850.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 846.000 169.650 850.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 846.000 177.470 850.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 846.000 185.290 850.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 846.000 193.110 850.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 846.000 200.930 850.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 846.000 209.210 850.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 846.000 217.030 850.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 846.000 224.850 850.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 846.000 232.670 850.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 846.000 19.690 850.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 846.000 240.490 850.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 846.000 248.310 850.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 846.000 256.590 850.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 846.000 264.410 850.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 846.000 272.230 850.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 846.000 280.050 850.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 846.000 287.870 850.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 846.000 295.690 850.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 846.000 27.510 850.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 846.000 35.330 850.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 846.000 43.150 850.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 846.000 50.970 850.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 846.000 59.250 850.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 846.000 67.070 850.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 846.000 74.890 850.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 846.000 303.970 850.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 846.000 382.630 850.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 846.000 390.450 850.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 846.000 398.270 850.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 846.000 406.550 850.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 846.000 414.370 850.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 846.000 422.190 850.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 846.000 430.010 850.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 846.000 437.830 850.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 846.000 445.650 850.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 846.000 453.930 850.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 846.000 311.790 850.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 846.000 461.750 850.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 846.000 469.570 850.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 846.000 477.390 850.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 846.000 485.210 850.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 846.000 493.030 850.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 846.000 500.850 850.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 846.000 509.130 850.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 846.000 516.950 850.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 846.000 524.770 850.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 846.000 532.590 850.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 846.000 319.610 850.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 846.000 540.410 850.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 846.000 548.230 850.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 846.000 556.510 850.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 846.000 564.330 850.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 846.000 572.150 850.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 846.000 579.970 850.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 846.000 587.790 850.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 846.000 595.610 850.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 846.000 327.430 850.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 846.000 335.250 850.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 846.000 343.070 850.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 846.000 350.890 850.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 846.000 359.170 850.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 846.000 366.990 850.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 846.000 374.810 850.000 ;
    END
  END io_out[9]
  PIN jtag_tck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 353.640 600.000 354.240 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 495.760 600.000 496.360 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 637.200 600.000 637.800 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 778.640 600.000 779.240 ;
    END
  END jtag_tms
  PIN probe_blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 70.760 600.000 71.360 ;
    END
  END probe_blink[0]
  PIN probe_blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 212.200 600.000 212.800 ;
    END
  END probe_blink[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 838.000 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 838.000 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.280 4.000 539.880 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.120 4.000 565.720 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.280 4.000 641.880 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.120 4.000 667.720 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.280 4.000 692.880 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.280 4.000 675.880 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.120 4.000 701.720 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.120 4.000 735.720 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.120 4.000 769.720 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.120 4.000 803.720 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 4.000 820.720 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.120 4.000 837.720 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.280 4.000 505.880 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.280 4.000 607.880 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.120 4.000 633.720 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.280 4.000 709.880 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.280 4.000 777.880 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 4.000 794.880 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.280 4.000 811.880 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.280 4.000 845.880 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 837.845 ;
      LAYER met1 ;
        RECT 5.130 8.200 597.470 839.080 ;
      LAYER met2 ;
        RECT 5.160 845.720 11.310 846.330 ;
        RECT 12.150 845.720 19.130 846.330 ;
        RECT 19.970 845.720 26.950 846.330 ;
        RECT 27.790 845.720 34.770 846.330 ;
        RECT 35.610 845.720 42.590 846.330 ;
        RECT 43.430 845.720 50.410 846.330 ;
        RECT 51.250 845.720 58.690 846.330 ;
        RECT 59.530 845.720 66.510 846.330 ;
        RECT 67.350 845.720 74.330 846.330 ;
        RECT 75.170 845.720 82.150 846.330 ;
        RECT 82.990 845.720 89.970 846.330 ;
        RECT 90.810 845.720 97.790 846.330 ;
        RECT 98.630 845.720 106.070 846.330 ;
        RECT 106.910 845.720 113.890 846.330 ;
        RECT 114.730 845.720 121.710 846.330 ;
        RECT 122.550 845.720 129.530 846.330 ;
        RECT 130.370 845.720 137.350 846.330 ;
        RECT 138.190 845.720 145.170 846.330 ;
        RECT 146.010 845.720 153.450 846.330 ;
        RECT 154.290 845.720 161.270 846.330 ;
        RECT 162.110 845.720 169.090 846.330 ;
        RECT 169.930 845.720 176.910 846.330 ;
        RECT 177.750 845.720 184.730 846.330 ;
        RECT 185.570 845.720 192.550 846.330 ;
        RECT 193.390 845.720 200.370 846.330 ;
        RECT 201.210 845.720 208.650 846.330 ;
        RECT 209.490 845.720 216.470 846.330 ;
        RECT 217.310 845.720 224.290 846.330 ;
        RECT 225.130 845.720 232.110 846.330 ;
        RECT 232.950 845.720 239.930 846.330 ;
        RECT 240.770 845.720 247.750 846.330 ;
        RECT 248.590 845.720 256.030 846.330 ;
        RECT 256.870 845.720 263.850 846.330 ;
        RECT 264.690 845.720 271.670 846.330 ;
        RECT 272.510 845.720 279.490 846.330 ;
        RECT 280.330 845.720 287.310 846.330 ;
        RECT 288.150 845.720 295.130 846.330 ;
        RECT 295.970 845.720 303.410 846.330 ;
        RECT 304.250 845.720 311.230 846.330 ;
        RECT 312.070 845.720 319.050 846.330 ;
        RECT 319.890 845.720 326.870 846.330 ;
        RECT 327.710 845.720 334.690 846.330 ;
        RECT 335.530 845.720 342.510 846.330 ;
        RECT 343.350 845.720 350.330 846.330 ;
        RECT 351.170 845.720 358.610 846.330 ;
        RECT 359.450 845.720 366.430 846.330 ;
        RECT 367.270 845.720 374.250 846.330 ;
        RECT 375.090 845.720 382.070 846.330 ;
        RECT 382.910 845.720 389.890 846.330 ;
        RECT 390.730 845.720 397.710 846.330 ;
        RECT 398.550 845.720 405.990 846.330 ;
        RECT 406.830 845.720 413.810 846.330 ;
        RECT 414.650 845.720 421.630 846.330 ;
        RECT 422.470 845.720 429.450 846.330 ;
        RECT 430.290 845.720 437.270 846.330 ;
        RECT 438.110 845.720 445.090 846.330 ;
        RECT 445.930 845.720 453.370 846.330 ;
        RECT 454.210 845.720 461.190 846.330 ;
        RECT 462.030 845.720 469.010 846.330 ;
        RECT 469.850 845.720 476.830 846.330 ;
        RECT 477.670 845.720 484.650 846.330 ;
        RECT 485.490 845.720 492.470 846.330 ;
        RECT 493.310 845.720 500.290 846.330 ;
        RECT 501.130 845.720 508.570 846.330 ;
        RECT 509.410 845.720 516.390 846.330 ;
        RECT 517.230 845.720 524.210 846.330 ;
        RECT 525.050 845.720 532.030 846.330 ;
        RECT 532.870 845.720 539.850 846.330 ;
        RECT 540.690 845.720 547.670 846.330 ;
        RECT 548.510 845.720 555.950 846.330 ;
        RECT 556.790 845.720 563.770 846.330 ;
        RECT 564.610 845.720 571.590 846.330 ;
        RECT 572.430 845.720 579.410 846.330 ;
        RECT 580.250 845.720 587.230 846.330 ;
        RECT 588.070 845.720 595.050 846.330 ;
        RECT 595.890 845.720 597.440 846.330 ;
        RECT 5.160 4.280 597.440 845.720 ;
        RECT 5.710 4.000 15.450 4.280 ;
        RECT 16.290 4.000 26.030 4.280 ;
        RECT 26.870 4.000 36.610 4.280 ;
        RECT 37.450 4.000 47.650 4.280 ;
        RECT 48.490 4.000 58.230 4.280 ;
        RECT 59.070 4.000 68.810 4.280 ;
        RECT 69.650 4.000 79.850 4.280 ;
        RECT 80.690 4.000 90.430 4.280 ;
        RECT 91.270 4.000 101.010 4.280 ;
        RECT 101.850 4.000 111.590 4.280 ;
        RECT 112.430 4.000 122.630 4.280 ;
        RECT 123.470 4.000 133.210 4.280 ;
        RECT 134.050 4.000 143.790 4.280 ;
        RECT 144.630 4.000 154.830 4.280 ;
        RECT 155.670 4.000 165.410 4.280 ;
        RECT 166.250 4.000 175.990 4.280 ;
        RECT 176.830 4.000 186.570 4.280 ;
        RECT 187.410 4.000 197.610 4.280 ;
        RECT 198.450 4.000 208.190 4.280 ;
        RECT 209.030 4.000 218.770 4.280 ;
        RECT 219.610 4.000 229.810 4.280 ;
        RECT 230.650 4.000 240.390 4.280 ;
        RECT 241.230 4.000 250.970 4.280 ;
        RECT 251.810 4.000 261.550 4.280 ;
        RECT 262.390 4.000 272.590 4.280 ;
        RECT 273.430 4.000 283.170 4.280 ;
        RECT 284.010 4.000 293.750 4.280 ;
        RECT 294.590 4.000 304.790 4.280 ;
        RECT 305.630 4.000 315.370 4.280 ;
        RECT 316.210 4.000 325.950 4.280 ;
        RECT 326.790 4.000 336.530 4.280 ;
        RECT 337.370 4.000 347.570 4.280 ;
        RECT 348.410 4.000 358.150 4.280 ;
        RECT 358.990 4.000 368.730 4.280 ;
        RECT 369.570 4.000 379.770 4.280 ;
        RECT 380.610 4.000 390.350 4.280 ;
        RECT 391.190 4.000 400.930 4.280 ;
        RECT 401.770 4.000 411.510 4.280 ;
        RECT 412.350 4.000 422.550 4.280 ;
        RECT 423.390 4.000 433.130 4.280 ;
        RECT 433.970 4.000 443.710 4.280 ;
        RECT 444.550 4.000 454.750 4.280 ;
        RECT 455.590 4.000 465.330 4.280 ;
        RECT 466.170 4.000 475.910 4.280 ;
        RECT 476.750 4.000 486.490 4.280 ;
        RECT 487.330 4.000 497.530 4.280 ;
        RECT 498.370 4.000 508.110 4.280 ;
        RECT 508.950 4.000 518.690 4.280 ;
        RECT 519.530 4.000 529.730 4.280 ;
        RECT 530.570 4.000 540.310 4.280 ;
        RECT 541.150 4.000 550.890 4.280 ;
        RECT 551.730 4.000 561.470 4.280 ;
        RECT 562.310 4.000 572.510 4.280 ;
        RECT 573.350 4.000 583.090 4.280 ;
        RECT 583.930 4.000 593.670 4.280 ;
        RECT 594.510 4.000 597.440 4.280 ;
      LAYER met3 ;
        RECT 4.400 844.880 596.000 845.745 ;
        RECT 4.000 838.120 596.000 844.880 ;
        RECT 4.400 836.720 596.000 838.120 ;
        RECT 4.000 829.280 596.000 836.720 ;
        RECT 4.400 827.880 596.000 829.280 ;
        RECT 4.000 821.120 596.000 827.880 ;
        RECT 4.400 819.720 596.000 821.120 ;
        RECT 4.000 812.280 596.000 819.720 ;
        RECT 4.400 810.880 596.000 812.280 ;
        RECT 4.000 804.120 596.000 810.880 ;
        RECT 4.400 802.720 596.000 804.120 ;
        RECT 4.000 795.280 596.000 802.720 ;
        RECT 4.400 793.880 596.000 795.280 ;
        RECT 4.000 787.120 596.000 793.880 ;
        RECT 4.400 785.720 596.000 787.120 ;
        RECT 4.000 779.640 596.000 785.720 ;
        RECT 4.000 778.280 595.600 779.640 ;
        RECT 4.400 778.240 595.600 778.280 ;
        RECT 4.400 776.880 596.000 778.240 ;
        RECT 4.000 770.120 596.000 776.880 ;
        RECT 4.400 768.720 596.000 770.120 ;
        RECT 4.000 761.280 596.000 768.720 ;
        RECT 4.400 759.880 596.000 761.280 ;
        RECT 4.000 753.120 596.000 759.880 ;
        RECT 4.400 751.720 596.000 753.120 ;
        RECT 4.000 744.280 596.000 751.720 ;
        RECT 4.400 742.880 596.000 744.280 ;
        RECT 4.000 736.120 596.000 742.880 ;
        RECT 4.400 734.720 596.000 736.120 ;
        RECT 4.000 727.280 596.000 734.720 ;
        RECT 4.400 725.880 596.000 727.280 ;
        RECT 4.000 719.120 596.000 725.880 ;
        RECT 4.400 717.720 596.000 719.120 ;
        RECT 4.000 710.280 596.000 717.720 ;
        RECT 4.400 708.880 596.000 710.280 ;
        RECT 4.000 702.120 596.000 708.880 ;
        RECT 4.400 700.720 596.000 702.120 ;
        RECT 4.000 693.280 596.000 700.720 ;
        RECT 4.400 691.880 596.000 693.280 ;
        RECT 4.000 685.120 596.000 691.880 ;
        RECT 4.400 683.720 596.000 685.120 ;
        RECT 4.000 676.280 596.000 683.720 ;
        RECT 4.400 674.880 596.000 676.280 ;
        RECT 4.000 668.120 596.000 674.880 ;
        RECT 4.400 666.720 596.000 668.120 ;
        RECT 4.000 659.280 596.000 666.720 ;
        RECT 4.400 657.880 596.000 659.280 ;
        RECT 4.000 651.120 596.000 657.880 ;
        RECT 4.400 649.720 596.000 651.120 ;
        RECT 4.000 642.280 596.000 649.720 ;
        RECT 4.400 640.880 596.000 642.280 ;
        RECT 4.000 638.200 596.000 640.880 ;
        RECT 4.000 636.800 595.600 638.200 ;
        RECT 4.000 634.120 596.000 636.800 ;
        RECT 4.400 632.720 596.000 634.120 ;
        RECT 4.000 625.280 596.000 632.720 ;
        RECT 4.400 623.880 596.000 625.280 ;
        RECT 4.000 617.120 596.000 623.880 ;
        RECT 4.400 615.720 596.000 617.120 ;
        RECT 4.000 608.280 596.000 615.720 ;
        RECT 4.400 606.880 596.000 608.280 ;
        RECT 4.000 600.120 596.000 606.880 ;
        RECT 4.400 598.720 596.000 600.120 ;
        RECT 4.000 591.280 596.000 598.720 ;
        RECT 4.400 589.880 596.000 591.280 ;
        RECT 4.000 583.120 596.000 589.880 ;
        RECT 4.400 581.720 596.000 583.120 ;
        RECT 4.000 574.280 596.000 581.720 ;
        RECT 4.400 572.880 596.000 574.280 ;
        RECT 4.000 566.120 596.000 572.880 ;
        RECT 4.400 564.720 596.000 566.120 ;
        RECT 4.000 557.280 596.000 564.720 ;
        RECT 4.400 555.880 596.000 557.280 ;
        RECT 4.000 549.120 596.000 555.880 ;
        RECT 4.400 547.720 596.000 549.120 ;
        RECT 4.000 540.280 596.000 547.720 ;
        RECT 4.400 538.880 596.000 540.280 ;
        RECT 4.000 532.120 596.000 538.880 ;
        RECT 4.400 530.720 596.000 532.120 ;
        RECT 4.000 523.280 596.000 530.720 ;
        RECT 4.400 521.880 596.000 523.280 ;
        RECT 4.000 515.120 596.000 521.880 ;
        RECT 4.400 513.720 596.000 515.120 ;
        RECT 4.000 506.280 596.000 513.720 ;
        RECT 4.400 504.880 596.000 506.280 ;
        RECT 4.000 498.120 596.000 504.880 ;
        RECT 4.400 496.760 596.000 498.120 ;
        RECT 4.400 496.720 595.600 496.760 ;
        RECT 4.000 495.360 595.600 496.720 ;
        RECT 4.000 489.280 596.000 495.360 ;
        RECT 4.400 487.880 596.000 489.280 ;
        RECT 4.000 481.120 596.000 487.880 ;
        RECT 4.400 479.720 596.000 481.120 ;
        RECT 4.000 472.280 596.000 479.720 ;
        RECT 4.400 470.880 596.000 472.280 ;
        RECT 4.000 464.120 596.000 470.880 ;
        RECT 4.400 462.720 596.000 464.120 ;
        RECT 4.000 455.280 596.000 462.720 ;
        RECT 4.400 453.880 596.000 455.280 ;
        RECT 4.000 447.120 596.000 453.880 ;
        RECT 4.400 445.720 596.000 447.120 ;
        RECT 4.000 438.280 596.000 445.720 ;
        RECT 4.400 436.880 596.000 438.280 ;
        RECT 4.000 430.120 596.000 436.880 ;
        RECT 4.400 428.720 596.000 430.120 ;
        RECT 4.000 421.280 596.000 428.720 ;
        RECT 4.400 419.880 596.000 421.280 ;
        RECT 4.000 413.120 596.000 419.880 ;
        RECT 4.400 411.720 596.000 413.120 ;
        RECT 4.000 404.280 596.000 411.720 ;
        RECT 4.400 402.880 596.000 404.280 ;
        RECT 4.000 396.120 596.000 402.880 ;
        RECT 4.400 394.720 596.000 396.120 ;
        RECT 4.000 387.280 596.000 394.720 ;
        RECT 4.400 385.880 596.000 387.280 ;
        RECT 4.000 379.120 596.000 385.880 ;
        RECT 4.400 377.720 596.000 379.120 ;
        RECT 4.000 370.280 596.000 377.720 ;
        RECT 4.400 368.880 596.000 370.280 ;
        RECT 4.000 362.120 596.000 368.880 ;
        RECT 4.400 360.720 596.000 362.120 ;
        RECT 4.000 354.640 596.000 360.720 ;
        RECT 4.000 353.280 595.600 354.640 ;
        RECT 4.400 353.240 595.600 353.280 ;
        RECT 4.400 351.880 596.000 353.240 ;
        RECT 4.000 345.120 596.000 351.880 ;
        RECT 4.400 343.720 596.000 345.120 ;
        RECT 4.000 336.280 596.000 343.720 ;
        RECT 4.400 334.880 596.000 336.280 ;
        RECT 4.000 328.120 596.000 334.880 ;
        RECT 4.400 326.720 596.000 328.120 ;
        RECT 4.000 319.280 596.000 326.720 ;
        RECT 4.400 317.880 596.000 319.280 ;
        RECT 4.000 311.120 596.000 317.880 ;
        RECT 4.400 309.720 596.000 311.120 ;
        RECT 4.000 302.280 596.000 309.720 ;
        RECT 4.400 300.880 596.000 302.280 ;
        RECT 4.000 294.120 596.000 300.880 ;
        RECT 4.400 292.720 596.000 294.120 ;
        RECT 4.000 285.280 596.000 292.720 ;
        RECT 4.400 283.880 596.000 285.280 ;
        RECT 4.000 277.120 596.000 283.880 ;
        RECT 4.400 275.720 596.000 277.120 ;
        RECT 4.000 268.280 596.000 275.720 ;
        RECT 4.400 266.880 596.000 268.280 ;
        RECT 4.000 260.120 596.000 266.880 ;
        RECT 4.400 258.720 596.000 260.120 ;
        RECT 4.000 251.280 596.000 258.720 ;
        RECT 4.400 249.880 596.000 251.280 ;
        RECT 4.000 243.120 596.000 249.880 ;
        RECT 4.400 241.720 596.000 243.120 ;
        RECT 4.000 234.280 596.000 241.720 ;
        RECT 4.400 232.880 596.000 234.280 ;
        RECT 4.000 226.120 596.000 232.880 ;
        RECT 4.400 224.720 596.000 226.120 ;
        RECT 4.000 217.280 596.000 224.720 ;
        RECT 4.400 215.880 596.000 217.280 ;
        RECT 4.000 213.200 596.000 215.880 ;
        RECT 4.000 211.800 595.600 213.200 ;
        RECT 4.000 209.120 596.000 211.800 ;
        RECT 4.400 207.720 596.000 209.120 ;
        RECT 4.000 200.280 596.000 207.720 ;
        RECT 4.400 198.880 596.000 200.280 ;
        RECT 4.000 192.120 596.000 198.880 ;
        RECT 4.400 190.720 596.000 192.120 ;
        RECT 4.000 183.280 596.000 190.720 ;
        RECT 4.400 181.880 596.000 183.280 ;
        RECT 4.000 175.120 596.000 181.880 ;
        RECT 4.400 173.720 596.000 175.120 ;
        RECT 4.000 166.280 596.000 173.720 ;
        RECT 4.400 164.880 596.000 166.280 ;
        RECT 4.000 158.120 596.000 164.880 ;
        RECT 4.400 156.720 596.000 158.120 ;
        RECT 4.000 149.280 596.000 156.720 ;
        RECT 4.400 147.880 596.000 149.280 ;
        RECT 4.000 141.120 596.000 147.880 ;
        RECT 4.400 139.720 596.000 141.120 ;
        RECT 4.000 132.280 596.000 139.720 ;
        RECT 4.400 130.880 596.000 132.280 ;
        RECT 4.000 124.120 596.000 130.880 ;
        RECT 4.400 122.720 596.000 124.120 ;
        RECT 4.000 115.280 596.000 122.720 ;
        RECT 4.400 113.880 596.000 115.280 ;
        RECT 4.000 107.120 596.000 113.880 ;
        RECT 4.400 105.720 596.000 107.120 ;
        RECT 4.000 98.280 596.000 105.720 ;
        RECT 4.400 96.880 596.000 98.280 ;
        RECT 4.000 90.120 596.000 96.880 ;
        RECT 4.400 88.720 596.000 90.120 ;
        RECT 4.000 81.280 596.000 88.720 ;
        RECT 4.400 79.880 596.000 81.280 ;
        RECT 4.000 73.120 596.000 79.880 ;
        RECT 4.400 71.760 596.000 73.120 ;
        RECT 4.400 71.720 595.600 71.760 ;
        RECT 4.000 70.360 595.600 71.720 ;
        RECT 4.000 64.280 596.000 70.360 ;
        RECT 4.400 62.880 596.000 64.280 ;
        RECT 4.000 56.120 596.000 62.880 ;
        RECT 4.400 54.720 596.000 56.120 ;
        RECT 4.000 47.280 596.000 54.720 ;
        RECT 4.400 45.880 596.000 47.280 ;
        RECT 4.000 39.120 596.000 45.880 ;
        RECT 4.400 37.720 596.000 39.120 ;
        RECT 4.000 30.280 596.000 37.720 ;
        RECT 4.400 28.880 596.000 30.280 ;
        RECT 4.000 22.120 596.000 28.880 ;
        RECT 4.400 20.720 596.000 22.120 ;
        RECT 4.000 13.280 596.000 20.720 ;
        RECT 4.400 11.880 596.000 13.280 ;
        RECT 4.000 5.120 596.000 11.880 ;
        RECT 4.400 4.255 596.000 5.120 ;
      LAYER met4 ;
        RECT 46.295 12.415 97.440 835.545 ;
        RECT 99.840 12.415 174.240 835.545 ;
        RECT 176.640 12.415 251.040 835.545 ;
        RECT 253.440 12.415 327.840 835.545 ;
        RECT 330.240 12.415 404.640 835.545 ;
        RECT 407.040 12.415 481.440 835.545 ;
        RECT 483.840 12.415 558.240 835.545 ;
        RECT 560.640 12.415 573.785 835.545 ;
  END
END Peripherals
END LIBRARY

