magic
tech sky130A
magscale 1 2
timestamp 1653087023
<< obsli1 >>
rect 1104 2159 118864 137649
<< obsm1 >>
rect 1026 1640 119126 137680
<< metal2 >>
rect 754 139200 810 140000
rect 2318 139200 2374 140000
rect 3882 139200 3938 140000
rect 5446 139200 5502 140000
rect 7010 139200 7066 140000
rect 8574 139200 8630 140000
rect 10138 139200 10194 140000
rect 11794 139200 11850 140000
rect 13358 139200 13414 140000
rect 14922 139200 14978 140000
rect 16486 139200 16542 140000
rect 18050 139200 18106 140000
rect 19614 139200 19670 140000
rect 21270 139200 21326 140000
rect 22834 139200 22890 140000
rect 24398 139200 24454 140000
rect 25962 139200 26018 140000
rect 27526 139200 27582 140000
rect 29090 139200 29146 140000
rect 30746 139200 30802 140000
rect 32310 139200 32366 140000
rect 33874 139200 33930 140000
rect 35438 139200 35494 140000
rect 37002 139200 37058 140000
rect 38566 139200 38622 140000
rect 40130 139200 40186 140000
rect 41786 139200 41842 140000
rect 43350 139200 43406 140000
rect 44914 139200 44970 140000
rect 46478 139200 46534 140000
rect 48042 139200 48098 140000
rect 49606 139200 49662 140000
rect 51262 139200 51318 140000
rect 52826 139200 52882 140000
rect 54390 139200 54446 140000
rect 55954 139200 56010 140000
rect 57518 139200 57574 140000
rect 59082 139200 59138 140000
rect 60738 139200 60794 140000
rect 62302 139200 62358 140000
rect 63866 139200 63922 140000
rect 65430 139200 65486 140000
rect 66994 139200 67050 140000
rect 68558 139200 68614 140000
rect 70122 139200 70178 140000
rect 71778 139200 71834 140000
rect 73342 139200 73398 140000
rect 74906 139200 74962 140000
rect 76470 139200 76526 140000
rect 78034 139200 78090 140000
rect 79598 139200 79654 140000
rect 81254 139200 81310 140000
rect 82818 139200 82874 140000
rect 84382 139200 84438 140000
rect 85946 139200 86002 140000
rect 87510 139200 87566 140000
rect 89074 139200 89130 140000
rect 90730 139200 90786 140000
rect 92294 139200 92350 140000
rect 93858 139200 93914 140000
rect 95422 139200 95478 140000
rect 96986 139200 97042 140000
rect 98550 139200 98606 140000
rect 100114 139200 100170 140000
rect 101770 139200 101826 140000
rect 103334 139200 103390 140000
rect 104898 139200 104954 140000
rect 106462 139200 106518 140000
rect 108026 139200 108082 140000
rect 109590 139200 109646 140000
rect 111246 139200 111302 140000
rect 112810 139200 112866 140000
rect 114374 139200 114430 140000
rect 115938 139200 115994 140000
rect 117502 139200 117558 140000
rect 119066 139200 119122 140000
rect 1030 0 1086 800
rect 3146 0 3202 800
rect 5262 0 5318 800
rect 7378 0 7434 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 16026 0 16082 800
rect 18142 0 18198 800
rect 20258 0 20314 800
rect 22374 0 22430 800
rect 24582 0 24638 800
rect 26698 0 26754 800
rect 28814 0 28870 800
rect 31022 0 31078 800
rect 33138 0 33194 800
rect 35254 0 35310 800
rect 37370 0 37426 800
rect 39578 0 39634 800
rect 41694 0 41750 800
rect 43810 0 43866 800
rect 46018 0 46074 800
rect 48134 0 48190 800
rect 50250 0 50306 800
rect 52366 0 52422 800
rect 54574 0 54630 800
rect 56690 0 56746 800
rect 58806 0 58862 800
rect 61014 0 61070 800
rect 63130 0 63186 800
rect 65246 0 65302 800
rect 67362 0 67418 800
rect 69570 0 69626 800
rect 71686 0 71742 800
rect 73802 0 73858 800
rect 76010 0 76066 800
rect 78126 0 78182 800
rect 80242 0 80298 800
rect 82358 0 82414 800
rect 84566 0 84622 800
rect 86682 0 86738 800
rect 88798 0 88854 800
rect 91006 0 91062 800
rect 93122 0 93178 800
rect 95238 0 95294 800
rect 97354 0 97410 800
rect 99562 0 99618 800
rect 101678 0 101734 800
rect 103794 0 103850 800
rect 106002 0 106058 800
rect 108118 0 108174 800
rect 110234 0 110290 800
rect 112350 0 112406 800
rect 114558 0 114614 800
rect 116674 0 116730 800
rect 118790 0 118846 800
<< obsm2 >>
rect 1032 139144 2262 139346
rect 2430 139144 3826 139346
rect 3994 139144 5390 139346
rect 5558 139144 6954 139346
rect 7122 139144 8518 139346
rect 8686 139144 10082 139346
rect 10250 139144 11738 139346
rect 11906 139144 13302 139346
rect 13470 139144 14866 139346
rect 15034 139144 16430 139346
rect 16598 139144 17994 139346
rect 18162 139144 19558 139346
rect 19726 139144 21214 139346
rect 21382 139144 22778 139346
rect 22946 139144 24342 139346
rect 24510 139144 25906 139346
rect 26074 139144 27470 139346
rect 27638 139144 29034 139346
rect 29202 139144 30690 139346
rect 30858 139144 32254 139346
rect 32422 139144 33818 139346
rect 33986 139144 35382 139346
rect 35550 139144 36946 139346
rect 37114 139144 38510 139346
rect 38678 139144 40074 139346
rect 40242 139144 41730 139346
rect 41898 139144 43294 139346
rect 43462 139144 44858 139346
rect 45026 139144 46422 139346
rect 46590 139144 47986 139346
rect 48154 139144 49550 139346
rect 49718 139144 51206 139346
rect 51374 139144 52770 139346
rect 52938 139144 54334 139346
rect 54502 139144 55898 139346
rect 56066 139144 57462 139346
rect 57630 139144 59026 139346
rect 59194 139144 60682 139346
rect 60850 139144 62246 139346
rect 62414 139144 63810 139346
rect 63978 139144 65374 139346
rect 65542 139144 66938 139346
rect 67106 139144 68502 139346
rect 68670 139144 70066 139346
rect 70234 139144 71722 139346
rect 71890 139144 73286 139346
rect 73454 139144 74850 139346
rect 75018 139144 76414 139346
rect 76582 139144 77978 139346
rect 78146 139144 79542 139346
rect 79710 139144 81198 139346
rect 81366 139144 82762 139346
rect 82930 139144 84326 139346
rect 84494 139144 85890 139346
rect 86058 139144 87454 139346
rect 87622 139144 89018 139346
rect 89186 139144 90674 139346
rect 90842 139144 92238 139346
rect 92406 139144 93802 139346
rect 93970 139144 95366 139346
rect 95534 139144 96930 139346
rect 97098 139144 98494 139346
rect 98662 139144 100058 139346
rect 100226 139144 101714 139346
rect 101882 139144 103278 139346
rect 103446 139144 104842 139346
rect 105010 139144 106406 139346
rect 106574 139144 107970 139346
rect 108138 139144 109534 139346
rect 109702 139144 111190 139346
rect 111358 139144 112754 139346
rect 112922 139144 114318 139346
rect 114486 139144 115882 139346
rect 116050 139144 117446 139346
rect 117614 139144 119010 139346
rect 1032 856 119120 139144
rect 1142 711 3090 856
rect 3258 711 5206 856
rect 5374 711 7322 856
rect 7490 711 9530 856
rect 9698 711 11646 856
rect 11814 711 13762 856
rect 13930 711 15970 856
rect 16138 711 18086 856
rect 18254 711 20202 856
rect 20370 711 22318 856
rect 22486 711 24526 856
rect 24694 711 26642 856
rect 26810 711 28758 856
rect 28926 711 30966 856
rect 31134 711 33082 856
rect 33250 711 35198 856
rect 35366 711 37314 856
rect 37482 711 39522 856
rect 39690 711 41638 856
rect 41806 711 43754 856
rect 43922 711 45962 856
rect 46130 711 48078 856
rect 48246 711 50194 856
rect 50362 711 52310 856
rect 52478 711 54518 856
rect 54686 711 56634 856
rect 56802 711 58750 856
rect 58918 711 60958 856
rect 61126 711 63074 856
rect 63242 711 65190 856
rect 65358 711 67306 856
rect 67474 711 69514 856
rect 69682 711 71630 856
rect 71798 711 73746 856
rect 73914 711 75954 856
rect 76122 711 78070 856
rect 78238 711 80186 856
rect 80354 711 82302 856
rect 82470 711 84510 856
rect 84678 711 86626 856
rect 86794 711 88742 856
rect 88910 711 90950 856
rect 91118 711 93066 856
rect 93234 711 95182 856
rect 95350 711 97298 856
rect 97466 711 99506 856
rect 99674 711 101622 856
rect 101790 711 103738 856
rect 103906 711 105946 856
rect 106114 711 108062 856
rect 108230 711 110178 856
rect 110346 711 112294 856
rect 112462 711 114502 856
rect 114670 711 116618 856
rect 116786 711 118734 856
rect 118902 711 119120 856
<< metal3 >>
rect 0 139136 800 139256
rect 0 137776 800 137896
rect 0 136416 800 136536
rect 0 134920 800 135040
rect 0 133560 800 133680
rect 0 132200 800 132320
rect 0 130704 800 130824
rect 0 129344 800 129464
rect 0 127984 800 128104
rect 119200 128120 120000 128240
rect 0 126624 800 126744
rect 0 125128 800 125248
rect 0 123768 800 123888
rect 0 122408 800 122528
rect 0 120912 800 121032
rect 0 119552 800 119672
rect 0 118192 800 118312
rect 0 116832 800 116952
rect 0 115336 800 115456
rect 0 113976 800 114096
rect 0 112616 800 112736
rect 0 111120 800 111240
rect 0 109760 800 109880
rect 0 108400 800 108520
rect 0 107040 800 107160
rect 0 105544 800 105664
rect 119200 104864 120000 104984
rect 0 104184 800 104304
rect 0 102824 800 102944
rect 0 101328 800 101448
rect 0 99968 800 100088
rect 0 98608 800 98728
rect 0 97248 800 97368
rect 0 95752 800 95872
rect 0 94392 800 94512
rect 0 93032 800 93152
rect 0 91536 800 91656
rect 0 90176 800 90296
rect 0 88816 800 88936
rect 0 87320 800 87440
rect 0 85960 800 86080
rect 0 84600 800 84720
rect 0 83240 800 83360
rect 0 81744 800 81864
rect 119200 81472 120000 81592
rect 0 80384 800 80504
rect 0 79024 800 79144
rect 0 77528 800 77648
rect 0 76168 800 76288
rect 0 74808 800 74928
rect 0 73448 800 73568
rect 0 71952 800 72072
rect 0 70592 800 70712
rect 0 69232 800 69352
rect 0 67736 800 67856
rect 0 66376 800 66496
rect 0 65016 800 65136
rect 0 63656 800 63776
rect 0 62160 800 62280
rect 0 60800 800 60920
rect 0 59440 800 59560
rect 119200 58216 120000 58336
rect 0 57944 800 58064
rect 0 56584 800 56704
rect 0 55224 800 55344
rect 0 53864 800 53984
rect 0 52368 800 52488
rect 0 51008 800 51128
rect 0 49648 800 49768
rect 0 48152 800 48272
rect 0 46792 800 46912
rect 0 45432 800 45552
rect 0 43936 800 44056
rect 0 42576 800 42696
rect 0 41216 800 41336
rect 0 39856 800 39976
rect 0 38360 800 38480
rect 0 37000 800 37120
rect 0 35640 800 35760
rect 119200 34824 120000 34944
rect 0 34144 800 34264
rect 0 32784 800 32904
rect 0 31424 800 31544
rect 0 30064 800 30184
rect 0 28568 800 28688
rect 0 27208 800 27328
rect 0 25848 800 25968
rect 0 24352 800 24472
rect 0 22992 800 23112
rect 0 21632 800 21752
rect 0 20272 800 20392
rect 0 18776 800 18896
rect 0 17416 800 17536
rect 0 16056 800 16176
rect 0 14560 800 14680
rect 0 13200 800 13320
rect 0 11840 800 11960
rect 119200 11568 120000 11688
rect 0 10480 800 10600
rect 0 8984 800 9104
rect 0 7624 800 7744
rect 0 6264 800 6384
rect 0 4768 800 4888
rect 0 3408 800 3528
rect 0 2048 800 2168
rect 0 688 800 808
<< obsm3 >>
rect 880 139056 119200 139229
rect 800 137976 119200 139056
rect 880 137696 119200 137976
rect 800 136616 119200 137696
rect 880 136336 119200 136616
rect 800 135120 119200 136336
rect 880 134840 119200 135120
rect 800 133760 119200 134840
rect 880 133480 119200 133760
rect 800 132400 119200 133480
rect 880 132120 119200 132400
rect 800 130904 119200 132120
rect 880 130624 119200 130904
rect 800 129544 119200 130624
rect 880 129264 119200 129544
rect 800 128320 119200 129264
rect 800 128184 119120 128320
rect 880 128040 119120 128184
rect 880 127904 119200 128040
rect 800 126824 119200 127904
rect 880 126544 119200 126824
rect 800 125328 119200 126544
rect 880 125048 119200 125328
rect 800 123968 119200 125048
rect 880 123688 119200 123968
rect 800 122608 119200 123688
rect 880 122328 119200 122608
rect 800 121112 119200 122328
rect 880 120832 119200 121112
rect 800 119752 119200 120832
rect 880 119472 119200 119752
rect 800 118392 119200 119472
rect 880 118112 119200 118392
rect 800 117032 119200 118112
rect 880 116752 119200 117032
rect 800 115536 119200 116752
rect 880 115256 119200 115536
rect 800 114176 119200 115256
rect 880 113896 119200 114176
rect 800 112816 119200 113896
rect 880 112536 119200 112816
rect 800 111320 119200 112536
rect 880 111040 119200 111320
rect 800 109960 119200 111040
rect 880 109680 119200 109960
rect 800 108600 119200 109680
rect 880 108320 119200 108600
rect 800 107240 119200 108320
rect 880 106960 119200 107240
rect 800 105744 119200 106960
rect 880 105464 119200 105744
rect 800 105064 119200 105464
rect 800 104784 119120 105064
rect 800 104384 119200 104784
rect 880 104104 119200 104384
rect 800 103024 119200 104104
rect 880 102744 119200 103024
rect 800 101528 119200 102744
rect 880 101248 119200 101528
rect 800 100168 119200 101248
rect 880 99888 119200 100168
rect 800 98808 119200 99888
rect 880 98528 119200 98808
rect 800 97448 119200 98528
rect 880 97168 119200 97448
rect 800 95952 119200 97168
rect 880 95672 119200 95952
rect 800 94592 119200 95672
rect 880 94312 119200 94592
rect 800 93232 119200 94312
rect 880 92952 119200 93232
rect 800 91736 119200 92952
rect 880 91456 119200 91736
rect 800 90376 119200 91456
rect 880 90096 119200 90376
rect 800 89016 119200 90096
rect 880 88736 119200 89016
rect 800 87520 119200 88736
rect 880 87240 119200 87520
rect 800 86160 119200 87240
rect 880 85880 119200 86160
rect 800 84800 119200 85880
rect 880 84520 119200 84800
rect 800 83440 119200 84520
rect 880 83160 119200 83440
rect 800 81944 119200 83160
rect 880 81672 119200 81944
rect 880 81664 119120 81672
rect 800 81392 119120 81664
rect 800 80584 119200 81392
rect 880 80304 119200 80584
rect 800 79224 119200 80304
rect 880 78944 119200 79224
rect 800 77728 119200 78944
rect 880 77448 119200 77728
rect 800 76368 119200 77448
rect 880 76088 119200 76368
rect 800 75008 119200 76088
rect 880 74728 119200 75008
rect 800 73648 119200 74728
rect 880 73368 119200 73648
rect 800 72152 119200 73368
rect 880 71872 119200 72152
rect 800 70792 119200 71872
rect 880 70512 119200 70792
rect 800 69432 119200 70512
rect 880 69152 119200 69432
rect 800 67936 119200 69152
rect 880 67656 119200 67936
rect 800 66576 119200 67656
rect 880 66296 119200 66576
rect 800 65216 119200 66296
rect 880 64936 119200 65216
rect 800 63856 119200 64936
rect 880 63576 119200 63856
rect 800 62360 119200 63576
rect 880 62080 119200 62360
rect 800 61000 119200 62080
rect 880 60720 119200 61000
rect 800 59640 119200 60720
rect 880 59360 119200 59640
rect 800 58416 119200 59360
rect 800 58144 119120 58416
rect 880 58136 119120 58144
rect 880 57864 119200 58136
rect 800 56784 119200 57864
rect 880 56504 119200 56784
rect 800 55424 119200 56504
rect 880 55144 119200 55424
rect 800 54064 119200 55144
rect 880 53784 119200 54064
rect 800 52568 119200 53784
rect 880 52288 119200 52568
rect 800 51208 119200 52288
rect 880 50928 119200 51208
rect 800 49848 119200 50928
rect 880 49568 119200 49848
rect 800 48352 119200 49568
rect 880 48072 119200 48352
rect 800 46992 119200 48072
rect 880 46712 119200 46992
rect 800 45632 119200 46712
rect 880 45352 119200 45632
rect 800 44136 119200 45352
rect 880 43856 119200 44136
rect 800 42776 119200 43856
rect 880 42496 119200 42776
rect 800 41416 119200 42496
rect 880 41136 119200 41416
rect 800 40056 119200 41136
rect 880 39776 119200 40056
rect 800 38560 119200 39776
rect 880 38280 119200 38560
rect 800 37200 119200 38280
rect 880 36920 119200 37200
rect 800 35840 119200 36920
rect 880 35560 119200 35840
rect 800 35024 119200 35560
rect 800 34744 119120 35024
rect 800 34344 119200 34744
rect 880 34064 119200 34344
rect 800 32984 119200 34064
rect 880 32704 119200 32984
rect 800 31624 119200 32704
rect 880 31344 119200 31624
rect 800 30264 119200 31344
rect 880 29984 119200 30264
rect 800 28768 119200 29984
rect 880 28488 119200 28768
rect 800 27408 119200 28488
rect 880 27128 119200 27408
rect 800 26048 119200 27128
rect 880 25768 119200 26048
rect 800 24552 119200 25768
rect 880 24272 119200 24552
rect 800 23192 119200 24272
rect 880 22912 119200 23192
rect 800 21832 119200 22912
rect 880 21552 119200 21832
rect 800 20472 119200 21552
rect 880 20192 119200 20472
rect 800 18976 119200 20192
rect 880 18696 119200 18976
rect 800 17616 119200 18696
rect 880 17336 119200 17616
rect 800 16256 119200 17336
rect 880 15976 119200 16256
rect 800 14760 119200 15976
rect 880 14480 119200 14760
rect 800 13400 119200 14480
rect 880 13120 119200 13400
rect 800 12040 119200 13120
rect 880 11768 119200 12040
rect 880 11760 119120 11768
rect 800 11488 119120 11760
rect 800 10680 119200 11488
rect 880 10400 119200 10680
rect 800 9184 119200 10400
rect 880 8904 119200 9184
rect 800 7824 119200 8904
rect 880 7544 119200 7824
rect 800 6464 119200 7544
rect 880 6184 119200 6464
rect 800 4968 119200 6184
rect 880 4688 119200 4968
rect 800 3608 119200 4688
rect 880 3328 119200 3608
rect 800 2248 119200 3328
rect 880 1968 119200 2248
rect 800 888 119200 1968
rect 880 715 119200 888
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
<< obsm4 >>
rect 4659 19891 19488 137053
rect 19968 19891 34848 137053
rect 35328 19891 50208 137053
rect 50688 19891 65568 137053
rect 66048 19891 80928 137053
rect 81408 19891 88813 137053
<< labels >>
rlabel metal2 s 86682 0 86738 800 6 flash_csb
port 1 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 flash_io0_read
port 2 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 flash_io0_we
port 3 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 flash_io0_write
port 4 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 flash_io1_read
port 5 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 flash_io1_we
port 6 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 flash_io1_write
port 7 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 flash_sck
port 8 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 internal_uart_rx
port 9 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 internal_uart_tx
port 10 nsew signal output
rlabel metal2 s 754 139200 810 140000 6 io_in[0]
port 11 nsew signal input
rlabel metal2 s 16486 139200 16542 140000 6 io_in[10]
port 12 nsew signal input
rlabel metal2 s 18050 139200 18106 140000 6 io_in[11]
port 13 nsew signal input
rlabel metal2 s 19614 139200 19670 140000 6 io_in[12]
port 14 nsew signal input
rlabel metal2 s 21270 139200 21326 140000 6 io_in[13]
port 15 nsew signal input
rlabel metal2 s 22834 139200 22890 140000 6 io_in[14]
port 16 nsew signal input
rlabel metal2 s 24398 139200 24454 140000 6 io_in[15]
port 17 nsew signal input
rlabel metal2 s 25962 139200 26018 140000 6 io_in[16]
port 18 nsew signal input
rlabel metal2 s 27526 139200 27582 140000 6 io_in[17]
port 19 nsew signal input
rlabel metal2 s 29090 139200 29146 140000 6 io_in[18]
port 20 nsew signal input
rlabel metal2 s 30746 139200 30802 140000 6 io_in[19]
port 21 nsew signal input
rlabel metal2 s 2318 139200 2374 140000 6 io_in[1]
port 22 nsew signal input
rlabel metal2 s 32310 139200 32366 140000 6 io_in[20]
port 23 nsew signal input
rlabel metal2 s 33874 139200 33930 140000 6 io_in[21]
port 24 nsew signal input
rlabel metal2 s 35438 139200 35494 140000 6 io_in[22]
port 25 nsew signal input
rlabel metal2 s 37002 139200 37058 140000 6 io_in[23]
port 26 nsew signal input
rlabel metal2 s 38566 139200 38622 140000 6 io_in[24]
port 27 nsew signal input
rlabel metal2 s 40130 139200 40186 140000 6 io_in[25]
port 28 nsew signal input
rlabel metal2 s 41786 139200 41842 140000 6 io_in[26]
port 29 nsew signal input
rlabel metal2 s 43350 139200 43406 140000 6 io_in[27]
port 30 nsew signal input
rlabel metal2 s 44914 139200 44970 140000 6 io_in[28]
port 31 nsew signal input
rlabel metal2 s 46478 139200 46534 140000 6 io_in[29]
port 32 nsew signal input
rlabel metal2 s 3882 139200 3938 140000 6 io_in[2]
port 33 nsew signal input
rlabel metal2 s 48042 139200 48098 140000 6 io_in[30]
port 34 nsew signal input
rlabel metal2 s 49606 139200 49662 140000 6 io_in[31]
port 35 nsew signal input
rlabel metal2 s 51262 139200 51318 140000 6 io_in[32]
port 36 nsew signal input
rlabel metal2 s 52826 139200 52882 140000 6 io_in[33]
port 37 nsew signal input
rlabel metal2 s 54390 139200 54446 140000 6 io_in[34]
port 38 nsew signal input
rlabel metal2 s 55954 139200 56010 140000 6 io_in[35]
port 39 nsew signal input
rlabel metal2 s 57518 139200 57574 140000 6 io_in[36]
port 40 nsew signal input
rlabel metal2 s 59082 139200 59138 140000 6 io_in[37]
port 41 nsew signal input
rlabel metal2 s 5446 139200 5502 140000 6 io_in[3]
port 42 nsew signal input
rlabel metal2 s 7010 139200 7066 140000 6 io_in[4]
port 43 nsew signal input
rlabel metal2 s 8574 139200 8630 140000 6 io_in[5]
port 44 nsew signal input
rlabel metal2 s 10138 139200 10194 140000 6 io_in[6]
port 45 nsew signal input
rlabel metal2 s 11794 139200 11850 140000 6 io_in[7]
port 46 nsew signal input
rlabel metal2 s 13358 139200 13414 140000 6 io_in[8]
port 47 nsew signal input
rlabel metal2 s 14922 139200 14978 140000 6 io_in[9]
port 48 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 io_oeb[0]
port 49 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 io_oeb[10]
port 50 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 io_oeb[11]
port 51 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 io_oeb[12]
port 52 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 io_oeb[13]
port 53 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 io_oeb[14]
port 54 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 io_oeb[15]
port 55 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 io_oeb[16]
port 56 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 io_oeb[17]
port 57 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 io_oeb[18]
port 58 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 io_oeb[19]
port 59 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 io_oeb[1]
port 60 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 io_oeb[20]
port 61 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 io_oeb[21]
port 62 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 io_oeb[22]
port 63 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 io_oeb[23]
port 64 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 io_oeb[24]
port 65 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 io_oeb[25]
port 66 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 io_oeb[26]
port 67 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 io_oeb[27]
port 68 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 io_oeb[28]
port 69 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 io_oeb[29]
port 70 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 io_oeb[2]
port 71 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 io_oeb[30]
port 72 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 io_oeb[31]
port 73 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 io_oeb[32]
port 74 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 io_oeb[33]
port 75 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 io_oeb[34]
port 76 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 io_oeb[35]
port 77 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 io_oeb[36]
port 78 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 io_oeb[37]
port 79 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 io_oeb[3]
port 80 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 io_oeb[4]
port 81 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 io_oeb[5]
port 82 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 io_oeb[6]
port 83 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 io_oeb[7]
port 84 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 io_oeb[8]
port 85 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 60738 139200 60794 140000 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 76470 139200 76526 140000 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 78034 139200 78090 140000 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 79598 139200 79654 140000 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 81254 139200 81310 140000 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 82818 139200 82874 140000 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 84382 139200 84438 140000 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 85946 139200 86002 140000 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 87510 139200 87566 140000 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 89074 139200 89130 140000 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 90730 139200 90786 140000 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 62302 139200 62358 140000 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 92294 139200 92350 140000 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 93858 139200 93914 140000 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 95422 139200 95478 140000 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 96986 139200 97042 140000 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 98550 139200 98606 140000 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 100114 139200 100170 140000 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 101770 139200 101826 140000 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 103334 139200 103390 140000 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 104898 139200 104954 140000 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 106462 139200 106518 140000 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 63866 139200 63922 140000 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 108026 139200 108082 140000 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 109590 139200 109646 140000 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 111246 139200 111302 140000 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 112810 139200 112866 140000 6 io_out[33]
port 113 nsew signal output
rlabel metal2 s 114374 139200 114430 140000 6 io_out[34]
port 114 nsew signal output
rlabel metal2 s 115938 139200 115994 140000 6 io_out[35]
port 115 nsew signal output
rlabel metal2 s 117502 139200 117558 140000 6 io_out[36]
port 116 nsew signal output
rlabel metal2 s 119066 139200 119122 140000 6 io_out[37]
port 117 nsew signal output
rlabel metal2 s 65430 139200 65486 140000 6 io_out[3]
port 118 nsew signal output
rlabel metal2 s 66994 139200 67050 140000 6 io_out[4]
port 119 nsew signal output
rlabel metal2 s 68558 139200 68614 140000 6 io_out[5]
port 120 nsew signal output
rlabel metal2 s 70122 139200 70178 140000 6 io_out[6]
port 121 nsew signal output
rlabel metal2 s 71778 139200 71834 140000 6 io_out[7]
port 122 nsew signal output
rlabel metal2 s 73342 139200 73398 140000 6 io_out[8]
port 123 nsew signal output
rlabel metal2 s 74906 139200 74962 140000 6 io_out[9]
port 124 nsew signal output
rlabel metal3 s 119200 58216 120000 58336 6 jtag_tck
port 125 nsew signal output
rlabel metal3 s 119200 81472 120000 81592 6 jtag_tdi
port 126 nsew signal output
rlabel metal3 s 119200 104864 120000 104984 6 jtag_tdo
port 127 nsew signal input
rlabel metal3 s 119200 128120 120000 128240 6 jtag_tms
port 128 nsew signal output
rlabel metal3 s 119200 11568 120000 11688 6 probe_blink[0]
port 129 nsew signal output
rlabel metal3 s 119200 34824 120000 34944 6 probe_blink[1]
port 130 nsew signal output
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal2 s 108118 0 108174 800 6 vga_b[0]
port 132 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 vga_b[1]
port 133 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 vga_g[0]
port 134 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 vga_g[1]
port 135 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 vga_hsync
port 136 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 vga_r[0]
port 137 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 vga_r[1]
port 138 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 vga_vsync
port 139 nsew signal input
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal3 s 0 688 800 808 6 wb_ack_o
port 141 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 wb_adr_i[0]
port 142 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 wb_adr_i[10]
port 143 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 wb_adr_i[11]
port 144 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 wb_adr_i[12]
port 145 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 wb_adr_i[13]
port 146 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 wb_adr_i[14]
port 147 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 wb_adr_i[15]
port 148 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 wb_adr_i[16]
port 149 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 wb_adr_i[17]
port 150 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 wb_adr_i[18]
port 151 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 wb_adr_i[19]
port 152 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 wb_adr_i[1]
port 153 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 wb_adr_i[20]
port 154 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 wb_adr_i[21]
port 155 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 wb_adr_i[22]
port 156 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 wb_adr_i[23]
port 157 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 wb_adr_i[2]
port 158 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 wb_adr_i[3]
port 159 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wb_adr_i[4]
port 160 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 wb_adr_i[5]
port 161 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 wb_adr_i[6]
port 162 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 wb_adr_i[7]
port 163 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 wb_adr_i[8]
port 164 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 wb_adr_i[9]
port 165 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 wb_clk_i
port 166 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 wb_cyc_i
port 167 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 wb_data_i[0]
port 168 nsew signal input
rlabel metal3 s 0 60800 800 60920 6 wb_data_i[10]
port 169 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 wb_data_i[11]
port 170 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 wb_data_i[12]
port 171 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 wb_data_i[13]
port 172 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wb_data_i[14]
port 173 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 wb_data_i[15]
port 174 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 wb_data_i[16]
port 175 nsew signal input
rlabel metal3 s 0 90176 800 90296 6 wb_data_i[17]
port 176 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 wb_data_i[18]
port 177 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 wb_data_i[19]
port 178 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 wb_data_i[1]
port 179 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 wb_data_i[20]
port 180 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 wb_data_i[21]
port 181 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 wb_data_i[22]
port 182 nsew signal input
rlabel metal3 s 0 115336 800 115456 6 wb_data_i[23]
port 183 nsew signal input
rlabel metal3 s 0 118192 800 118312 6 wb_data_i[24]
port 184 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 wb_data_i[25]
port 185 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 wb_data_i[26]
port 186 nsew signal input
rlabel metal3 s 0 126624 800 126744 6 wb_data_i[27]
port 187 nsew signal input
rlabel metal3 s 0 129344 800 129464 6 wb_data_i[28]
port 188 nsew signal input
rlabel metal3 s 0 132200 800 132320 6 wb_data_i[29]
port 189 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 wb_data_i[2]
port 190 nsew signal input
rlabel metal3 s 0 134920 800 135040 6 wb_data_i[30]
port 191 nsew signal input
rlabel metal3 s 0 137776 800 137896 6 wb_data_i[31]
port 192 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 wb_data_i[3]
port 193 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 wb_data_i[4]
port 194 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 wb_data_i[5]
port 195 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 wb_data_i[6]
port 196 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 wb_data_i[7]
port 197 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 wb_data_i[8]
port 198 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 wb_data_i[9]
port 199 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 wb_data_o[0]
port 200 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 wb_data_o[10]
port 201 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 wb_data_o[11]
port 202 nsew signal output
rlabel metal3 s 0 70592 800 70712 6 wb_data_o[12]
port 203 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 wb_data_o[13]
port 204 nsew signal output
rlabel metal3 s 0 79024 800 79144 6 wb_data_o[14]
port 205 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 wb_data_o[15]
port 206 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 wb_data_o[16]
port 207 nsew signal output
rlabel metal3 s 0 91536 800 91656 6 wb_data_o[17]
port 208 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 wb_data_o[18]
port 209 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 wb_data_o[19]
port 210 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 wb_data_o[1]
port 211 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 wb_data_o[20]
port 212 nsew signal output
rlabel metal3 s 0 108400 800 108520 6 wb_data_o[21]
port 213 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 wb_data_o[22]
port 214 nsew signal output
rlabel metal3 s 0 116832 800 116952 6 wb_data_o[23]
port 215 nsew signal output
rlabel metal3 s 0 119552 800 119672 6 wb_data_o[24]
port 216 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 wb_data_o[25]
port 217 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 wb_data_o[26]
port 218 nsew signal output
rlabel metal3 s 0 127984 800 128104 6 wb_data_o[27]
port 219 nsew signal output
rlabel metal3 s 0 130704 800 130824 6 wb_data_o[28]
port 220 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 wb_data_o[29]
port 221 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 wb_data_o[2]
port 222 nsew signal output
rlabel metal3 s 0 136416 800 136536 6 wb_data_o[30]
port 223 nsew signal output
rlabel metal3 s 0 139136 800 139256 6 wb_data_o[31]
port 224 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 wb_data_o[3]
port 225 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 wb_data_o[4]
port 226 nsew signal output
rlabel metal3 s 0 41216 800 41336 6 wb_data_o[5]
port 227 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 wb_data_o[6]
port 228 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 wb_data_o[7]
port 229 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 wb_data_o[8]
port 230 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 wb_data_o[9]
port 231 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 wb_error_o
port 232 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 wb_rst_i
port 233 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 wb_sel_i[0]
port 234 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 wb_sel_i[1]
port 235 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 wb_sel_i[2]
port 236 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 wb_sel_i[3]
port 237 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 wb_stall_o
port 238 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 wb_stb_i
port 239 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 wb_we_i
port 240 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29559574
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripherals_Flat/runs/Peripherals_Flat/results/signoff/Peripherals.magic.gds
string GDS_START 1002462
<< end >>

