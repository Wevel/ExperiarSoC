magic
tech sky130A
magscale 1 2
timestamp 1652654225
<< nwell >>
rect 1066 22021 8870 22342
rect 1066 20933 8870 21499
rect 1066 19845 8870 20411
rect 1066 18757 8870 19323
rect 1066 17669 8870 18235
rect 1066 16581 8870 17147
rect 1066 15493 8870 16059
rect 1066 14405 8870 14971
rect 1066 13317 8870 13883
rect 1066 12229 8870 12795
rect 1066 11141 8870 11707
rect 1066 10053 8870 10619
rect 1066 8965 8870 9531
rect 1066 7877 8870 8443
rect 1066 6789 8870 7355
rect 1066 5701 8870 6267
rect 1066 4613 8870 5179
rect 1066 3525 8870 4091
rect 1066 2437 8870 3003
<< obsli1 >>
rect 1104 2159 8832 22321
<< obsm1 >>
rect 1104 2128 8832 22352
<< metal2 >>
rect 4986 0 5042 800
<< obsm2 >>
rect 2248 856 8262 24721
rect 2248 167 4930 856
rect 5098 167 8262 856
<< metal3 >>
rect 9200 24624 10000 24744
rect 9200 24080 10000 24200
rect 9200 23536 10000 23656
rect 9200 22992 10000 23112
rect 9200 22448 10000 22568
rect 9200 21904 10000 22024
rect 9200 21360 10000 21480
rect 9200 20816 10000 20936
rect 9200 20272 10000 20392
rect 9200 19728 10000 19848
rect 9200 19184 10000 19304
rect 9200 18776 10000 18896
rect 9200 18232 10000 18352
rect 9200 17688 10000 17808
rect 9200 17144 10000 17264
rect 9200 16600 10000 16720
rect 9200 16056 10000 16176
rect 9200 15512 10000 15632
rect 9200 14968 10000 15088
rect 9200 14424 10000 14544
rect 9200 13880 10000 14000
rect 9200 13336 10000 13456
rect 9200 12792 10000 12912
rect 9200 12384 10000 12504
rect 9200 11840 10000 11960
rect 9200 11296 10000 11416
rect 9200 10752 10000 10872
rect 9200 10208 10000 10328
rect 9200 9664 10000 9784
rect 9200 9120 10000 9240
rect 9200 8576 10000 8696
rect 9200 8032 10000 8152
rect 9200 7488 10000 7608
rect 9200 6944 10000 7064
rect 9200 6400 10000 6520
rect 9200 5992 10000 6112
rect 9200 5448 10000 5568
rect 9200 4904 10000 5024
rect 9200 4360 10000 4480
rect 9200 3816 10000 3936
rect 9200 3272 10000 3392
rect 9200 2728 10000 2848
rect 9200 2184 10000 2304
rect 9200 1640 10000 1760
rect 9200 1096 10000 1216
rect 9200 552 10000 672
rect 9200 144 10000 264
<< obsm3 >>
rect 2242 24544 9120 24717
rect 2242 24280 9200 24544
rect 2242 24000 9120 24280
rect 2242 23736 9200 24000
rect 2242 23456 9120 23736
rect 2242 23192 9200 23456
rect 2242 22912 9120 23192
rect 2242 22648 9200 22912
rect 2242 22368 9120 22648
rect 2242 22104 9200 22368
rect 2242 21824 9120 22104
rect 2242 21560 9200 21824
rect 2242 21280 9120 21560
rect 2242 21016 9200 21280
rect 2242 20736 9120 21016
rect 2242 20472 9200 20736
rect 2242 20192 9120 20472
rect 2242 19928 9200 20192
rect 2242 19648 9120 19928
rect 2242 19384 9200 19648
rect 2242 19104 9120 19384
rect 2242 18976 9200 19104
rect 2242 18696 9120 18976
rect 2242 18432 9200 18696
rect 2242 18152 9120 18432
rect 2242 17888 9200 18152
rect 2242 17608 9120 17888
rect 2242 17344 9200 17608
rect 2242 17064 9120 17344
rect 2242 16800 9200 17064
rect 2242 16520 9120 16800
rect 2242 16256 9200 16520
rect 2242 15976 9120 16256
rect 2242 15712 9200 15976
rect 2242 15432 9120 15712
rect 2242 15168 9200 15432
rect 2242 14888 9120 15168
rect 2242 14624 9200 14888
rect 2242 14344 9120 14624
rect 2242 14080 9200 14344
rect 2242 13800 9120 14080
rect 2242 13536 9200 13800
rect 2242 13256 9120 13536
rect 2242 12992 9200 13256
rect 2242 12712 9120 12992
rect 2242 12584 9200 12712
rect 2242 12304 9120 12584
rect 2242 12040 9200 12304
rect 2242 11760 9120 12040
rect 2242 11496 9200 11760
rect 2242 11216 9120 11496
rect 2242 10952 9200 11216
rect 2242 10672 9120 10952
rect 2242 10408 9200 10672
rect 2242 10128 9120 10408
rect 2242 9864 9200 10128
rect 2242 9584 9120 9864
rect 2242 9320 9200 9584
rect 2242 9040 9120 9320
rect 2242 8776 9200 9040
rect 2242 8496 9120 8776
rect 2242 8232 9200 8496
rect 2242 7952 9120 8232
rect 2242 7688 9200 7952
rect 2242 7408 9120 7688
rect 2242 7144 9200 7408
rect 2242 6864 9120 7144
rect 2242 6600 9200 6864
rect 2242 6320 9120 6600
rect 2242 6192 9200 6320
rect 2242 5912 9120 6192
rect 2242 5648 9200 5912
rect 2242 5368 9120 5648
rect 2242 5104 9200 5368
rect 2242 4824 9120 5104
rect 2242 4560 9200 4824
rect 2242 4280 9120 4560
rect 2242 4016 9200 4280
rect 2242 3736 9120 4016
rect 2242 3472 9200 3736
rect 2242 3192 9120 3472
rect 2242 2928 9200 3192
rect 2242 2648 9120 2928
rect 2242 2384 9200 2648
rect 2242 2104 9120 2384
rect 2242 1840 9200 2104
rect 2242 1560 9120 1840
rect 2242 1296 9200 1560
rect 2242 1016 9120 1296
rect 2242 752 9200 1016
rect 2242 472 9120 752
rect 2242 344 9200 472
rect 2242 171 9120 344
<< metal4 >>
rect 2242 2128 2562 22352
rect 3542 2128 3862 22352
rect 4840 2128 5160 22352
rect 6139 2128 6459 22352
rect 7437 2128 7757 22352
<< obsm4 >>
rect 3942 2128 4760 22352
rect 5240 2128 6059 22352
<< labels >>
rlabel metal2 s 4986 0 5042 800 6 clk
port 1 nsew signal input
rlabel metal3 s 9200 144 10000 264 6 core0Index[0]
port 2 nsew signal output
rlabel metal3 s 9200 552 10000 672 6 core0Index[1]
port 3 nsew signal output
rlabel metal3 s 9200 1096 10000 1216 6 core0Index[2]
port 4 nsew signal output
rlabel metal3 s 9200 1640 10000 1760 6 core0Index[3]
port 5 nsew signal output
rlabel metal3 s 9200 2184 10000 2304 6 core0Index[4]
port 6 nsew signal output
rlabel metal3 s 9200 2728 10000 2848 6 core0Index[5]
port 7 nsew signal output
rlabel metal3 s 9200 3272 10000 3392 6 core0Index[6]
port 8 nsew signal output
rlabel metal3 s 9200 3816 10000 3936 6 core0Index[7]
port 9 nsew signal output
rlabel metal3 s 9200 4360 10000 4480 6 core1Index[0]
port 10 nsew signal output
rlabel metal3 s 9200 4904 10000 5024 6 core1Index[1]
port 11 nsew signal output
rlabel metal3 s 9200 5448 10000 5568 6 core1Index[2]
port 12 nsew signal output
rlabel metal3 s 9200 5992 10000 6112 6 core1Index[3]
port 13 nsew signal output
rlabel metal3 s 9200 6400 10000 6520 6 core1Index[4]
port 14 nsew signal output
rlabel metal3 s 9200 6944 10000 7064 6 core1Index[5]
port 15 nsew signal output
rlabel metal3 s 9200 7488 10000 7608 6 core1Index[6]
port 16 nsew signal output
rlabel metal3 s 9200 8032 10000 8152 6 core1Index[7]
port 17 nsew signal output
rlabel metal3 s 9200 8576 10000 8696 6 manufacturerID[0]
port 18 nsew signal output
rlabel metal3 s 9200 13880 10000 14000 6 manufacturerID[10]
port 19 nsew signal output
rlabel metal3 s 9200 9120 10000 9240 6 manufacturerID[1]
port 20 nsew signal output
rlabel metal3 s 9200 9664 10000 9784 6 manufacturerID[2]
port 21 nsew signal output
rlabel metal3 s 9200 10208 10000 10328 6 manufacturerID[3]
port 22 nsew signal output
rlabel metal3 s 9200 10752 10000 10872 6 manufacturerID[4]
port 23 nsew signal output
rlabel metal3 s 9200 11296 10000 11416 6 manufacturerID[5]
port 24 nsew signal output
rlabel metal3 s 9200 11840 10000 11960 6 manufacturerID[6]
port 25 nsew signal output
rlabel metal3 s 9200 12384 10000 12504 6 manufacturerID[7]
port 26 nsew signal output
rlabel metal3 s 9200 12792 10000 12912 6 manufacturerID[8]
port 27 nsew signal output
rlabel metal3 s 9200 13336 10000 13456 6 manufacturerID[9]
port 28 nsew signal output
rlabel metal3 s 9200 14424 10000 14544 6 partID[0]
port 29 nsew signal output
rlabel metal3 s 9200 19728 10000 19848 6 partID[10]
port 30 nsew signal output
rlabel metal3 s 9200 20272 10000 20392 6 partID[11]
port 31 nsew signal output
rlabel metal3 s 9200 20816 10000 20936 6 partID[12]
port 32 nsew signal output
rlabel metal3 s 9200 21360 10000 21480 6 partID[13]
port 33 nsew signal output
rlabel metal3 s 9200 21904 10000 22024 6 partID[14]
port 34 nsew signal output
rlabel metal3 s 9200 22448 10000 22568 6 partID[15]
port 35 nsew signal output
rlabel metal3 s 9200 14968 10000 15088 6 partID[1]
port 36 nsew signal output
rlabel metal3 s 9200 15512 10000 15632 6 partID[2]
port 37 nsew signal output
rlabel metal3 s 9200 16056 10000 16176 6 partID[3]
port 38 nsew signal output
rlabel metal3 s 9200 16600 10000 16720 6 partID[4]
port 39 nsew signal output
rlabel metal3 s 9200 17144 10000 17264 6 partID[5]
port 40 nsew signal output
rlabel metal3 s 9200 17688 10000 17808 6 partID[6]
port 41 nsew signal output
rlabel metal3 s 9200 18232 10000 18352 6 partID[7]
port 42 nsew signal output
rlabel metal3 s 9200 18776 10000 18896 6 partID[8]
port 43 nsew signal output
rlabel metal3 s 9200 19184 10000 19304 6 partID[9]
port 44 nsew signal output
rlabel metal4 s 2242 2128 2562 22352 6 vccd1
port 45 nsew power input
rlabel metal4 s 4840 2128 5160 22352 6 vccd1
port 45 nsew power input
rlabel metal4 s 7437 2128 7757 22352 6 vccd1
port 45 nsew power input
rlabel metal3 s 9200 22992 10000 23112 6 versionID[0]
port 46 nsew signal output
rlabel metal3 s 9200 23536 10000 23656 6 versionID[1]
port 47 nsew signal output
rlabel metal3 s 9200 24080 10000 24200 6 versionID[2]
port 48 nsew signal output
rlabel metal3 s 9200 24624 10000 24744 6 versionID[3]
port 49 nsew signal output
rlabel metal4 s 3542 2128 3862 22352 6 vssd1
port 50 nsew ground input
rlabel metal4 s 6139 2128 6459 22352 6 vssd1
port 50 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 10000 25000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 206044
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Configuration/runs/Configuration/results/finishing/Configuration.magic.gds
string GDS_START 20970
<< end >>

