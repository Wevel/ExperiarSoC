VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO IOMultiplexer
  CLASS BLOCK ;
  FOREIGN IOMultiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 230.000 BY 200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END clk
  PIN config_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END config_address[0]
  PIN config_address[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END config_address[10]
  PIN config_address[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END config_address[11]
  PIN config_address[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END config_address[12]
  PIN config_address[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END config_address[13]
  PIN config_address[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END config_address[14]
  PIN config_address[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END config_address[15]
  PIN config_address[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END config_address[16]
  PIN config_address[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END config_address[17]
  PIN config_address[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END config_address[18]
  PIN config_address[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END config_address[19]
  PIN config_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END config_address[1]
  PIN config_address[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END config_address[20]
  PIN config_address[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END config_address[21]
  PIN config_address[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END config_address[22]
  PIN config_address[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END config_address[23]
  PIN config_address[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END config_address[24]
  PIN config_address[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END config_address[25]
  PIN config_address[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END config_address[26]
  PIN config_address[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END config_address[27]
  PIN config_address[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END config_address[28]
  PIN config_address[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END config_address[29]
  PIN config_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END config_address[2]
  PIN config_address[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END config_address[30]
  PIN config_address[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END config_address[31]
  PIN config_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END config_address[3]
  PIN config_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END config_address[4]
  PIN config_address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END config_address[5]
  PIN config_address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END config_address[6]
  PIN config_address[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END config_address[7]
  PIN config_address[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END config_address[8]
  PIN config_address[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END config_address[9]
  PIN config_data[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END config_data[0]
  PIN config_data[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END config_data[10]
  PIN config_data[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END config_data[11]
  PIN config_data[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END config_data[12]
  PIN config_data[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END config_data[13]
  PIN config_data[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END config_data[14]
  PIN config_data[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END config_data[15]
  PIN config_data[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END config_data[16]
  PIN config_data[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END config_data[17]
  PIN config_data[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END config_data[18]
  PIN config_data[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END config_data[19]
  PIN config_data[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END config_data[1]
  PIN config_data[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END config_data[20]
  PIN config_data[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END config_data[21]
  PIN config_data[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END config_data[22]
  PIN config_data[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END config_data[23]
  PIN config_data[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END config_data[24]
  PIN config_data[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END config_data[25]
  PIN config_data[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END config_data[26]
  PIN config_data[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END config_data[27]
  PIN config_data[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END config_data[28]
  PIN config_data[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END config_data[29]
  PIN config_data[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END config_data[2]
  PIN config_data[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END config_data[30]
  PIN config_data[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END config_data[31]
  PIN config_data[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END config_data[3]
  PIN config_data[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END config_data[4]
  PIN config_data[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END config_data[5]
  PIN config_data[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END config_data[6]
  PIN config_data[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END config_data[7]
  PIN config_data[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END config_data[8]
  PIN config_data[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END config_data[9]
  PIN config_oe
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END config_oe
  PIN config_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END config_we
  PIN gpio0_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END gpio0_input[0]
  PIN gpio0_input[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END gpio0_input[10]
  PIN gpio0_input[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END gpio0_input[11]
  PIN gpio0_input[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END gpio0_input[12]
  PIN gpio0_input[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END gpio0_input[13]
  PIN gpio0_input[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END gpio0_input[14]
  PIN gpio0_input[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END gpio0_input[15]
  PIN gpio0_input[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END gpio0_input[16]
  PIN gpio0_input[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END gpio0_input[17]
  PIN gpio0_input[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END gpio0_input[18]
  PIN gpio0_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END gpio0_input[1]
  PIN gpio0_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END gpio0_input[2]
  PIN gpio0_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END gpio0_input[3]
  PIN gpio0_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END gpio0_input[4]
  PIN gpio0_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END gpio0_input[5]
  PIN gpio0_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END gpio0_input[6]
  PIN gpio0_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END gpio0_input[7]
  PIN gpio0_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END gpio0_input[8]
  PIN gpio0_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END gpio0_input[9]
  PIN gpio0_oe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END gpio0_oe[0]
  PIN gpio0_oe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END gpio0_oe[10]
  PIN gpio0_oe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END gpio0_oe[11]
  PIN gpio0_oe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END gpio0_oe[12]
  PIN gpio0_oe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END gpio0_oe[13]
  PIN gpio0_oe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END gpio0_oe[14]
  PIN gpio0_oe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END gpio0_oe[15]
  PIN gpio0_oe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END gpio0_oe[16]
  PIN gpio0_oe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END gpio0_oe[17]
  PIN gpio0_oe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END gpio0_oe[18]
  PIN gpio0_oe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END gpio0_oe[1]
  PIN gpio0_oe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END gpio0_oe[2]
  PIN gpio0_oe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END gpio0_oe[3]
  PIN gpio0_oe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END gpio0_oe[4]
  PIN gpio0_oe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END gpio0_oe[5]
  PIN gpio0_oe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END gpio0_oe[6]
  PIN gpio0_oe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END gpio0_oe[7]
  PIN gpio0_oe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END gpio0_oe[8]
  PIN gpio0_oe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END gpio0_oe[9]
  PIN gpio0_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END gpio0_output[0]
  PIN gpio0_output[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END gpio0_output[10]
  PIN gpio0_output[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END gpio0_output[11]
  PIN gpio0_output[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END gpio0_output[12]
  PIN gpio0_output[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END gpio0_output[13]
  PIN gpio0_output[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END gpio0_output[14]
  PIN gpio0_output[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END gpio0_output[15]
  PIN gpio0_output[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END gpio0_output[16]
  PIN gpio0_output[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END gpio0_output[17]
  PIN gpio0_output[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END gpio0_output[18]
  PIN gpio0_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END gpio0_output[1]
  PIN gpio0_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END gpio0_output[2]
  PIN gpio0_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END gpio0_output[3]
  PIN gpio0_output[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END gpio0_output[4]
  PIN gpio0_output[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END gpio0_output[5]
  PIN gpio0_output[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END gpio0_output[6]
  PIN gpio0_output[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END gpio0_output[7]
  PIN gpio0_output[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END gpio0_output[8]
  PIN gpio0_output[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END gpio0_output[9]
  PIN gpio1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END gpio1_input[0]
  PIN gpio1_input[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END gpio1_input[10]
  PIN gpio1_input[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END gpio1_input[11]
  PIN gpio1_input[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END gpio1_input[12]
  PIN gpio1_input[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END gpio1_input[13]
  PIN gpio1_input[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END gpio1_input[14]
  PIN gpio1_input[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END gpio1_input[15]
  PIN gpio1_input[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END gpio1_input[16]
  PIN gpio1_input[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END gpio1_input[17]
  PIN gpio1_input[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END gpio1_input[18]
  PIN gpio1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END gpio1_input[1]
  PIN gpio1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END gpio1_input[2]
  PIN gpio1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END gpio1_input[3]
  PIN gpio1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END gpio1_input[4]
  PIN gpio1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END gpio1_input[5]
  PIN gpio1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END gpio1_input[6]
  PIN gpio1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END gpio1_input[7]
  PIN gpio1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END gpio1_input[8]
  PIN gpio1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END gpio1_input[9]
  PIN gpio1_oe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END gpio1_oe[0]
  PIN gpio1_oe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END gpio1_oe[10]
  PIN gpio1_oe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END gpio1_oe[11]
  PIN gpio1_oe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END gpio1_oe[12]
  PIN gpio1_oe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END gpio1_oe[13]
  PIN gpio1_oe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END gpio1_oe[14]
  PIN gpio1_oe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END gpio1_oe[15]
  PIN gpio1_oe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END gpio1_oe[16]
  PIN gpio1_oe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END gpio1_oe[17]
  PIN gpio1_oe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END gpio1_oe[18]
  PIN gpio1_oe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END gpio1_oe[1]
  PIN gpio1_oe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END gpio1_oe[2]
  PIN gpio1_oe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END gpio1_oe[3]
  PIN gpio1_oe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END gpio1_oe[4]
  PIN gpio1_oe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END gpio1_oe[5]
  PIN gpio1_oe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END gpio1_oe[6]
  PIN gpio1_oe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END gpio1_oe[7]
  PIN gpio1_oe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END gpio1_oe[8]
  PIN gpio1_oe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END gpio1_oe[9]
  PIN gpio1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END gpio1_output[0]
  PIN gpio1_output[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END gpio1_output[10]
  PIN gpio1_output[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END gpio1_output[11]
  PIN gpio1_output[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END gpio1_output[12]
  PIN gpio1_output[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END gpio1_output[13]
  PIN gpio1_output[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END gpio1_output[14]
  PIN gpio1_output[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END gpio1_output[15]
  PIN gpio1_output[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END gpio1_output[16]
  PIN gpio1_output[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END gpio1_output[17]
  PIN gpio1_output[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END gpio1_output[18]
  PIN gpio1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END gpio1_output[1]
  PIN gpio1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END gpio1_output[2]
  PIN gpio1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END gpio1_output[3]
  PIN gpio1_output[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END gpio1_output[4]
  PIN gpio1_output[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END gpio1_output[5]
  PIN gpio1_output[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END gpio1_output[6]
  PIN gpio1_output[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END gpio1_output[7]
  PIN gpio1_output[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END gpio1_output[8]
  PIN gpio1_output[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END gpio1_output[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 196.000 1.290 200.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 196.000 61.550 200.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 196.000 67.530 200.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 196.000 73.510 200.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 196.000 79.950 200.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 196.000 85.930 200.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 196.000 91.910 200.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 196.000 97.890 200.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 196.000 103.870 200.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 196.000 109.850 200.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 196.000 116.290 200.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 196.000 7.270 200.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 196.000 122.270 200.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 196.000 128.250 200.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 196.000 134.230 200.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 196.000 140.210 200.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 196.000 146.190 200.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 196.000 152.170 200.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 196.000 158.610 200.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 196.000 164.590 200.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 196.000 170.570 200.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 196.000 176.550 200.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 196.000 13.250 200.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 196.000 182.530 200.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 196.000 188.510 200.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 196.000 194.950 200.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 196.000 200.930 200.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 196.000 206.910 200.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 196.000 212.890 200.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 196.000 218.870 200.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 196.000 224.850 200.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 196.000 19.230 200.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 196.000 25.210 200.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 196.000 31.190 200.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 196.000 37.170 200.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 196.000 43.610 200.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 196.000 49.590 200.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 196.000 55.570 200.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 196.000 3.130 200.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 196.000 63.390 200.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 196.000 69.830 200.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 196.000 75.810 200.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 196.000 81.790 200.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 196.000 87.770 200.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 196.000 93.750 200.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 196.000 99.730 200.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 196.000 106.170 200.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 196.000 112.150 200.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 196.000 118.130 200.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 196.000 9.110 200.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 196.000 124.110 200.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 196.000 130.090 200.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 196.000 136.070 200.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 196.000 142.510 200.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 196.000 148.490 200.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 196.000 154.470 200.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 196.000 160.450 200.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 196.000 166.430 200.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 196.000 172.410 200.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 196.000 178.390 200.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 196.000 15.090 200.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 196.000 184.830 200.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 196.000 190.810 200.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 196.000 196.790 200.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 196.000 202.770 200.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 196.000 208.750 200.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 196.000 214.730 200.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 196.000 221.170 200.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 196.000 227.150 200.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 196.000 21.070 200.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 196.000 27.510 200.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 196.000 33.490 200.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 196.000 39.470 200.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 196.000 45.450 200.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 196.000 51.430 200.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 196.000 57.410 200.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 196.000 4.970 200.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 196.000 65.690 200.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 196.000 71.670 200.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 196.000 77.650 200.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 196.000 83.630 200.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 196.000 89.610 200.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 196.000 96.050 200.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 196.000 102.030 200.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 196.000 108.010 200.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 196.000 113.990 200.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 196.000 119.970 200.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 196.000 10.950 200.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 196.000 125.950 200.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 196.000 132.390 200.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 196.000 138.370 200.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 196.000 144.350 200.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 196.000 150.330 200.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 196.000 156.310 200.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 196.000 162.290 200.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 196.000 168.730 200.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 196.000 174.710 200.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 196.000 180.690 200.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 196.000 17.390 200.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 196.000 186.670 200.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 196.000 192.650 200.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 196.000 198.630 200.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 196.000 204.610 200.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 196.000 211.050 200.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 196.000 217.030 200.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 196.000 223.010 200.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 196.000 228.990 200.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 196.000 23.370 200.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 196.000 29.350 200.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 196.000 35.330 200.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 196.000 41.310 200.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 196.000 47.290 200.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 196.000 53.730 200.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 196.000 59.710 200.000 ;
    END
  END io_out[9]
  PIN la_blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 49.680 230.000 50.280 ;
    END
  END la_blink[0]
  PIN la_blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 149.640 230.000 150.240 ;
    END
  END la_blink[1]
  PIN pwm_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END pwm_out[0]
  PIN pwm_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END pwm_out[10]
  PIN pwm_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END pwm_out[11]
  PIN pwm_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END pwm_out[12]
  PIN pwm_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END pwm_out[13]
  PIN pwm_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END pwm_out[14]
  PIN pwm_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END pwm_out[15]
  PIN pwm_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END pwm_out[1]
  PIN pwm_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END pwm_out[2]
  PIN pwm_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END pwm_out[3]
  PIN pwm_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END pwm_out[4]
  PIN pwm_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END pwm_out[5]
  PIN pwm_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END pwm_out[6]
  PIN pwm_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END pwm_out[7]
  PIN pwm_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END pwm_out[8]
  PIN pwm_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END pwm_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END rst
  PIN spi_clk[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END spi_clk[0]
  PIN spi_clk[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END spi_clk[1]
  PIN spi_cs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END spi_cs[0]
  PIN spi_cs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END spi_cs[1]
  PIN spi_miso[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END spi_miso[0]
  PIN spi_miso[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END spi_miso[1]
  PIN spi_mosi[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END spi_mosi[0]
  PIN spi_mosi[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END spi_mosi[1]
  PIN uart_rx[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END uart_rx[0]
  PIN uart_rx[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END uart_rx[1]
  PIN uart_rx[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END uart_rx[2]
  PIN uart_rx[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END uart_rx[3]
  PIN uart_tx[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END uart_tx[0]
  PIN uart_tx[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END uart_tx[1]
  PIN uart_tx[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END uart_tx[2]
  PIN uart_tx[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END uart_tx[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 224.480 187.765 ;
      LAYER met1 ;
        RECT 0.070 0.040 229.010 190.360 ;
      LAYER met2 ;
        RECT 0.090 195.720 0.730 198.405 ;
        RECT 1.570 195.720 2.570 198.405 ;
        RECT 3.410 195.720 4.410 198.405 ;
        RECT 5.250 195.720 6.710 198.405 ;
        RECT 7.550 195.720 8.550 198.405 ;
        RECT 9.390 195.720 10.390 198.405 ;
        RECT 11.230 195.720 12.690 198.405 ;
        RECT 13.530 195.720 14.530 198.405 ;
        RECT 15.370 195.720 16.830 198.405 ;
        RECT 17.670 195.720 18.670 198.405 ;
        RECT 19.510 195.720 20.510 198.405 ;
        RECT 21.350 195.720 22.810 198.405 ;
        RECT 23.650 195.720 24.650 198.405 ;
        RECT 25.490 195.720 26.950 198.405 ;
        RECT 27.790 195.720 28.790 198.405 ;
        RECT 29.630 195.720 30.630 198.405 ;
        RECT 31.470 195.720 32.930 198.405 ;
        RECT 33.770 195.720 34.770 198.405 ;
        RECT 35.610 195.720 36.610 198.405 ;
        RECT 37.450 195.720 38.910 198.405 ;
        RECT 39.750 195.720 40.750 198.405 ;
        RECT 41.590 195.720 43.050 198.405 ;
        RECT 43.890 195.720 44.890 198.405 ;
        RECT 45.730 195.720 46.730 198.405 ;
        RECT 47.570 195.720 49.030 198.405 ;
        RECT 49.870 195.720 50.870 198.405 ;
        RECT 51.710 195.720 53.170 198.405 ;
        RECT 54.010 195.720 55.010 198.405 ;
        RECT 55.850 195.720 56.850 198.405 ;
        RECT 57.690 195.720 59.150 198.405 ;
        RECT 59.990 195.720 60.990 198.405 ;
        RECT 61.830 195.720 62.830 198.405 ;
        RECT 63.670 195.720 65.130 198.405 ;
        RECT 65.970 195.720 66.970 198.405 ;
        RECT 67.810 195.720 69.270 198.405 ;
        RECT 70.110 195.720 71.110 198.405 ;
        RECT 71.950 195.720 72.950 198.405 ;
        RECT 73.790 195.720 75.250 198.405 ;
        RECT 76.090 195.720 77.090 198.405 ;
        RECT 77.930 195.720 79.390 198.405 ;
        RECT 80.230 195.720 81.230 198.405 ;
        RECT 82.070 195.720 83.070 198.405 ;
        RECT 83.910 195.720 85.370 198.405 ;
        RECT 86.210 195.720 87.210 198.405 ;
        RECT 88.050 195.720 89.050 198.405 ;
        RECT 89.890 195.720 91.350 198.405 ;
        RECT 92.190 195.720 93.190 198.405 ;
        RECT 94.030 195.720 95.490 198.405 ;
        RECT 96.330 195.720 97.330 198.405 ;
        RECT 98.170 195.720 99.170 198.405 ;
        RECT 100.010 195.720 101.470 198.405 ;
        RECT 102.310 195.720 103.310 198.405 ;
        RECT 104.150 195.720 105.610 198.405 ;
        RECT 106.450 195.720 107.450 198.405 ;
        RECT 108.290 195.720 109.290 198.405 ;
        RECT 110.130 195.720 111.590 198.405 ;
        RECT 112.430 195.720 113.430 198.405 ;
        RECT 114.270 195.720 115.730 198.405 ;
        RECT 116.570 195.720 117.570 198.405 ;
        RECT 118.410 195.720 119.410 198.405 ;
        RECT 120.250 195.720 121.710 198.405 ;
        RECT 122.550 195.720 123.550 198.405 ;
        RECT 124.390 195.720 125.390 198.405 ;
        RECT 126.230 195.720 127.690 198.405 ;
        RECT 128.530 195.720 129.530 198.405 ;
        RECT 130.370 195.720 131.830 198.405 ;
        RECT 132.670 195.720 133.670 198.405 ;
        RECT 134.510 195.720 135.510 198.405 ;
        RECT 136.350 195.720 137.810 198.405 ;
        RECT 138.650 195.720 139.650 198.405 ;
        RECT 140.490 195.720 141.950 198.405 ;
        RECT 142.790 195.720 143.790 198.405 ;
        RECT 144.630 195.720 145.630 198.405 ;
        RECT 146.470 195.720 147.930 198.405 ;
        RECT 148.770 195.720 149.770 198.405 ;
        RECT 150.610 195.720 151.610 198.405 ;
        RECT 152.450 195.720 153.910 198.405 ;
        RECT 154.750 195.720 155.750 198.405 ;
        RECT 156.590 195.720 158.050 198.405 ;
        RECT 158.890 195.720 159.890 198.405 ;
        RECT 160.730 195.720 161.730 198.405 ;
        RECT 162.570 195.720 164.030 198.405 ;
        RECT 164.870 195.720 165.870 198.405 ;
        RECT 166.710 195.720 168.170 198.405 ;
        RECT 169.010 195.720 170.010 198.405 ;
        RECT 170.850 195.720 171.850 198.405 ;
        RECT 172.690 195.720 174.150 198.405 ;
        RECT 174.990 195.720 175.990 198.405 ;
        RECT 176.830 195.720 177.830 198.405 ;
        RECT 178.670 195.720 180.130 198.405 ;
        RECT 180.970 195.720 181.970 198.405 ;
        RECT 182.810 195.720 184.270 198.405 ;
        RECT 185.110 195.720 186.110 198.405 ;
        RECT 186.950 195.720 187.950 198.405 ;
        RECT 188.790 195.720 190.250 198.405 ;
        RECT 191.090 195.720 192.090 198.405 ;
        RECT 192.930 195.720 194.390 198.405 ;
        RECT 195.230 195.720 196.230 198.405 ;
        RECT 197.070 195.720 198.070 198.405 ;
        RECT 198.910 195.720 200.370 198.405 ;
        RECT 201.210 195.720 202.210 198.405 ;
        RECT 203.050 195.720 204.050 198.405 ;
        RECT 204.890 195.720 206.350 198.405 ;
        RECT 207.190 195.720 208.190 198.405 ;
        RECT 209.030 195.720 210.490 198.405 ;
        RECT 211.330 195.720 212.330 198.405 ;
        RECT 213.170 195.720 214.170 198.405 ;
        RECT 215.010 195.720 216.470 198.405 ;
        RECT 217.310 195.720 218.310 198.405 ;
        RECT 219.150 195.720 220.610 198.405 ;
        RECT 221.450 195.720 222.450 198.405 ;
        RECT 223.290 195.720 224.290 198.405 ;
        RECT 225.130 195.720 226.590 198.405 ;
        RECT 227.430 195.720 228.430 198.405 ;
        RECT 0.090 4.280 228.980 195.720 ;
        RECT 0.090 0.010 0.270 4.280 ;
        RECT 1.110 0.010 1.650 4.280 ;
        RECT 2.490 0.010 3.030 4.280 ;
        RECT 3.870 0.010 4.870 4.280 ;
        RECT 5.710 0.010 6.250 4.280 ;
        RECT 7.090 0.010 8.090 4.280 ;
        RECT 8.930 0.010 9.470 4.280 ;
        RECT 10.310 0.010 10.850 4.280 ;
        RECT 11.690 0.010 12.690 4.280 ;
        RECT 13.530 0.010 14.070 4.280 ;
        RECT 14.910 0.010 15.910 4.280 ;
        RECT 16.750 0.010 17.290 4.280 ;
        RECT 18.130 0.010 19.130 4.280 ;
        RECT 19.970 0.010 20.510 4.280 ;
        RECT 21.350 0.010 21.890 4.280 ;
        RECT 22.730 0.010 23.730 4.280 ;
        RECT 24.570 0.010 25.110 4.280 ;
        RECT 25.950 0.010 26.950 4.280 ;
        RECT 27.790 0.010 28.330 4.280 ;
        RECT 29.170 0.010 30.170 4.280 ;
        RECT 31.010 0.010 31.550 4.280 ;
        RECT 32.390 0.010 32.930 4.280 ;
        RECT 33.770 0.010 34.770 4.280 ;
        RECT 35.610 0.010 36.150 4.280 ;
        RECT 36.990 0.010 37.990 4.280 ;
        RECT 38.830 0.010 39.370 4.280 ;
        RECT 40.210 0.010 41.210 4.280 ;
        RECT 42.050 0.010 42.590 4.280 ;
        RECT 43.430 0.010 43.970 4.280 ;
        RECT 44.810 0.010 45.810 4.280 ;
        RECT 46.650 0.010 47.190 4.280 ;
        RECT 48.030 0.010 49.030 4.280 ;
        RECT 49.870 0.010 50.410 4.280 ;
        RECT 51.250 0.010 52.250 4.280 ;
        RECT 53.090 0.010 53.630 4.280 ;
        RECT 54.470 0.010 55.010 4.280 ;
        RECT 55.850 0.010 56.850 4.280 ;
        RECT 57.690 0.010 58.230 4.280 ;
        RECT 59.070 0.010 60.070 4.280 ;
        RECT 60.910 0.010 61.450 4.280 ;
        RECT 62.290 0.010 62.830 4.280 ;
        RECT 63.670 0.010 64.670 4.280 ;
        RECT 65.510 0.010 66.050 4.280 ;
        RECT 66.890 0.010 67.890 4.280 ;
        RECT 68.730 0.010 69.270 4.280 ;
        RECT 70.110 0.010 71.110 4.280 ;
        RECT 71.950 0.010 72.490 4.280 ;
        RECT 73.330 0.010 73.870 4.280 ;
        RECT 74.710 0.010 75.710 4.280 ;
        RECT 76.550 0.010 77.090 4.280 ;
        RECT 77.930 0.010 78.930 4.280 ;
        RECT 79.770 0.010 80.310 4.280 ;
        RECT 81.150 0.010 82.150 4.280 ;
        RECT 82.990 0.010 83.530 4.280 ;
        RECT 84.370 0.010 84.910 4.280 ;
        RECT 85.750 0.010 86.750 4.280 ;
        RECT 87.590 0.010 88.130 4.280 ;
        RECT 88.970 0.010 89.970 4.280 ;
        RECT 90.810 0.010 91.350 4.280 ;
        RECT 92.190 0.010 93.190 4.280 ;
        RECT 94.030 0.010 94.570 4.280 ;
        RECT 95.410 0.010 95.950 4.280 ;
        RECT 96.790 0.010 97.790 4.280 ;
        RECT 98.630 0.010 99.170 4.280 ;
        RECT 100.010 0.010 101.010 4.280 ;
        RECT 101.850 0.010 102.390 4.280 ;
        RECT 103.230 0.010 104.230 4.280 ;
        RECT 105.070 0.010 105.610 4.280 ;
        RECT 106.450 0.010 106.990 4.280 ;
        RECT 107.830 0.010 108.830 4.280 ;
        RECT 109.670 0.010 110.210 4.280 ;
        RECT 111.050 0.010 112.050 4.280 ;
        RECT 112.890 0.010 113.430 4.280 ;
        RECT 114.270 0.010 115.270 4.280 ;
        RECT 116.110 0.010 116.650 4.280 ;
        RECT 117.490 0.010 118.030 4.280 ;
        RECT 118.870 0.010 119.870 4.280 ;
        RECT 120.710 0.010 121.250 4.280 ;
        RECT 122.090 0.010 123.090 4.280 ;
        RECT 123.930 0.010 124.470 4.280 ;
        RECT 125.310 0.010 125.850 4.280 ;
        RECT 126.690 0.010 127.690 4.280 ;
        RECT 128.530 0.010 129.070 4.280 ;
        RECT 129.910 0.010 130.910 4.280 ;
        RECT 131.750 0.010 132.290 4.280 ;
        RECT 133.130 0.010 134.130 4.280 ;
        RECT 134.970 0.010 135.510 4.280 ;
        RECT 136.350 0.010 136.890 4.280 ;
        RECT 137.730 0.010 138.730 4.280 ;
        RECT 139.570 0.010 140.110 4.280 ;
        RECT 140.950 0.010 141.950 4.280 ;
        RECT 142.790 0.010 143.330 4.280 ;
        RECT 144.170 0.010 145.170 4.280 ;
        RECT 146.010 0.010 146.550 4.280 ;
        RECT 147.390 0.010 147.930 4.280 ;
        RECT 148.770 0.010 149.770 4.280 ;
        RECT 150.610 0.010 151.150 4.280 ;
        RECT 151.990 0.010 152.990 4.280 ;
        RECT 153.830 0.010 154.370 4.280 ;
        RECT 155.210 0.010 156.210 4.280 ;
        RECT 157.050 0.010 157.590 4.280 ;
        RECT 158.430 0.010 158.970 4.280 ;
        RECT 159.810 0.010 160.810 4.280 ;
        RECT 161.650 0.010 162.190 4.280 ;
        RECT 163.030 0.010 164.030 4.280 ;
        RECT 164.870 0.010 165.410 4.280 ;
        RECT 166.250 0.010 167.250 4.280 ;
        RECT 168.090 0.010 168.630 4.280 ;
        RECT 169.470 0.010 170.010 4.280 ;
        RECT 170.850 0.010 171.850 4.280 ;
        RECT 172.690 0.010 173.230 4.280 ;
        RECT 174.070 0.010 175.070 4.280 ;
        RECT 175.910 0.010 176.450 4.280 ;
        RECT 177.290 0.010 177.830 4.280 ;
        RECT 178.670 0.010 179.670 4.280 ;
        RECT 180.510 0.010 181.050 4.280 ;
        RECT 181.890 0.010 182.890 4.280 ;
        RECT 183.730 0.010 184.270 4.280 ;
        RECT 185.110 0.010 186.110 4.280 ;
        RECT 186.950 0.010 187.490 4.280 ;
        RECT 188.330 0.010 188.870 4.280 ;
        RECT 189.710 0.010 190.710 4.280 ;
        RECT 191.550 0.010 192.090 4.280 ;
        RECT 192.930 0.010 193.930 4.280 ;
        RECT 194.770 0.010 195.310 4.280 ;
        RECT 196.150 0.010 197.150 4.280 ;
        RECT 197.990 0.010 198.530 4.280 ;
        RECT 199.370 0.010 199.910 4.280 ;
        RECT 200.750 0.010 201.750 4.280 ;
        RECT 202.590 0.010 203.130 4.280 ;
        RECT 203.970 0.010 204.970 4.280 ;
        RECT 205.810 0.010 206.350 4.280 ;
        RECT 207.190 0.010 208.190 4.280 ;
        RECT 209.030 0.010 209.570 4.280 ;
        RECT 210.410 0.010 210.950 4.280 ;
        RECT 211.790 0.010 212.790 4.280 ;
        RECT 213.630 0.010 214.170 4.280 ;
        RECT 215.010 0.010 216.010 4.280 ;
        RECT 216.850 0.010 217.390 4.280 ;
        RECT 218.230 0.010 219.230 4.280 ;
        RECT 220.070 0.010 220.610 4.280 ;
        RECT 221.450 0.010 221.990 4.280 ;
        RECT 222.830 0.010 223.830 4.280 ;
        RECT 224.670 0.010 225.210 4.280 ;
        RECT 226.050 0.010 227.050 4.280 ;
        RECT 227.890 0.010 228.430 4.280 ;
      LAYER met3 ;
        RECT 4.400 197.520 226.000 198.385 ;
        RECT 0.065 196.200 226.000 197.520 ;
        RECT 4.400 194.800 226.000 196.200 ;
        RECT 0.065 193.480 226.000 194.800 ;
        RECT 4.400 192.080 226.000 193.480 ;
        RECT 0.065 190.080 226.000 192.080 ;
        RECT 4.400 188.680 226.000 190.080 ;
        RECT 0.065 187.360 226.000 188.680 ;
        RECT 4.400 185.960 226.000 187.360 ;
        RECT 0.065 184.640 226.000 185.960 ;
        RECT 4.400 183.240 226.000 184.640 ;
        RECT 0.065 181.240 226.000 183.240 ;
        RECT 4.400 179.840 226.000 181.240 ;
        RECT 0.065 178.520 226.000 179.840 ;
        RECT 4.400 177.120 226.000 178.520 ;
        RECT 0.065 175.800 226.000 177.120 ;
        RECT 4.400 174.400 226.000 175.800 ;
        RECT 0.065 172.400 226.000 174.400 ;
        RECT 4.400 171.000 226.000 172.400 ;
        RECT 0.065 169.680 226.000 171.000 ;
        RECT 4.400 168.280 226.000 169.680 ;
        RECT 0.065 166.960 226.000 168.280 ;
        RECT 4.400 165.560 226.000 166.960 ;
        RECT 0.065 163.560 226.000 165.560 ;
        RECT 4.400 162.160 226.000 163.560 ;
        RECT 0.065 160.840 226.000 162.160 ;
        RECT 4.400 159.440 226.000 160.840 ;
        RECT 0.065 158.120 226.000 159.440 ;
        RECT 4.400 156.720 226.000 158.120 ;
        RECT 0.065 154.720 226.000 156.720 ;
        RECT 4.400 153.320 226.000 154.720 ;
        RECT 0.065 152.000 226.000 153.320 ;
        RECT 4.400 150.640 226.000 152.000 ;
        RECT 4.400 150.600 225.600 150.640 ;
        RECT 0.065 149.280 225.600 150.600 ;
        RECT 4.400 149.240 225.600 149.280 ;
        RECT 4.400 147.880 226.000 149.240 ;
        RECT 0.065 145.880 226.000 147.880 ;
        RECT 4.400 144.480 226.000 145.880 ;
        RECT 0.065 143.160 226.000 144.480 ;
        RECT 4.400 141.760 226.000 143.160 ;
        RECT 0.065 140.440 226.000 141.760 ;
        RECT 4.400 139.040 226.000 140.440 ;
        RECT 0.065 137.040 226.000 139.040 ;
        RECT 4.400 135.640 226.000 137.040 ;
        RECT 0.065 134.320 226.000 135.640 ;
        RECT 4.400 132.920 226.000 134.320 ;
        RECT 0.065 131.600 226.000 132.920 ;
        RECT 4.400 130.200 226.000 131.600 ;
        RECT 0.065 128.200 226.000 130.200 ;
        RECT 4.400 126.800 226.000 128.200 ;
        RECT 0.065 125.480 226.000 126.800 ;
        RECT 4.400 124.080 226.000 125.480 ;
        RECT 0.065 122.760 226.000 124.080 ;
        RECT 4.400 121.360 226.000 122.760 ;
        RECT 0.065 119.360 226.000 121.360 ;
        RECT 4.400 117.960 226.000 119.360 ;
        RECT 0.065 116.640 226.000 117.960 ;
        RECT 4.400 115.240 226.000 116.640 ;
        RECT 0.065 113.920 226.000 115.240 ;
        RECT 4.400 112.520 226.000 113.920 ;
        RECT 0.065 110.520 226.000 112.520 ;
        RECT 4.400 109.120 226.000 110.520 ;
        RECT 0.065 107.800 226.000 109.120 ;
        RECT 4.400 106.400 226.000 107.800 ;
        RECT 0.065 105.080 226.000 106.400 ;
        RECT 4.400 103.680 226.000 105.080 ;
        RECT 0.065 102.360 226.000 103.680 ;
        RECT 4.400 100.960 226.000 102.360 ;
        RECT 0.065 98.960 226.000 100.960 ;
        RECT 4.400 97.560 226.000 98.960 ;
        RECT 0.065 96.240 226.000 97.560 ;
        RECT 4.400 94.840 226.000 96.240 ;
        RECT 0.065 93.520 226.000 94.840 ;
        RECT 4.400 92.120 226.000 93.520 ;
        RECT 0.065 90.120 226.000 92.120 ;
        RECT 4.400 88.720 226.000 90.120 ;
        RECT 0.065 87.400 226.000 88.720 ;
        RECT 4.400 86.000 226.000 87.400 ;
        RECT 0.065 84.680 226.000 86.000 ;
        RECT 4.400 83.280 226.000 84.680 ;
        RECT 0.065 81.280 226.000 83.280 ;
        RECT 4.400 79.880 226.000 81.280 ;
        RECT 0.065 78.560 226.000 79.880 ;
        RECT 4.400 77.160 226.000 78.560 ;
        RECT 0.065 75.840 226.000 77.160 ;
        RECT 4.400 74.440 226.000 75.840 ;
        RECT 0.065 72.440 226.000 74.440 ;
        RECT 4.400 71.040 226.000 72.440 ;
        RECT 0.065 69.720 226.000 71.040 ;
        RECT 4.400 68.320 226.000 69.720 ;
        RECT 0.065 67.000 226.000 68.320 ;
        RECT 4.400 65.600 226.000 67.000 ;
        RECT 0.065 63.600 226.000 65.600 ;
        RECT 4.400 62.200 226.000 63.600 ;
        RECT 0.065 60.880 226.000 62.200 ;
        RECT 4.400 59.480 226.000 60.880 ;
        RECT 0.065 58.160 226.000 59.480 ;
        RECT 4.400 56.760 226.000 58.160 ;
        RECT 0.065 54.760 226.000 56.760 ;
        RECT 4.400 53.360 226.000 54.760 ;
        RECT 0.065 52.040 226.000 53.360 ;
        RECT 4.400 50.680 226.000 52.040 ;
        RECT 4.400 50.640 225.600 50.680 ;
        RECT 0.065 49.320 225.600 50.640 ;
        RECT 4.400 49.280 225.600 49.320 ;
        RECT 4.400 47.920 226.000 49.280 ;
        RECT 0.065 45.920 226.000 47.920 ;
        RECT 4.400 44.520 226.000 45.920 ;
        RECT 0.065 43.200 226.000 44.520 ;
        RECT 4.400 41.800 226.000 43.200 ;
        RECT 0.065 40.480 226.000 41.800 ;
        RECT 4.400 39.080 226.000 40.480 ;
        RECT 0.065 37.080 226.000 39.080 ;
        RECT 4.400 35.680 226.000 37.080 ;
        RECT 0.065 34.360 226.000 35.680 ;
        RECT 4.400 32.960 226.000 34.360 ;
        RECT 0.065 31.640 226.000 32.960 ;
        RECT 4.400 30.240 226.000 31.640 ;
        RECT 0.065 28.240 226.000 30.240 ;
        RECT 4.400 26.840 226.000 28.240 ;
        RECT 0.065 25.520 226.000 26.840 ;
        RECT 4.400 24.120 226.000 25.520 ;
        RECT 0.065 22.800 226.000 24.120 ;
        RECT 4.400 21.400 226.000 22.800 ;
        RECT 0.065 19.400 226.000 21.400 ;
        RECT 4.400 18.000 226.000 19.400 ;
        RECT 0.065 16.680 226.000 18.000 ;
        RECT 4.400 15.280 226.000 16.680 ;
        RECT 0.065 13.960 226.000 15.280 ;
        RECT 4.400 12.560 226.000 13.960 ;
        RECT 0.065 10.560 226.000 12.560 ;
        RECT 4.400 9.160 226.000 10.560 ;
        RECT 0.065 7.840 226.000 9.160 ;
        RECT 4.400 6.440 226.000 7.840 ;
        RECT 0.065 5.120 226.000 6.440 ;
        RECT 4.400 3.720 226.000 5.120 ;
        RECT 0.065 2.400 226.000 3.720 ;
        RECT 4.400 1.000 226.000 2.400 ;
        RECT 0.065 0.175 226.000 1.000 ;
      LAYER met4 ;
        RECT 3.975 188.320 169.905 189.545 ;
        RECT 3.975 10.240 20.640 188.320 ;
        RECT 23.040 10.240 97.440 188.320 ;
        RECT 99.840 10.240 169.905 188.320 ;
        RECT 3.975 0.175 169.905 10.240 ;
  END
END IOMultiplexer
END LIBRARY

