VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CaravelHost
  CLASS BLOCK ;
  FOREIGN CaravelHost ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 425.000 ;
  PIN caravel_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 421.000 385.850 425.000 ;
    END
  END caravel_irq[0]
  PIN caravel_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 421.000 389.530 425.000 ;
    END
  END caravel_irq[1]
  PIN caravel_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 421.000 393.210 425.000 ;
    END
  END caravel_irq[2]
  PIN caravel_irq[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 421.000 396.890 425.000 ;
    END
  END caravel_irq[3]
  PIN caravel_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 421.000 378.490 425.000 ;
    END
  END caravel_uart_rx
  PIN caravel_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 421.000 382.170 425.000 ;
    END
  END caravel_uart_tx
  PIN caravel_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 421.000 3.130 425.000 ;
    END
  END caravel_wb_ack_i
  PIN caravel_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 421.000 25.210 425.000 ;
    END
  END caravel_wb_adr_o[0]
  PIN caravel_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 421.000 150.330 425.000 ;
    END
  END caravel_wb_adr_o[10]
  PIN caravel_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 421.000 161.370 425.000 ;
    END
  END caravel_wb_adr_o[11]
  PIN caravel_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 421.000 172.410 425.000 ;
    END
  END caravel_wb_adr_o[12]
  PIN caravel_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 421.000 183.450 425.000 ;
    END
  END caravel_wb_adr_o[13]
  PIN caravel_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 421.000 194.490 425.000 ;
    END
  END caravel_wb_adr_o[14]
  PIN caravel_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 421.000 205.530 425.000 ;
    END
  END caravel_wb_adr_o[15]
  PIN caravel_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 421.000 216.570 425.000 ;
    END
  END caravel_wb_adr_o[16]
  PIN caravel_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 421.000 227.610 425.000 ;
    END
  END caravel_wb_adr_o[17]
  PIN caravel_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 421.000 238.650 425.000 ;
    END
  END caravel_wb_adr_o[18]
  PIN caravel_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 421.000 249.690 425.000 ;
    END
  END caravel_wb_adr_o[19]
  PIN caravel_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 421.000 39.930 425.000 ;
    END
  END caravel_wb_adr_o[1]
  PIN caravel_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 421.000 260.730 425.000 ;
    END
  END caravel_wb_adr_o[20]
  PIN caravel_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 421.000 271.770 425.000 ;
    END
  END caravel_wb_adr_o[21]
  PIN caravel_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 421.000 282.810 425.000 ;
    END
  END caravel_wb_adr_o[22]
  PIN caravel_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 421.000 293.850 425.000 ;
    END
  END caravel_wb_adr_o[23]
  PIN caravel_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 421.000 304.890 425.000 ;
    END
  END caravel_wb_adr_o[24]
  PIN caravel_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 421.000 315.930 425.000 ;
    END
  END caravel_wb_adr_o[25]
  PIN caravel_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 421.000 326.970 425.000 ;
    END
  END caravel_wb_adr_o[26]
  PIN caravel_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 421.000 338.010 425.000 ;
    END
  END caravel_wb_adr_o[27]
  PIN caravel_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 421.000 54.650 425.000 ;
    END
  END caravel_wb_adr_o[2]
  PIN caravel_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 421.000 69.370 425.000 ;
    END
  END caravel_wb_adr_o[3]
  PIN caravel_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 421.000 84.090 425.000 ;
    END
  END caravel_wb_adr_o[4]
  PIN caravel_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 421.000 95.130 425.000 ;
    END
  END caravel_wb_adr_o[5]
  PIN caravel_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 421.000 106.170 425.000 ;
    END
  END caravel_wb_adr_o[6]
  PIN caravel_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 421.000 117.210 425.000 ;
    END
  END caravel_wb_adr_o[7]
  PIN caravel_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 421.000 128.250 425.000 ;
    END
  END caravel_wb_adr_o[8]
  PIN caravel_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 421.000 139.290 425.000 ;
    END
  END caravel_wb_adr_o[9]
  PIN caravel_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 421.000 6.810 425.000 ;
    END
  END caravel_wb_cyc_o
  PIN caravel_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 421.000 28.890 425.000 ;
    END
  END caravel_wb_data_i[0]
  PIN caravel_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 421.000 154.010 425.000 ;
    END
  END caravel_wb_data_i[10]
  PIN caravel_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 421.000 165.050 425.000 ;
    END
  END caravel_wb_data_i[11]
  PIN caravel_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 421.000 176.090 425.000 ;
    END
  END caravel_wb_data_i[12]
  PIN caravel_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 421.000 187.130 425.000 ;
    END
  END caravel_wb_data_i[13]
  PIN caravel_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 421.000 198.170 425.000 ;
    END
  END caravel_wb_data_i[14]
  PIN caravel_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 421.000 209.210 425.000 ;
    END
  END caravel_wb_data_i[15]
  PIN caravel_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 421.000 220.250 425.000 ;
    END
  END caravel_wb_data_i[16]
  PIN caravel_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 421.000 231.290 425.000 ;
    END
  END caravel_wb_data_i[17]
  PIN caravel_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 421.000 242.330 425.000 ;
    END
  END caravel_wb_data_i[18]
  PIN caravel_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 421.000 253.370 425.000 ;
    END
  END caravel_wb_data_i[19]
  PIN caravel_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 421.000 43.610 425.000 ;
    END
  END caravel_wb_data_i[1]
  PIN caravel_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 421.000 264.410 425.000 ;
    END
  END caravel_wb_data_i[20]
  PIN caravel_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 421.000 275.450 425.000 ;
    END
  END caravel_wb_data_i[21]
  PIN caravel_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 421.000 286.490 425.000 ;
    END
  END caravel_wb_data_i[22]
  PIN caravel_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 421.000 297.530 425.000 ;
    END
  END caravel_wb_data_i[23]
  PIN caravel_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 421.000 308.570 425.000 ;
    END
  END caravel_wb_data_i[24]
  PIN caravel_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 421.000 319.610 425.000 ;
    END
  END caravel_wb_data_i[25]
  PIN caravel_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 421.000 330.650 425.000 ;
    END
  END caravel_wb_data_i[26]
  PIN caravel_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 421.000 341.690 425.000 ;
    END
  END caravel_wb_data_i[27]
  PIN caravel_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 421.000 349.050 425.000 ;
    END
  END caravel_wb_data_i[28]
  PIN caravel_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 421.000 356.410 425.000 ;
    END
  END caravel_wb_data_i[29]
  PIN caravel_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 421.000 58.330 425.000 ;
    END
  END caravel_wb_data_i[2]
  PIN caravel_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 421.000 363.770 425.000 ;
    END
  END caravel_wb_data_i[30]
  PIN caravel_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 421.000 371.130 425.000 ;
    END
  END caravel_wb_data_i[31]
  PIN caravel_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 421.000 73.050 425.000 ;
    END
  END caravel_wb_data_i[3]
  PIN caravel_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 421.000 87.770 425.000 ;
    END
  END caravel_wb_data_i[4]
  PIN caravel_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 421.000 98.810 425.000 ;
    END
  END caravel_wb_data_i[5]
  PIN caravel_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 421.000 109.850 425.000 ;
    END
  END caravel_wb_data_i[6]
  PIN caravel_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 421.000 120.890 425.000 ;
    END
  END caravel_wb_data_i[7]
  PIN caravel_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 421.000 131.930 425.000 ;
    END
  END caravel_wb_data_i[8]
  PIN caravel_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 421.000 142.970 425.000 ;
    END
  END caravel_wb_data_i[9]
  PIN caravel_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 421.000 32.570 425.000 ;
    END
  END caravel_wb_data_o[0]
  PIN caravel_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 421.000 157.690 425.000 ;
    END
  END caravel_wb_data_o[10]
  PIN caravel_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 421.000 168.730 425.000 ;
    END
  END caravel_wb_data_o[11]
  PIN caravel_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 421.000 179.770 425.000 ;
    END
  END caravel_wb_data_o[12]
  PIN caravel_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 421.000 190.810 425.000 ;
    END
  END caravel_wb_data_o[13]
  PIN caravel_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 421.000 201.850 425.000 ;
    END
  END caravel_wb_data_o[14]
  PIN caravel_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 421.000 212.890 425.000 ;
    END
  END caravel_wb_data_o[15]
  PIN caravel_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 421.000 223.930 425.000 ;
    END
  END caravel_wb_data_o[16]
  PIN caravel_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 421.000 234.970 425.000 ;
    END
  END caravel_wb_data_o[17]
  PIN caravel_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 421.000 246.010 425.000 ;
    END
  END caravel_wb_data_o[18]
  PIN caravel_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 421.000 257.050 425.000 ;
    END
  END caravel_wb_data_o[19]
  PIN caravel_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 421.000 47.290 425.000 ;
    END
  END caravel_wb_data_o[1]
  PIN caravel_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 421.000 268.090 425.000 ;
    END
  END caravel_wb_data_o[20]
  PIN caravel_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 421.000 279.130 425.000 ;
    END
  END caravel_wb_data_o[21]
  PIN caravel_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 421.000 290.170 425.000 ;
    END
  END caravel_wb_data_o[22]
  PIN caravel_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 421.000 301.210 425.000 ;
    END
  END caravel_wb_data_o[23]
  PIN caravel_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 421.000 312.250 425.000 ;
    END
  END caravel_wb_data_o[24]
  PIN caravel_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 421.000 323.290 425.000 ;
    END
  END caravel_wb_data_o[25]
  PIN caravel_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 421.000 334.330 425.000 ;
    END
  END caravel_wb_data_o[26]
  PIN caravel_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 421.000 345.370 425.000 ;
    END
  END caravel_wb_data_o[27]
  PIN caravel_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 421.000 352.730 425.000 ;
    END
  END caravel_wb_data_o[28]
  PIN caravel_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 421.000 360.090 425.000 ;
    END
  END caravel_wb_data_o[29]
  PIN caravel_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 421.000 62.010 425.000 ;
    END
  END caravel_wb_data_o[2]
  PIN caravel_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 421.000 367.450 425.000 ;
    END
  END caravel_wb_data_o[30]
  PIN caravel_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 421.000 374.810 425.000 ;
    END
  END caravel_wb_data_o[31]
  PIN caravel_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 421.000 76.730 425.000 ;
    END
  END caravel_wb_data_o[3]
  PIN caravel_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 421.000 91.450 425.000 ;
    END
  END caravel_wb_data_o[4]
  PIN caravel_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 421.000 102.490 425.000 ;
    END
  END caravel_wb_data_o[5]
  PIN caravel_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 421.000 113.530 425.000 ;
    END
  END caravel_wb_data_o[6]
  PIN caravel_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 421.000 124.570 425.000 ;
    END
  END caravel_wb_data_o[7]
  PIN caravel_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 421.000 135.610 425.000 ;
    END
  END caravel_wb_data_o[8]
  PIN caravel_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 421.000 146.650 425.000 ;
    END
  END caravel_wb_data_o[9]
  PIN caravel_wb_error_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 421.000 10.490 425.000 ;
    END
  END caravel_wb_error_i
  PIN caravel_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 421.000 36.250 425.000 ;
    END
  END caravel_wb_sel_o[0]
  PIN caravel_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 421.000 50.970 425.000 ;
    END
  END caravel_wb_sel_o[1]
  PIN caravel_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 421.000 65.690 425.000 ;
    END
  END caravel_wb_sel_o[2]
  PIN caravel_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 421.000 80.410 425.000 ;
    END
  END caravel_wb_sel_o[3]
  PIN caravel_wb_stall_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 421.000 14.170 425.000 ;
    END
  END caravel_wb_stall_i
  PIN caravel_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 421.000 17.850 425.000 ;
    END
  END caravel_wb_stb_o
  PIN caravel_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 421.000 21.530 425.000 ;
    END
  END caravel_wb_we_o
  PIN core0Index[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END core0Index[0]
  PIN core0Index[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END core0Index[1]
  PIN core0Index[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END core0Index[2]
  PIN core0Index[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END core0Index[3]
  PIN core0Index[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END core0Index[4]
  PIN core0Index[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END core0Index[5]
  PIN core0Index[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END core0Index[6]
  PIN core0Index[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END core0Index[7]
  PIN core1Index[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END core1Index[0]
  PIN core1Index[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END core1Index[1]
  PIN core1Index[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END core1Index[2]
  PIN core1Index[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END core1Index[3]
  PIN core1Index[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END core1Index[4]
  PIN core1Index[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END core1Index[5]
  PIN core1Index[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END core1Index[6]
  PIN core1Index[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END core1Index[7]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 59.200 400.000 59.800 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 195.200 400.000 195.800 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 196.560 400.000 197.160 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.920 400.000 198.520 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 199.280 400.000 199.880 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 200.640 400.000 201.240 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 202.000 400.000 202.600 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 203.360 400.000 203.960 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.720 400.000 205.320 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 206.080 400.000 206.680 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 207.440 400.000 208.040 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 72.800 400.000 73.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 208.800 400.000 209.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 210.160 400.000 210.760 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 211.520 400.000 212.120 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 212.880 400.000 213.480 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.240 400.000 214.840 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 215.600 400.000 216.200 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 216.960 400.000 217.560 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 218.320 400.000 218.920 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 219.680 400.000 220.280 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.040 400.000 221.640 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 74.160 400.000 74.760 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 222.400 400.000 223.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 223.760 400.000 224.360 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 225.120 400.000 225.720 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 226.480 400.000 227.080 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 227.840 400.000 228.440 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 229.200 400.000 229.800 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 230.560 400.000 231.160 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 231.920 400.000 232.520 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 75.520 400.000 76.120 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 76.880 400.000 77.480 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 78.240 400.000 78.840 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 79.600 400.000 80.200 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 80.960 400.000 81.560 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 82.320 400.000 82.920 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 83.680 400.000 84.280 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 85.040 400.000 85.640 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 60.560 400.000 61.160 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 86.400 400.000 87.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 87.760 400.000 88.360 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 89.120 400.000 89.720 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 90.480 400.000 91.080 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 91.840 400.000 92.440 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 93.200 400.000 93.800 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 94.560 400.000 95.160 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.920 400.000 96.520 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 97.280 400.000 97.880 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 98.640 400.000 99.240 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 61.920 400.000 62.520 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 100.000 400.000 100.600 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 101.360 400.000 101.960 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 102.720 400.000 103.320 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 104.080 400.000 104.680 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 105.440 400.000 106.040 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 106.800 400.000 107.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 108.160 400.000 108.760 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 109.520 400.000 110.120 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 110.880 400.000 111.480 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.240 400.000 112.840 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 63.280 400.000 63.880 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 113.600 400.000 114.200 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 114.960 400.000 115.560 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 116.320 400.000 116.920 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 117.680 400.000 118.280 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 119.040 400.000 119.640 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 120.400 400.000 121.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 121.760 400.000 122.360 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 123.120 400.000 123.720 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 124.480 400.000 125.080 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 125.840 400.000 126.440 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 64.640 400.000 65.240 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 127.200 400.000 127.800 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 128.560 400.000 129.160 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 129.920 400.000 130.520 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 131.280 400.000 131.880 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 132.640 400.000 133.240 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 134.000 400.000 134.600 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 135.360 400.000 135.960 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 136.720 400.000 137.320 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 138.080 400.000 138.680 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 139.440 400.000 140.040 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 66.000 400.000 66.600 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 140.800 400.000 141.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 142.160 400.000 142.760 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 143.520 400.000 144.120 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 144.880 400.000 145.480 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 146.240 400.000 146.840 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 147.600 400.000 148.200 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 148.960 400.000 149.560 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 150.320 400.000 150.920 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 151.680 400.000 152.280 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 153.040 400.000 153.640 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 67.360 400.000 67.960 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 154.400 400.000 155.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 155.760 400.000 156.360 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 157.120 400.000 157.720 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 158.480 400.000 159.080 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 159.840 400.000 160.440 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 161.200 400.000 161.800 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 162.560 400.000 163.160 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 163.920 400.000 164.520 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 165.280 400.000 165.880 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 166.640 400.000 167.240 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.720 400.000 69.320 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 168.000 400.000 168.600 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 169.360 400.000 169.960 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.720 400.000 171.320 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 172.080 400.000 172.680 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 173.440 400.000 174.040 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 174.800 400.000 175.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 176.160 400.000 176.760 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 177.520 400.000 178.120 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 178.880 400.000 179.480 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.240 400.000 180.840 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 70.080 400.000 70.680 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 181.600 400.000 182.200 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 182.960 400.000 183.560 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 184.320 400.000 184.920 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 185.680 400.000 186.280 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 187.040 400.000 187.640 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 188.400 400.000 189.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 189.760 400.000 190.360 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 191.120 400.000 191.720 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 192.480 400.000 193.080 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.840 400.000 194.440 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 71.440 400.000 72.040 ;
    END
  END la_data_out[9]
  PIN manufacturerID[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END partID[9]
  PIN probe_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 233.280 400.000 233.880 ;
    END
  END probe_out[0]
  PIN probe_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 246.880 400.000 247.480 ;
    END
  END probe_out[10]
  PIN probe_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 248.240 400.000 248.840 ;
    END
  END probe_out[11]
  PIN probe_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 249.600 400.000 250.200 ;
    END
  END probe_out[12]
  PIN probe_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 250.960 400.000 251.560 ;
    END
  END probe_out[13]
  PIN probe_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 252.320 400.000 252.920 ;
    END
  END probe_out[14]
  PIN probe_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 253.680 400.000 254.280 ;
    END
  END probe_out[15]
  PIN probe_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 255.040 400.000 255.640 ;
    END
  END probe_out[16]
  PIN probe_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 256.400 400.000 257.000 ;
    END
  END probe_out[17]
  PIN probe_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 257.760 400.000 258.360 ;
    END
  END probe_out[18]
  PIN probe_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 259.120 400.000 259.720 ;
    END
  END probe_out[19]
  PIN probe_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 234.640 400.000 235.240 ;
    END
  END probe_out[1]
  PIN probe_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 260.480 400.000 261.080 ;
    END
  END probe_out[20]
  PIN probe_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 261.840 400.000 262.440 ;
    END
  END probe_out[21]
  PIN probe_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 263.200 400.000 263.800 ;
    END
  END probe_out[22]
  PIN probe_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 264.560 400.000 265.160 ;
    END
  END probe_out[23]
  PIN probe_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 265.920 400.000 266.520 ;
    END
  END probe_out[24]
  PIN probe_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 267.280 400.000 267.880 ;
    END
  END probe_out[25]
  PIN probe_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 268.640 400.000 269.240 ;
    END
  END probe_out[26]
  PIN probe_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 270.000 400.000 270.600 ;
    END
  END probe_out[27]
  PIN probe_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 271.360 400.000 271.960 ;
    END
  END probe_out[28]
  PIN probe_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 272.720 400.000 273.320 ;
    END
  END probe_out[29]
  PIN probe_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 236.000 400.000 236.600 ;
    END
  END probe_out[2]
  PIN probe_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 274.080 400.000 274.680 ;
    END
  END probe_out[30]
  PIN probe_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 275.440 400.000 276.040 ;
    END
  END probe_out[31]
  PIN probe_out[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 276.800 400.000 277.400 ;
    END
  END probe_out[32]
  PIN probe_out[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.160 400.000 278.760 ;
    END
  END probe_out[33]
  PIN probe_out[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 279.520 400.000 280.120 ;
    END
  END probe_out[34]
  PIN probe_out[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 280.880 400.000 281.480 ;
    END
  END probe_out[35]
  PIN probe_out[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 282.240 400.000 282.840 ;
    END
  END probe_out[36]
  PIN probe_out[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 283.600 400.000 284.200 ;
    END
  END probe_out[37]
  PIN probe_out[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 284.960 400.000 285.560 ;
    END
  END probe_out[38]
  PIN probe_out[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 286.320 400.000 286.920 ;
    END
  END probe_out[39]
  PIN probe_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 237.360 400.000 237.960 ;
    END
  END probe_out[3]
  PIN probe_out[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 287.680 400.000 288.280 ;
    END
  END probe_out[40]
  PIN probe_out[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 289.040 400.000 289.640 ;
    END
  END probe_out[41]
  PIN probe_out[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 290.400 400.000 291.000 ;
    END
  END probe_out[42]
  PIN probe_out[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 291.760 400.000 292.360 ;
    END
  END probe_out[43]
  PIN probe_out[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 293.120 400.000 293.720 ;
    END
  END probe_out[44]
  PIN probe_out[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 294.480 400.000 295.080 ;
    END
  END probe_out[45]
  PIN probe_out[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 295.840 400.000 296.440 ;
    END
  END probe_out[46]
  PIN probe_out[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 297.200 400.000 297.800 ;
    END
  END probe_out[47]
  PIN probe_out[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 298.560 400.000 299.160 ;
    END
  END probe_out[48]
  PIN probe_out[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 299.920 400.000 300.520 ;
    END
  END probe_out[49]
  PIN probe_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.720 400.000 239.320 ;
    END
  END probe_out[4]
  PIN probe_out[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 301.280 400.000 301.880 ;
    END
  END probe_out[50]
  PIN probe_out[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 302.640 400.000 303.240 ;
    END
  END probe_out[51]
  PIN probe_out[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 304.000 400.000 304.600 ;
    END
  END probe_out[52]
  PIN probe_out[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 305.360 400.000 305.960 ;
    END
  END probe_out[53]
  PIN probe_out[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.720 400.000 307.320 ;
    END
  END probe_out[54]
  PIN probe_out[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 308.080 400.000 308.680 ;
    END
  END probe_out[55]
  PIN probe_out[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 309.440 400.000 310.040 ;
    END
  END probe_out[56]
  PIN probe_out[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 310.800 400.000 311.400 ;
    END
  END probe_out[57]
  PIN probe_out[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 312.160 400.000 312.760 ;
    END
  END probe_out[58]
  PIN probe_out[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 313.520 400.000 314.120 ;
    END
  END probe_out[59]
  PIN probe_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 240.080 400.000 240.680 ;
    END
  END probe_out[5]
  PIN probe_out[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 314.880 400.000 315.480 ;
    END
  END probe_out[60]
  PIN probe_out[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 316.240 400.000 316.840 ;
    END
  END probe_out[61]
  PIN probe_out[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 317.600 400.000 318.200 ;
    END
  END probe_out[62]
  PIN probe_out[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 318.960 400.000 319.560 ;
    END
  END probe_out[63]
  PIN probe_out[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 320.320 400.000 320.920 ;
    END
  END probe_out[64]
  PIN probe_out[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 321.680 400.000 322.280 ;
    END
  END probe_out[65]
  PIN probe_out[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 323.040 400.000 323.640 ;
    END
  END probe_out[66]
  PIN probe_out[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 324.400 400.000 325.000 ;
    END
  END probe_out[67]
  PIN probe_out[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 325.760 400.000 326.360 ;
    END
  END probe_out[68]
  PIN probe_out[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 327.120 400.000 327.720 ;
    END
  END probe_out[69]
  PIN probe_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 241.440 400.000 242.040 ;
    END
  END probe_out[6]
  PIN probe_out[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 328.480 400.000 329.080 ;
    END
  END probe_out[70]
  PIN probe_out[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 329.840 400.000 330.440 ;
    END
  END probe_out[71]
  PIN probe_out[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 331.200 400.000 331.800 ;
    END
  END probe_out[72]
  PIN probe_out[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 332.560 400.000 333.160 ;
    END
  END probe_out[73]
  PIN probe_out[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.920 400.000 334.520 ;
    END
  END probe_out[74]
  PIN probe_out[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 335.280 400.000 335.880 ;
    END
  END probe_out[75]
  PIN probe_out[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 336.640 400.000 337.240 ;
    END
  END probe_out[76]
  PIN probe_out[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 338.000 400.000 338.600 ;
    END
  END probe_out[77]
  PIN probe_out[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 339.360 400.000 339.960 ;
    END
  END probe_out[78]
  PIN probe_out[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 340.720 400.000 341.320 ;
    END
  END probe_out[79]
  PIN probe_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 242.800 400.000 243.400 ;
    END
  END probe_out[7]
  PIN probe_out[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 342.080 400.000 342.680 ;
    END
  END probe_out[80]
  PIN probe_out[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 343.440 400.000 344.040 ;
    END
  END probe_out[81]
  PIN probe_out[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 344.800 400.000 345.400 ;
    END
  END probe_out[82]
  PIN probe_out[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 346.160 400.000 346.760 ;
    END
  END probe_out[83]
  PIN probe_out[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 347.520 400.000 348.120 ;
    END
  END probe_out[84]
  PIN probe_out[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 348.880 400.000 349.480 ;
    END
  END probe_out[85]
  PIN probe_out[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 350.240 400.000 350.840 ;
    END
  END probe_out[86]
  PIN probe_out[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 351.600 400.000 352.200 ;
    END
  END probe_out[87]
  PIN probe_out[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 352.960 400.000 353.560 ;
    END
  END probe_out[88]
  PIN probe_out[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 354.320 400.000 354.920 ;
    END
  END probe_out[89]
  PIN probe_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 244.160 400.000 244.760 ;
    END
  END probe_out[8]
  PIN probe_out[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 355.680 400.000 356.280 ;
    END
  END probe_out[90]
  PIN probe_out[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 357.040 400.000 357.640 ;
    END
  END probe_out[91]
  PIN probe_out[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 358.400 400.000 359.000 ;
    END
  END probe_out[92]
  PIN probe_out[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 359.760 400.000 360.360 ;
    END
  END probe_out[93]
  PIN probe_out[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 361.120 400.000 361.720 ;
    END
  END probe_out[94]
  PIN probe_out[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 362.480 400.000 363.080 ;
    END
  END probe_out[95]
  PIN probe_out[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 363.840 400.000 364.440 ;
    END
  END probe_out[96]
  PIN probe_out[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 365.200 400.000 365.800 ;
    END
  END probe_out[97]
  PIN probe_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 245.520 400.000 246.120 ;
    END
  END probe_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 413.680 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 413.680 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wbs_data_i[0]
  PIN wbs_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END wbs_data_i[10]
  PIN wbs_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_data_i[11]
  PIN wbs_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wbs_data_i[12]
  PIN wbs_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END wbs_data_i[13]
  PIN wbs_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END wbs_data_i[14]
  PIN wbs_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wbs_data_i[15]
  PIN wbs_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END wbs_data_i[16]
  PIN wbs_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END wbs_data_i[17]
  PIN wbs_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END wbs_data_i[18]
  PIN wbs_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END wbs_data_i[19]
  PIN wbs_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END wbs_data_i[1]
  PIN wbs_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END wbs_data_i[20]
  PIN wbs_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END wbs_data_i[21]
  PIN wbs_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END wbs_data_i[22]
  PIN wbs_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END wbs_data_i[23]
  PIN wbs_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END wbs_data_i[24]
  PIN wbs_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END wbs_data_i[25]
  PIN wbs_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_data_i[26]
  PIN wbs_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END wbs_data_i[27]
  PIN wbs_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END wbs_data_i[28]
  PIN wbs_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END wbs_data_i[29]
  PIN wbs_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_data_i[2]
  PIN wbs_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END wbs_data_i[30]
  PIN wbs_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END wbs_data_i[31]
  PIN wbs_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END wbs_data_i[3]
  PIN wbs_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END wbs_data_i[4]
  PIN wbs_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_data_i[5]
  PIN wbs_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END wbs_data_i[6]
  PIN wbs_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_data_i[7]
  PIN wbs_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_data_i[8]
  PIN wbs_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END wbs_data_i[9]
  PIN wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END wbs_data_o[0]
  PIN wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END wbs_data_o[10]
  PIN wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END wbs_data_o[11]
  PIN wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END wbs_data_o[12]
  PIN wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END wbs_data_o[13]
  PIN wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END wbs_data_o[14]
  PIN wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END wbs_data_o[15]
  PIN wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END wbs_data_o[16]
  PIN wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END wbs_data_o[17]
  PIN wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END wbs_data_o[18]
  PIN wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END wbs_data_o[19]
  PIN wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END wbs_data_o[1]
  PIN wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END wbs_data_o[20]
  PIN wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END wbs_data_o[21]
  PIN wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_data_o[22]
  PIN wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END wbs_data_o[23]
  PIN wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END wbs_data_o[24]
  PIN wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END wbs_data_o[25]
  PIN wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END wbs_data_o[26]
  PIN wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END wbs_data_o[27]
  PIN wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END wbs_data_o[28]
  PIN wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END wbs_data_o[29]
  PIN wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END wbs_data_o[2]
  PIN wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END wbs_data_o[30]
  PIN wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END wbs_data_o[31]
  PIN wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END wbs_data_o[3]
  PIN wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END wbs_data_o[4]
  PIN wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END wbs_data_o[5]
  PIN wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_data_o[6]
  PIN wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_data_o[7]
  PIN wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wbs_data_o[8]
  PIN wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END wbs_data_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 413.525 ;
      LAYER met1 ;
        RECT 2.830 0.380 399.670 420.540 ;
      LAYER met2 ;
        RECT 3.410 420.720 6.250 421.330 ;
        RECT 7.090 420.720 9.930 421.330 ;
        RECT 10.770 420.720 13.610 421.330 ;
        RECT 14.450 420.720 17.290 421.330 ;
        RECT 18.130 420.720 20.970 421.330 ;
        RECT 21.810 420.720 24.650 421.330 ;
        RECT 25.490 420.720 28.330 421.330 ;
        RECT 29.170 420.720 32.010 421.330 ;
        RECT 32.850 420.720 35.690 421.330 ;
        RECT 36.530 420.720 39.370 421.330 ;
        RECT 40.210 420.720 43.050 421.330 ;
        RECT 43.890 420.720 46.730 421.330 ;
        RECT 47.570 420.720 50.410 421.330 ;
        RECT 51.250 420.720 54.090 421.330 ;
        RECT 54.930 420.720 57.770 421.330 ;
        RECT 58.610 420.720 61.450 421.330 ;
        RECT 62.290 420.720 65.130 421.330 ;
        RECT 65.970 420.720 68.810 421.330 ;
        RECT 69.650 420.720 72.490 421.330 ;
        RECT 73.330 420.720 76.170 421.330 ;
        RECT 77.010 420.720 79.850 421.330 ;
        RECT 80.690 420.720 83.530 421.330 ;
        RECT 84.370 420.720 87.210 421.330 ;
        RECT 88.050 420.720 90.890 421.330 ;
        RECT 91.730 420.720 94.570 421.330 ;
        RECT 95.410 420.720 98.250 421.330 ;
        RECT 99.090 420.720 101.930 421.330 ;
        RECT 102.770 420.720 105.610 421.330 ;
        RECT 106.450 420.720 109.290 421.330 ;
        RECT 110.130 420.720 112.970 421.330 ;
        RECT 113.810 420.720 116.650 421.330 ;
        RECT 117.490 420.720 120.330 421.330 ;
        RECT 121.170 420.720 124.010 421.330 ;
        RECT 124.850 420.720 127.690 421.330 ;
        RECT 128.530 420.720 131.370 421.330 ;
        RECT 132.210 420.720 135.050 421.330 ;
        RECT 135.890 420.720 138.730 421.330 ;
        RECT 139.570 420.720 142.410 421.330 ;
        RECT 143.250 420.720 146.090 421.330 ;
        RECT 146.930 420.720 149.770 421.330 ;
        RECT 150.610 420.720 153.450 421.330 ;
        RECT 154.290 420.720 157.130 421.330 ;
        RECT 157.970 420.720 160.810 421.330 ;
        RECT 161.650 420.720 164.490 421.330 ;
        RECT 165.330 420.720 168.170 421.330 ;
        RECT 169.010 420.720 171.850 421.330 ;
        RECT 172.690 420.720 175.530 421.330 ;
        RECT 176.370 420.720 179.210 421.330 ;
        RECT 180.050 420.720 182.890 421.330 ;
        RECT 183.730 420.720 186.570 421.330 ;
        RECT 187.410 420.720 190.250 421.330 ;
        RECT 191.090 420.720 193.930 421.330 ;
        RECT 194.770 420.720 197.610 421.330 ;
        RECT 198.450 420.720 201.290 421.330 ;
        RECT 202.130 420.720 204.970 421.330 ;
        RECT 205.810 420.720 208.650 421.330 ;
        RECT 209.490 420.720 212.330 421.330 ;
        RECT 213.170 420.720 216.010 421.330 ;
        RECT 216.850 420.720 219.690 421.330 ;
        RECT 220.530 420.720 223.370 421.330 ;
        RECT 224.210 420.720 227.050 421.330 ;
        RECT 227.890 420.720 230.730 421.330 ;
        RECT 231.570 420.720 234.410 421.330 ;
        RECT 235.250 420.720 238.090 421.330 ;
        RECT 238.930 420.720 241.770 421.330 ;
        RECT 242.610 420.720 245.450 421.330 ;
        RECT 246.290 420.720 249.130 421.330 ;
        RECT 249.970 420.720 252.810 421.330 ;
        RECT 253.650 420.720 256.490 421.330 ;
        RECT 257.330 420.720 260.170 421.330 ;
        RECT 261.010 420.720 263.850 421.330 ;
        RECT 264.690 420.720 267.530 421.330 ;
        RECT 268.370 420.720 271.210 421.330 ;
        RECT 272.050 420.720 274.890 421.330 ;
        RECT 275.730 420.720 278.570 421.330 ;
        RECT 279.410 420.720 282.250 421.330 ;
        RECT 283.090 420.720 285.930 421.330 ;
        RECT 286.770 420.720 289.610 421.330 ;
        RECT 290.450 420.720 293.290 421.330 ;
        RECT 294.130 420.720 296.970 421.330 ;
        RECT 297.810 420.720 300.650 421.330 ;
        RECT 301.490 420.720 304.330 421.330 ;
        RECT 305.170 420.720 308.010 421.330 ;
        RECT 308.850 420.720 311.690 421.330 ;
        RECT 312.530 420.720 315.370 421.330 ;
        RECT 316.210 420.720 319.050 421.330 ;
        RECT 319.890 420.720 322.730 421.330 ;
        RECT 323.570 420.720 326.410 421.330 ;
        RECT 327.250 420.720 330.090 421.330 ;
        RECT 330.930 420.720 333.770 421.330 ;
        RECT 334.610 420.720 337.450 421.330 ;
        RECT 338.290 420.720 341.130 421.330 ;
        RECT 341.970 420.720 344.810 421.330 ;
        RECT 345.650 420.720 348.490 421.330 ;
        RECT 349.330 420.720 352.170 421.330 ;
        RECT 353.010 420.720 355.850 421.330 ;
        RECT 356.690 420.720 359.530 421.330 ;
        RECT 360.370 420.720 363.210 421.330 ;
        RECT 364.050 420.720 366.890 421.330 ;
        RECT 367.730 420.720 370.570 421.330 ;
        RECT 371.410 420.720 374.250 421.330 ;
        RECT 375.090 420.720 377.930 421.330 ;
        RECT 378.770 420.720 381.610 421.330 ;
        RECT 382.450 420.720 385.290 421.330 ;
        RECT 386.130 420.720 388.970 421.330 ;
        RECT 389.810 420.720 392.650 421.330 ;
        RECT 393.490 420.720 396.330 421.330 ;
        RECT 397.170 420.720 399.640 421.330 ;
        RECT 2.860 4.280 399.640 420.720 ;
        RECT 2.860 0.350 6.250 4.280 ;
        RECT 7.090 0.350 9.930 4.280 ;
        RECT 10.770 0.350 13.610 4.280 ;
        RECT 14.450 0.350 17.290 4.280 ;
        RECT 18.130 0.350 20.970 4.280 ;
        RECT 21.810 0.350 24.650 4.280 ;
        RECT 25.490 0.350 28.330 4.280 ;
        RECT 29.170 0.350 32.010 4.280 ;
        RECT 32.850 0.350 35.690 4.280 ;
        RECT 36.530 0.350 39.370 4.280 ;
        RECT 40.210 0.350 43.050 4.280 ;
        RECT 43.890 0.350 46.730 4.280 ;
        RECT 47.570 0.350 50.410 4.280 ;
        RECT 51.250 0.350 54.090 4.280 ;
        RECT 54.930 0.350 57.770 4.280 ;
        RECT 58.610 0.350 61.450 4.280 ;
        RECT 62.290 0.350 65.130 4.280 ;
        RECT 65.970 0.350 68.810 4.280 ;
        RECT 69.650 0.350 72.490 4.280 ;
        RECT 73.330 0.350 76.170 4.280 ;
        RECT 77.010 0.350 79.850 4.280 ;
        RECT 80.690 0.350 83.530 4.280 ;
        RECT 84.370 0.350 87.210 4.280 ;
        RECT 88.050 0.350 90.890 4.280 ;
        RECT 91.730 0.350 94.570 4.280 ;
        RECT 95.410 0.350 98.250 4.280 ;
        RECT 99.090 0.350 101.930 4.280 ;
        RECT 102.770 0.350 105.610 4.280 ;
        RECT 106.450 0.350 109.290 4.280 ;
        RECT 110.130 0.350 112.970 4.280 ;
        RECT 113.810 0.350 116.650 4.280 ;
        RECT 117.490 0.350 120.330 4.280 ;
        RECT 121.170 0.350 124.010 4.280 ;
        RECT 124.850 0.350 127.690 4.280 ;
        RECT 128.530 0.350 131.370 4.280 ;
        RECT 132.210 0.350 135.050 4.280 ;
        RECT 135.890 0.350 138.730 4.280 ;
        RECT 139.570 0.350 142.410 4.280 ;
        RECT 143.250 0.350 146.090 4.280 ;
        RECT 146.930 0.350 149.770 4.280 ;
        RECT 150.610 0.350 153.450 4.280 ;
        RECT 154.290 0.350 157.130 4.280 ;
        RECT 157.970 0.350 160.810 4.280 ;
        RECT 161.650 0.350 164.490 4.280 ;
        RECT 165.330 0.350 168.170 4.280 ;
        RECT 169.010 0.350 171.850 4.280 ;
        RECT 172.690 0.350 175.530 4.280 ;
        RECT 176.370 0.350 179.210 4.280 ;
        RECT 180.050 0.350 182.890 4.280 ;
        RECT 183.730 0.350 186.570 4.280 ;
        RECT 187.410 0.350 190.250 4.280 ;
        RECT 191.090 0.350 193.930 4.280 ;
        RECT 194.770 0.350 197.610 4.280 ;
        RECT 198.450 0.350 201.290 4.280 ;
        RECT 202.130 0.350 204.970 4.280 ;
        RECT 205.810 0.350 208.650 4.280 ;
        RECT 209.490 0.350 212.330 4.280 ;
        RECT 213.170 0.350 216.010 4.280 ;
        RECT 216.850 0.350 219.690 4.280 ;
        RECT 220.530 0.350 223.370 4.280 ;
        RECT 224.210 0.350 227.050 4.280 ;
        RECT 227.890 0.350 230.730 4.280 ;
        RECT 231.570 0.350 234.410 4.280 ;
        RECT 235.250 0.350 238.090 4.280 ;
        RECT 238.930 0.350 241.770 4.280 ;
        RECT 242.610 0.350 245.450 4.280 ;
        RECT 246.290 0.350 249.130 4.280 ;
        RECT 249.970 0.350 252.810 4.280 ;
        RECT 253.650 0.350 256.490 4.280 ;
        RECT 257.330 0.350 260.170 4.280 ;
        RECT 261.010 0.350 263.850 4.280 ;
        RECT 264.690 0.350 267.530 4.280 ;
        RECT 268.370 0.350 271.210 4.280 ;
        RECT 272.050 0.350 274.890 4.280 ;
        RECT 275.730 0.350 278.570 4.280 ;
        RECT 279.410 0.350 282.250 4.280 ;
        RECT 283.090 0.350 285.930 4.280 ;
        RECT 286.770 0.350 289.610 4.280 ;
        RECT 290.450 0.350 293.290 4.280 ;
        RECT 294.130 0.350 296.970 4.280 ;
        RECT 297.810 0.350 300.650 4.280 ;
        RECT 301.490 0.350 304.330 4.280 ;
        RECT 305.170 0.350 308.010 4.280 ;
        RECT 308.850 0.350 311.690 4.280 ;
        RECT 312.530 0.350 315.370 4.280 ;
        RECT 316.210 0.350 319.050 4.280 ;
        RECT 319.890 0.350 322.730 4.280 ;
        RECT 323.570 0.350 326.410 4.280 ;
        RECT 327.250 0.350 330.090 4.280 ;
        RECT 330.930 0.350 333.770 4.280 ;
        RECT 334.610 0.350 337.450 4.280 ;
        RECT 338.290 0.350 341.130 4.280 ;
        RECT 341.970 0.350 344.810 4.280 ;
        RECT 345.650 0.350 348.490 4.280 ;
        RECT 349.330 0.350 352.170 4.280 ;
        RECT 353.010 0.350 355.850 4.280 ;
        RECT 356.690 0.350 359.530 4.280 ;
        RECT 360.370 0.350 363.210 4.280 ;
        RECT 364.050 0.350 366.890 4.280 ;
        RECT 367.730 0.350 370.570 4.280 ;
        RECT 371.410 0.350 374.250 4.280 ;
        RECT 375.090 0.350 377.930 4.280 ;
        RECT 378.770 0.350 381.610 4.280 ;
        RECT 382.450 0.350 385.290 4.280 ;
        RECT 386.130 0.350 388.970 4.280 ;
        RECT 389.810 0.350 392.650 4.280 ;
        RECT 393.490 0.350 399.640 4.280 ;
      LAYER met3 ;
        RECT 4.400 415.120 396.000 415.985 ;
        RECT 4.000 407.680 396.000 415.120 ;
        RECT 4.400 406.280 396.000 407.680 ;
        RECT 4.000 398.840 396.000 406.280 ;
        RECT 4.400 397.440 396.000 398.840 ;
        RECT 4.000 390.000 396.000 397.440 ;
        RECT 4.400 388.600 396.000 390.000 ;
        RECT 4.000 381.160 396.000 388.600 ;
        RECT 4.400 379.760 396.000 381.160 ;
        RECT 4.000 372.320 396.000 379.760 ;
        RECT 4.400 370.920 396.000 372.320 ;
        RECT 4.000 366.200 396.000 370.920 ;
        RECT 4.000 363.480 395.600 366.200 ;
        RECT 4.400 362.080 395.600 363.480 ;
        RECT 4.000 354.640 395.600 362.080 ;
        RECT 4.400 353.240 395.600 354.640 ;
        RECT 4.000 345.800 395.600 353.240 ;
        RECT 4.400 344.400 395.600 345.800 ;
        RECT 4.000 336.960 395.600 344.400 ;
        RECT 4.400 335.560 395.600 336.960 ;
        RECT 4.000 328.120 395.600 335.560 ;
        RECT 4.400 326.720 395.600 328.120 ;
        RECT 4.000 319.280 395.600 326.720 ;
        RECT 4.400 317.880 395.600 319.280 ;
        RECT 4.000 310.440 395.600 317.880 ;
        RECT 4.400 309.040 395.600 310.440 ;
        RECT 4.000 301.600 395.600 309.040 ;
        RECT 4.400 300.200 395.600 301.600 ;
        RECT 4.000 292.760 395.600 300.200 ;
        RECT 4.400 291.360 395.600 292.760 ;
        RECT 4.000 283.920 395.600 291.360 ;
        RECT 4.400 282.520 395.600 283.920 ;
        RECT 4.000 275.080 395.600 282.520 ;
        RECT 4.400 273.680 395.600 275.080 ;
        RECT 4.000 266.240 395.600 273.680 ;
        RECT 4.400 264.840 395.600 266.240 ;
        RECT 4.000 257.400 395.600 264.840 ;
        RECT 4.400 256.000 395.600 257.400 ;
        RECT 4.000 248.560 395.600 256.000 ;
        RECT 4.400 247.160 395.600 248.560 ;
        RECT 4.000 239.720 395.600 247.160 ;
        RECT 4.400 238.320 395.600 239.720 ;
        RECT 4.000 230.880 395.600 238.320 ;
        RECT 4.400 229.480 395.600 230.880 ;
        RECT 4.000 222.040 395.600 229.480 ;
        RECT 4.400 220.640 395.600 222.040 ;
        RECT 4.000 213.200 395.600 220.640 ;
        RECT 4.400 211.800 395.600 213.200 ;
        RECT 4.000 204.360 395.600 211.800 ;
        RECT 4.400 202.960 395.600 204.360 ;
        RECT 4.000 195.520 395.600 202.960 ;
        RECT 4.400 194.120 395.600 195.520 ;
        RECT 4.000 186.680 395.600 194.120 ;
        RECT 4.400 185.280 395.600 186.680 ;
        RECT 4.000 177.840 395.600 185.280 ;
        RECT 4.400 176.440 395.600 177.840 ;
        RECT 4.000 169.000 395.600 176.440 ;
        RECT 4.400 167.600 395.600 169.000 ;
        RECT 4.000 160.160 395.600 167.600 ;
        RECT 4.400 158.760 395.600 160.160 ;
        RECT 4.000 151.320 395.600 158.760 ;
        RECT 4.400 149.920 395.600 151.320 ;
        RECT 4.000 142.480 395.600 149.920 ;
        RECT 4.400 141.080 395.600 142.480 ;
        RECT 4.000 133.640 395.600 141.080 ;
        RECT 4.400 132.240 395.600 133.640 ;
        RECT 4.000 124.800 395.600 132.240 ;
        RECT 4.400 123.400 395.600 124.800 ;
        RECT 4.000 115.960 395.600 123.400 ;
        RECT 4.400 114.560 395.600 115.960 ;
        RECT 4.000 107.120 395.600 114.560 ;
        RECT 4.400 105.720 395.600 107.120 ;
        RECT 4.000 98.280 395.600 105.720 ;
        RECT 4.400 96.880 395.600 98.280 ;
        RECT 4.000 89.440 395.600 96.880 ;
        RECT 4.400 88.040 395.600 89.440 ;
        RECT 4.000 80.600 395.600 88.040 ;
        RECT 4.400 79.200 395.600 80.600 ;
        RECT 4.000 71.760 395.600 79.200 ;
        RECT 4.400 70.360 395.600 71.760 ;
        RECT 4.000 62.920 395.600 70.360 ;
        RECT 4.400 61.520 395.600 62.920 ;
        RECT 4.000 58.800 395.600 61.520 ;
        RECT 4.000 54.080 396.000 58.800 ;
        RECT 4.400 52.680 396.000 54.080 ;
        RECT 4.000 45.240 396.000 52.680 ;
        RECT 4.400 43.840 396.000 45.240 ;
        RECT 4.000 36.400 396.000 43.840 ;
        RECT 4.400 35.000 396.000 36.400 ;
        RECT 4.000 27.560 396.000 35.000 ;
        RECT 4.400 26.160 396.000 27.560 ;
        RECT 4.000 18.720 396.000 26.160 ;
        RECT 4.400 17.320 396.000 18.720 ;
        RECT 4.000 9.880 396.000 17.320 ;
        RECT 4.400 9.015 396.000 9.880 ;
      LAYER met4 ;
        RECT 8.575 11.735 20.640 407.825 ;
        RECT 23.040 11.735 97.440 407.825 ;
        RECT 99.840 11.735 174.240 407.825 ;
        RECT 176.640 11.735 251.040 407.825 ;
        RECT 253.440 11.735 327.840 407.825 ;
        RECT 330.240 11.735 385.185 407.825 ;
  END
END CaravelHost
END LIBRARY

