magic
tech sky130A
magscale 1 2
timestamp 1653404051
<< obsli1 >>
rect 1104 2159 68816 217617
<< obsm1 >>
rect 290 1980 69722 217648
<< metal2 >>
rect 294 219200 350 220000
rect 938 219200 994 220000
rect 1674 219200 1730 220000
rect 2410 219200 2466 220000
rect 3146 219200 3202 220000
rect 3790 219200 3846 220000
rect 4526 219200 4582 220000
rect 5262 219200 5318 220000
rect 5998 219200 6054 220000
rect 6642 219200 6698 220000
rect 7378 219200 7434 220000
rect 8114 219200 8170 220000
rect 8850 219200 8906 220000
rect 9494 219200 9550 220000
rect 10230 219200 10286 220000
rect 10966 219200 11022 220000
rect 11702 219200 11758 220000
rect 12438 219200 12494 220000
rect 13082 219200 13138 220000
rect 13818 219200 13874 220000
rect 14554 219200 14610 220000
rect 15290 219200 15346 220000
rect 15934 219200 15990 220000
rect 16670 219200 16726 220000
rect 17406 219200 17462 220000
rect 18142 219200 18198 220000
rect 18786 219200 18842 220000
rect 19522 219200 19578 220000
rect 20258 219200 20314 220000
rect 20994 219200 21050 220000
rect 21638 219200 21694 220000
rect 22374 219200 22430 220000
rect 23110 219200 23166 220000
rect 23846 219200 23902 220000
rect 24582 219200 24638 220000
rect 25226 219200 25282 220000
rect 25962 219200 26018 220000
rect 26698 219200 26754 220000
rect 27434 219200 27490 220000
rect 28078 219200 28134 220000
rect 28814 219200 28870 220000
rect 29550 219200 29606 220000
rect 30286 219200 30342 220000
rect 30930 219200 30986 220000
rect 31666 219200 31722 220000
rect 32402 219200 32458 220000
rect 33138 219200 33194 220000
rect 33782 219200 33838 220000
rect 34518 219200 34574 220000
rect 35254 219200 35310 220000
rect 35990 219200 36046 220000
rect 36726 219200 36782 220000
rect 37370 219200 37426 220000
rect 38106 219200 38162 220000
rect 38842 219200 38898 220000
rect 39578 219200 39634 220000
rect 40222 219200 40278 220000
rect 40958 219200 41014 220000
rect 41694 219200 41750 220000
rect 42430 219200 42486 220000
rect 43074 219200 43130 220000
rect 43810 219200 43866 220000
rect 44546 219200 44602 220000
rect 45282 219200 45338 220000
rect 45926 219200 45982 220000
rect 46662 219200 46718 220000
rect 47398 219200 47454 220000
rect 48134 219200 48190 220000
rect 48870 219200 48926 220000
rect 49514 219200 49570 220000
rect 50250 219200 50306 220000
rect 50986 219200 51042 220000
rect 51722 219200 51778 220000
rect 52366 219200 52422 220000
rect 53102 219200 53158 220000
rect 53838 219200 53894 220000
rect 54574 219200 54630 220000
rect 55218 219200 55274 220000
rect 55954 219200 56010 220000
rect 56690 219200 56746 220000
rect 57426 219200 57482 220000
rect 58070 219200 58126 220000
rect 58806 219200 58862 220000
rect 59542 219200 59598 220000
rect 60278 219200 60334 220000
rect 61014 219200 61070 220000
rect 61658 219200 61714 220000
rect 62394 219200 62450 220000
rect 63130 219200 63186 220000
rect 63866 219200 63922 220000
rect 64510 219200 64566 220000
rect 65246 219200 65302 220000
rect 65982 219200 66038 220000
rect 66718 219200 66774 220000
rect 67362 219200 67418 220000
rect 68098 219200 68154 220000
rect 68834 219200 68890 220000
rect 69570 219200 69626 220000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3146 0 3202 800
rect 3790 0 3846 800
rect 4342 0 4398 800
rect 4894 0 4950 800
rect 5538 0 5594 800
rect 6090 0 6146 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9586 0 9642 800
rect 10138 0 10194 800
rect 10782 0 10838 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15382 0 15438 800
rect 16026 0 16082 800
rect 16578 0 16634 800
rect 17130 0 17186 800
rect 17774 0 17830 800
rect 18326 0 18382 800
rect 18878 0 18934 800
rect 19522 0 19578 800
rect 20074 0 20130 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21822 0 21878 800
rect 22374 0 22430 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24214 0 24270 800
rect 24766 0 24822 800
rect 25318 0 25374 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28262 0 28318 800
rect 28814 0 28870 800
rect 29458 0 29514 800
rect 30010 0 30066 800
rect 30562 0 30618 800
rect 31206 0 31262 800
rect 31758 0 31814 800
rect 32310 0 32366 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34058 0 34114 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36450 0 36506 800
rect 37002 0 37058 800
rect 37554 0 37610 800
rect 38198 0 38254 800
rect 38750 0 38806 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40498 0 40554 800
rect 41050 0 41106 800
rect 41694 0 41750 800
rect 42246 0 42302 800
rect 42798 0 42854 800
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 45190 0 45246 800
rect 45742 0 45798 800
rect 46294 0 46350 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 48134 0 48190 800
rect 48686 0 48742 800
rect 49238 0 49294 800
rect 49882 0 49938 800
rect 50434 0 50490 800
rect 50986 0 51042 800
rect 51630 0 51686 800
rect 52182 0 52238 800
rect 52734 0 52790 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54482 0 54538 800
rect 55126 0 55182 800
rect 55678 0 55734 800
rect 56230 0 56286 800
rect 56874 0 56930 800
rect 57426 0 57482 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59174 0 59230 800
rect 59726 0 59782 800
rect 60370 0 60426 800
rect 60922 0 60978 800
rect 61474 0 61530 800
rect 62118 0 62174 800
rect 62670 0 62726 800
rect 63222 0 63278 800
rect 63866 0 63922 800
rect 64418 0 64474 800
rect 64970 0 65026 800
rect 65614 0 65670 800
rect 66166 0 66222 800
rect 66718 0 66774 800
rect 67362 0 67418 800
rect 67914 0 67970 800
rect 68466 0 68522 800
rect 69110 0 69166 800
rect 69662 0 69718 800
<< obsm2 >>
rect 406 219144 882 219745
rect 1050 219144 1618 219745
rect 1786 219144 2354 219745
rect 2522 219144 3090 219745
rect 3258 219144 3734 219745
rect 3902 219144 4470 219745
rect 4638 219144 5206 219745
rect 5374 219144 5942 219745
rect 6110 219144 6586 219745
rect 6754 219144 7322 219745
rect 7490 219144 8058 219745
rect 8226 219144 8794 219745
rect 8962 219144 9438 219745
rect 9606 219144 10174 219745
rect 10342 219144 10910 219745
rect 11078 219144 11646 219745
rect 11814 219144 12382 219745
rect 12550 219144 13026 219745
rect 13194 219144 13762 219745
rect 13930 219144 14498 219745
rect 14666 219144 15234 219745
rect 15402 219144 15878 219745
rect 16046 219144 16614 219745
rect 16782 219144 17350 219745
rect 17518 219144 18086 219745
rect 18254 219144 18730 219745
rect 18898 219144 19466 219745
rect 19634 219144 20202 219745
rect 20370 219144 20938 219745
rect 21106 219144 21582 219745
rect 21750 219144 22318 219745
rect 22486 219144 23054 219745
rect 23222 219144 23790 219745
rect 23958 219144 24526 219745
rect 24694 219144 25170 219745
rect 25338 219144 25906 219745
rect 26074 219144 26642 219745
rect 26810 219144 27378 219745
rect 27546 219144 28022 219745
rect 28190 219144 28758 219745
rect 28926 219144 29494 219745
rect 29662 219144 30230 219745
rect 30398 219144 30874 219745
rect 31042 219144 31610 219745
rect 31778 219144 32346 219745
rect 32514 219144 33082 219745
rect 33250 219144 33726 219745
rect 33894 219144 34462 219745
rect 34630 219144 35198 219745
rect 35366 219144 35934 219745
rect 36102 219144 36670 219745
rect 36838 219144 37314 219745
rect 37482 219144 38050 219745
rect 38218 219144 38786 219745
rect 38954 219144 39522 219745
rect 39690 219144 40166 219745
rect 40334 219144 40902 219745
rect 41070 219144 41638 219745
rect 41806 219144 42374 219745
rect 42542 219144 43018 219745
rect 43186 219144 43754 219745
rect 43922 219144 44490 219745
rect 44658 219144 45226 219745
rect 45394 219144 45870 219745
rect 46038 219144 46606 219745
rect 46774 219144 47342 219745
rect 47510 219144 48078 219745
rect 48246 219144 48814 219745
rect 48982 219144 49458 219745
rect 49626 219144 50194 219745
rect 50362 219144 50930 219745
rect 51098 219144 51666 219745
rect 51834 219144 52310 219745
rect 52478 219144 53046 219745
rect 53214 219144 53782 219745
rect 53950 219144 54518 219745
rect 54686 219144 55162 219745
rect 55330 219144 55898 219745
rect 56066 219144 56634 219745
rect 56802 219144 57370 219745
rect 57538 219144 58014 219745
rect 58182 219144 58750 219745
rect 58918 219144 59486 219745
rect 59654 219144 60222 219745
rect 60390 219144 60958 219745
rect 61126 219144 61602 219745
rect 61770 219144 62338 219745
rect 62506 219144 63074 219745
rect 63242 219144 63810 219745
rect 63978 219144 64454 219745
rect 64622 219144 65190 219745
rect 65358 219144 65926 219745
rect 66094 219144 66662 219745
rect 66830 219144 67306 219745
rect 67474 219144 68042 219745
rect 68210 219144 68778 219745
rect 68946 219144 69514 219745
rect 69682 219144 69716 219745
rect 294 856 69716 219144
rect 406 303 790 856
rect 958 303 1342 856
rect 1510 303 1986 856
rect 2154 303 2538 856
rect 2706 303 3090 856
rect 3258 303 3734 856
rect 3902 303 4286 856
rect 4454 303 4838 856
rect 5006 303 5482 856
rect 5650 303 6034 856
rect 6202 303 6586 856
rect 6754 303 7230 856
rect 7398 303 7782 856
rect 7950 303 8334 856
rect 8502 303 8978 856
rect 9146 303 9530 856
rect 9698 303 10082 856
rect 10250 303 10726 856
rect 10894 303 11278 856
rect 11446 303 11830 856
rect 11998 303 12474 856
rect 12642 303 13026 856
rect 13194 303 13578 856
rect 13746 303 14222 856
rect 14390 303 14774 856
rect 14942 303 15326 856
rect 15494 303 15970 856
rect 16138 303 16522 856
rect 16690 303 17074 856
rect 17242 303 17718 856
rect 17886 303 18270 856
rect 18438 303 18822 856
rect 18990 303 19466 856
rect 19634 303 20018 856
rect 20186 303 20570 856
rect 20738 303 21214 856
rect 21382 303 21766 856
rect 21934 303 22318 856
rect 22486 303 22962 856
rect 23130 303 23514 856
rect 23682 303 24158 856
rect 24326 303 24710 856
rect 24878 303 25262 856
rect 25430 303 25906 856
rect 26074 303 26458 856
rect 26626 303 27010 856
rect 27178 303 27654 856
rect 27822 303 28206 856
rect 28374 303 28758 856
rect 28926 303 29402 856
rect 29570 303 29954 856
rect 30122 303 30506 856
rect 30674 303 31150 856
rect 31318 303 31702 856
rect 31870 303 32254 856
rect 32422 303 32898 856
rect 33066 303 33450 856
rect 33618 303 34002 856
rect 34170 303 34646 856
rect 34814 303 35198 856
rect 35366 303 35750 856
rect 35918 303 36394 856
rect 36562 303 36946 856
rect 37114 303 37498 856
rect 37666 303 38142 856
rect 38310 303 38694 856
rect 38862 303 39246 856
rect 39414 303 39890 856
rect 40058 303 40442 856
rect 40610 303 40994 856
rect 41162 303 41638 856
rect 41806 303 42190 856
rect 42358 303 42742 856
rect 42910 303 43386 856
rect 43554 303 43938 856
rect 44106 303 44490 856
rect 44658 303 45134 856
rect 45302 303 45686 856
rect 45854 303 46238 856
rect 46406 303 46882 856
rect 47050 303 47434 856
rect 47602 303 48078 856
rect 48246 303 48630 856
rect 48798 303 49182 856
rect 49350 303 49826 856
rect 49994 303 50378 856
rect 50546 303 50930 856
rect 51098 303 51574 856
rect 51742 303 52126 856
rect 52294 303 52678 856
rect 52846 303 53322 856
rect 53490 303 53874 856
rect 54042 303 54426 856
rect 54594 303 55070 856
rect 55238 303 55622 856
rect 55790 303 56174 856
rect 56342 303 56818 856
rect 56986 303 57370 856
rect 57538 303 57922 856
rect 58090 303 58566 856
rect 58734 303 59118 856
rect 59286 303 59670 856
rect 59838 303 60314 856
rect 60482 303 60866 856
rect 61034 303 61418 856
rect 61586 303 62062 856
rect 62230 303 62614 856
rect 62782 303 63166 856
rect 63334 303 63810 856
rect 63978 303 64362 856
rect 64530 303 64914 856
rect 65082 303 65558 856
rect 65726 303 66110 856
rect 66278 303 66662 856
rect 66830 303 67306 856
rect 67474 303 67858 856
rect 68026 303 68410 856
rect 68578 303 69054 856
rect 69222 303 69606 856
<< metal3 >>
rect 0 219648 800 219768
rect 69200 219376 70000 219496
rect 0 219104 800 219224
rect 0 218560 800 218680
rect 69200 218288 70000 218408
rect 0 218016 800 218136
rect 0 217472 800 217592
rect 69200 217200 70000 217320
rect 0 216928 800 217048
rect 0 216384 800 216504
rect 0 215840 800 215960
rect 69200 215976 70000 216096
rect 0 215296 800 215416
rect 0 214752 800 214872
rect 69200 214888 70000 215008
rect 0 214208 800 214328
rect 0 213664 800 213784
rect 69200 213800 70000 213920
rect 0 213120 800 213240
rect 0 212576 800 212696
rect 69200 212712 70000 212832
rect 0 212032 800 212152
rect 0 211488 800 211608
rect 69200 211488 70000 211608
rect 0 210944 800 211064
rect 0 210400 800 210520
rect 69200 210400 70000 210520
rect 0 209856 800 209976
rect 0 209312 800 209432
rect 69200 209312 70000 209432
rect 0 208768 800 208888
rect 0 208224 800 208344
rect 69200 208224 70000 208344
rect 0 207544 800 207664
rect 0 207000 800 207120
rect 69200 207000 70000 207120
rect 0 206456 800 206576
rect 0 205912 800 206032
rect 69200 205912 70000 206032
rect 0 205368 800 205488
rect 0 204824 800 204944
rect 69200 204824 70000 204944
rect 0 204280 800 204400
rect 0 203736 800 203856
rect 69200 203736 70000 203856
rect 0 203192 800 203312
rect 0 202648 800 202768
rect 69200 202512 70000 202632
rect 0 202104 800 202224
rect 0 201560 800 201680
rect 69200 201424 70000 201544
rect 0 201016 800 201136
rect 0 200472 800 200592
rect 69200 200336 70000 200456
rect 0 199928 800 200048
rect 0 199384 800 199504
rect 69200 199248 70000 199368
rect 0 198840 800 198960
rect 0 198296 800 198416
rect 69200 198024 70000 198144
rect 0 197752 800 197872
rect 0 197208 800 197328
rect 69200 196936 70000 197056
rect 0 196664 800 196784
rect 0 196120 800 196240
rect 69200 195848 70000 195968
rect 0 195440 800 195560
rect 0 194896 800 195016
rect 69200 194760 70000 194880
rect 0 194352 800 194472
rect 0 193808 800 193928
rect 69200 193536 70000 193656
rect 0 193264 800 193384
rect 0 192720 800 192840
rect 69200 192448 70000 192568
rect 0 192176 800 192296
rect 0 191632 800 191752
rect 69200 191360 70000 191480
rect 0 191088 800 191208
rect 0 190544 800 190664
rect 69200 190272 70000 190392
rect 0 190000 800 190120
rect 0 189456 800 189576
rect 0 188912 800 189032
rect 69200 189048 70000 189168
rect 0 188368 800 188488
rect 0 187824 800 187944
rect 69200 187960 70000 188080
rect 0 187280 800 187400
rect 0 186736 800 186856
rect 69200 186872 70000 186992
rect 0 186192 800 186312
rect 0 185648 800 185768
rect 69200 185784 70000 185904
rect 0 185104 800 185224
rect 0 184560 800 184680
rect 69200 184560 70000 184680
rect 0 184016 800 184136
rect 0 183336 800 183456
rect 69200 183472 70000 183592
rect 0 182792 800 182912
rect 0 182248 800 182368
rect 69200 182384 70000 182504
rect 0 181704 800 181824
rect 0 181160 800 181280
rect 69200 181296 70000 181416
rect 0 180616 800 180736
rect 0 180072 800 180192
rect 69200 180072 70000 180192
rect 0 179528 800 179648
rect 0 178984 800 179104
rect 69200 178984 70000 179104
rect 0 178440 800 178560
rect 0 177896 800 178016
rect 69200 177896 70000 178016
rect 0 177352 800 177472
rect 0 176808 800 176928
rect 69200 176808 70000 176928
rect 0 176264 800 176384
rect 0 175720 800 175840
rect 69200 175584 70000 175704
rect 0 175176 800 175296
rect 0 174632 800 174752
rect 69200 174496 70000 174616
rect 0 174088 800 174208
rect 0 173544 800 173664
rect 69200 173408 70000 173528
rect 0 173000 800 173120
rect 0 172456 800 172576
rect 69200 172320 70000 172440
rect 0 171912 800 172032
rect 0 171232 800 171352
rect 69200 171096 70000 171216
rect 0 170688 800 170808
rect 0 170144 800 170264
rect 69200 170008 70000 170128
rect 0 169600 800 169720
rect 0 169056 800 169176
rect 69200 168920 70000 169040
rect 0 168512 800 168632
rect 0 167968 800 168088
rect 69200 167832 70000 167952
rect 0 167424 800 167544
rect 0 166880 800 167000
rect 69200 166608 70000 166728
rect 0 166336 800 166456
rect 0 165792 800 165912
rect 69200 165520 70000 165640
rect 0 165248 800 165368
rect 0 164704 800 164824
rect 69200 164432 70000 164552
rect 0 164160 800 164280
rect 0 163616 800 163736
rect 0 163072 800 163192
rect 69200 163208 70000 163328
rect 0 162528 800 162648
rect 0 161984 800 162104
rect 69200 162120 70000 162240
rect 0 161440 800 161560
rect 0 160896 800 161016
rect 69200 161032 70000 161152
rect 0 160352 800 160472
rect 0 159808 800 159928
rect 69200 159944 70000 160064
rect 0 159264 800 159384
rect 0 158584 800 158704
rect 69200 158720 70000 158840
rect 0 158040 800 158160
rect 0 157496 800 157616
rect 69200 157632 70000 157752
rect 0 156952 800 157072
rect 0 156408 800 156528
rect 69200 156544 70000 156664
rect 0 155864 800 155984
rect 0 155320 800 155440
rect 69200 155456 70000 155576
rect 0 154776 800 154896
rect 0 154232 800 154352
rect 69200 154232 70000 154352
rect 0 153688 800 153808
rect 0 153144 800 153264
rect 69200 153144 70000 153264
rect 0 152600 800 152720
rect 0 152056 800 152176
rect 69200 152056 70000 152176
rect 0 151512 800 151632
rect 0 150968 800 151088
rect 69200 150968 70000 151088
rect 0 150424 800 150544
rect 0 149880 800 150000
rect 69200 149744 70000 149864
rect 0 149336 800 149456
rect 0 148792 800 148912
rect 69200 148656 70000 148776
rect 0 148248 800 148368
rect 0 147704 800 147824
rect 69200 147568 70000 147688
rect 0 147160 800 147280
rect 0 146480 800 146600
rect 69200 146480 70000 146600
rect 0 145936 800 146056
rect 0 145392 800 145512
rect 69200 145256 70000 145376
rect 0 144848 800 144968
rect 0 144304 800 144424
rect 69200 144168 70000 144288
rect 0 143760 800 143880
rect 0 143216 800 143336
rect 69200 143080 70000 143200
rect 0 142672 800 142792
rect 0 142128 800 142248
rect 69200 141992 70000 142112
rect 0 141584 800 141704
rect 0 141040 800 141160
rect 69200 140768 70000 140888
rect 0 140496 800 140616
rect 0 139952 800 140072
rect 69200 139680 70000 139800
rect 0 139408 800 139528
rect 0 138864 800 138984
rect 69200 138592 70000 138712
rect 0 138320 800 138440
rect 0 137776 800 137896
rect 69200 137504 70000 137624
rect 0 137232 800 137352
rect 0 136688 800 136808
rect 0 136144 800 136264
rect 69200 136280 70000 136400
rect 0 135600 800 135720
rect 0 135056 800 135176
rect 69200 135192 70000 135312
rect 0 134376 800 134496
rect 69200 134104 70000 134224
rect 0 133832 800 133952
rect 0 133288 800 133408
rect 69200 133016 70000 133136
rect 0 132744 800 132864
rect 0 132200 800 132320
rect 0 131656 800 131776
rect 69200 131792 70000 131912
rect 0 131112 800 131232
rect 0 130568 800 130688
rect 69200 130704 70000 130824
rect 0 130024 800 130144
rect 0 129480 800 129600
rect 69200 129616 70000 129736
rect 0 128936 800 129056
rect 0 128392 800 128512
rect 69200 128528 70000 128648
rect 0 127848 800 127968
rect 0 127304 800 127424
rect 69200 127304 70000 127424
rect 0 126760 800 126880
rect 0 126216 800 126336
rect 69200 126216 70000 126336
rect 0 125672 800 125792
rect 0 125128 800 125248
rect 69200 125128 70000 125248
rect 0 124584 800 124704
rect 0 124040 800 124160
rect 69200 124040 70000 124160
rect 0 123496 800 123616
rect 0 122952 800 123072
rect 69200 122816 70000 122936
rect 0 122272 800 122392
rect 0 121728 800 121848
rect 69200 121728 70000 121848
rect 0 121184 800 121304
rect 0 120640 800 120760
rect 69200 120640 70000 120760
rect 0 120096 800 120216
rect 0 119552 800 119672
rect 69200 119552 70000 119672
rect 0 119008 800 119128
rect 0 118464 800 118584
rect 69200 118328 70000 118448
rect 0 117920 800 118040
rect 0 117376 800 117496
rect 69200 117240 70000 117360
rect 0 116832 800 116952
rect 0 116288 800 116408
rect 69200 116152 70000 116272
rect 0 115744 800 115864
rect 0 115200 800 115320
rect 69200 115064 70000 115184
rect 0 114656 800 114776
rect 0 114112 800 114232
rect 69200 113840 70000 113960
rect 0 113568 800 113688
rect 0 113024 800 113144
rect 69200 112752 70000 112872
rect 0 112480 800 112600
rect 0 111936 800 112056
rect 69200 111664 70000 111784
rect 0 111392 800 111512
rect 0 110848 800 110968
rect 69200 110576 70000 110696
rect 0 110304 800 110424
rect 0 109624 800 109744
rect 69200 109352 70000 109472
rect 0 109080 800 109200
rect 0 108536 800 108656
rect 69200 108264 70000 108384
rect 0 107992 800 108112
rect 0 107448 800 107568
rect 69200 107176 70000 107296
rect 0 106904 800 107024
rect 0 106360 800 106480
rect 0 105816 800 105936
rect 69200 105952 70000 106072
rect 0 105272 800 105392
rect 0 104728 800 104848
rect 69200 104864 70000 104984
rect 0 104184 800 104304
rect 0 103640 800 103760
rect 69200 103776 70000 103896
rect 0 103096 800 103216
rect 0 102552 800 102672
rect 69200 102688 70000 102808
rect 0 102008 800 102128
rect 0 101464 800 101584
rect 69200 101464 70000 101584
rect 0 100920 800 101040
rect 0 100376 800 100496
rect 69200 100376 70000 100496
rect 0 99832 800 99952
rect 0 99288 800 99408
rect 69200 99288 70000 99408
rect 0 98744 800 98864
rect 0 98200 800 98320
rect 69200 98200 70000 98320
rect 0 97520 800 97640
rect 0 96976 800 97096
rect 69200 96976 70000 97096
rect 0 96432 800 96552
rect 0 95888 800 96008
rect 69200 95888 70000 96008
rect 0 95344 800 95464
rect 0 94800 800 94920
rect 69200 94800 70000 94920
rect 0 94256 800 94376
rect 0 93712 800 93832
rect 69200 93712 70000 93832
rect 0 93168 800 93288
rect 0 92624 800 92744
rect 69200 92488 70000 92608
rect 0 92080 800 92200
rect 0 91536 800 91656
rect 69200 91400 70000 91520
rect 0 90992 800 91112
rect 0 90448 800 90568
rect 69200 90312 70000 90432
rect 0 89904 800 90024
rect 0 89360 800 89480
rect 69200 89224 70000 89344
rect 0 88816 800 88936
rect 0 88272 800 88392
rect 69200 88000 70000 88120
rect 0 87728 800 87848
rect 0 87184 800 87304
rect 69200 86912 70000 87032
rect 0 86640 800 86760
rect 0 86096 800 86216
rect 69200 85824 70000 85944
rect 0 85416 800 85536
rect 0 84872 800 84992
rect 69200 84736 70000 84856
rect 0 84328 800 84448
rect 0 83784 800 83904
rect 69200 83512 70000 83632
rect 0 83240 800 83360
rect 0 82696 800 82816
rect 69200 82424 70000 82544
rect 0 82152 800 82272
rect 0 81608 800 81728
rect 69200 81336 70000 81456
rect 0 81064 800 81184
rect 0 80520 800 80640
rect 69200 80248 70000 80368
rect 0 79976 800 80096
rect 0 79432 800 79552
rect 0 78888 800 79008
rect 69200 79024 70000 79144
rect 0 78344 800 78464
rect 0 77800 800 77920
rect 69200 77936 70000 78056
rect 0 77256 800 77376
rect 0 76712 800 76832
rect 69200 76848 70000 76968
rect 0 76168 800 76288
rect 0 75624 800 75744
rect 69200 75760 70000 75880
rect 0 75080 800 75200
rect 0 74536 800 74656
rect 69200 74536 70000 74656
rect 0 73992 800 74112
rect 0 73312 800 73432
rect 69200 73448 70000 73568
rect 0 72768 800 72888
rect 0 72224 800 72344
rect 69200 72360 70000 72480
rect 0 71680 800 71800
rect 0 71136 800 71256
rect 69200 71272 70000 71392
rect 0 70592 800 70712
rect 0 70048 800 70168
rect 69200 70048 70000 70168
rect 0 69504 800 69624
rect 0 68960 800 69080
rect 69200 68960 70000 69080
rect 0 68416 800 68536
rect 0 67872 800 67992
rect 69200 67872 70000 67992
rect 0 67328 800 67448
rect 0 66784 800 66904
rect 69200 66784 70000 66904
rect 0 66240 800 66360
rect 0 65696 800 65816
rect 69200 65560 70000 65680
rect 0 65152 800 65272
rect 0 64608 800 64728
rect 69200 64472 70000 64592
rect 0 64064 800 64184
rect 0 63520 800 63640
rect 69200 63384 70000 63504
rect 0 62976 800 63096
rect 0 62432 800 62552
rect 69200 62296 70000 62416
rect 0 61888 800 62008
rect 0 61208 800 61328
rect 69200 61072 70000 61192
rect 0 60664 800 60784
rect 0 60120 800 60240
rect 69200 59984 70000 60104
rect 0 59576 800 59696
rect 0 59032 800 59152
rect 69200 58896 70000 59016
rect 0 58488 800 58608
rect 0 57944 800 58064
rect 69200 57808 70000 57928
rect 0 57400 800 57520
rect 0 56856 800 56976
rect 69200 56584 70000 56704
rect 0 56312 800 56432
rect 0 55768 800 55888
rect 69200 55496 70000 55616
rect 0 55224 800 55344
rect 0 54680 800 54800
rect 69200 54408 70000 54528
rect 0 54136 800 54256
rect 0 53592 800 53712
rect 0 53048 800 53168
rect 69200 53184 70000 53304
rect 0 52504 800 52624
rect 0 51960 800 52080
rect 69200 52096 70000 52216
rect 0 51416 800 51536
rect 0 50872 800 50992
rect 69200 51008 70000 51128
rect 0 50328 800 50448
rect 0 49784 800 49904
rect 69200 49920 70000 50040
rect 0 49240 800 49360
rect 0 48560 800 48680
rect 69200 48696 70000 48816
rect 0 48016 800 48136
rect 0 47472 800 47592
rect 69200 47608 70000 47728
rect 0 46928 800 47048
rect 0 46384 800 46504
rect 69200 46520 70000 46640
rect 0 45840 800 45960
rect 0 45296 800 45416
rect 69200 45432 70000 45552
rect 0 44752 800 44872
rect 0 44208 800 44328
rect 69200 44208 70000 44328
rect 0 43664 800 43784
rect 0 43120 800 43240
rect 69200 43120 70000 43240
rect 0 42576 800 42696
rect 0 42032 800 42152
rect 69200 42032 70000 42152
rect 0 41488 800 41608
rect 0 40944 800 41064
rect 69200 40944 70000 41064
rect 0 40400 800 40520
rect 0 39856 800 39976
rect 69200 39720 70000 39840
rect 0 39312 800 39432
rect 0 38768 800 38888
rect 69200 38632 70000 38752
rect 0 38224 800 38344
rect 0 37680 800 37800
rect 69200 37544 70000 37664
rect 0 37136 800 37256
rect 0 36456 800 36576
rect 69200 36456 70000 36576
rect 0 35912 800 36032
rect 0 35368 800 35488
rect 69200 35232 70000 35352
rect 0 34824 800 34944
rect 0 34280 800 34400
rect 69200 34144 70000 34264
rect 0 33736 800 33856
rect 0 33192 800 33312
rect 69200 33056 70000 33176
rect 0 32648 800 32768
rect 0 32104 800 32224
rect 69200 31968 70000 32088
rect 0 31560 800 31680
rect 0 31016 800 31136
rect 69200 30744 70000 30864
rect 0 30472 800 30592
rect 0 29928 800 30048
rect 69200 29656 70000 29776
rect 0 29384 800 29504
rect 0 28840 800 28960
rect 69200 28568 70000 28688
rect 0 28296 800 28416
rect 0 27752 800 27872
rect 69200 27480 70000 27600
rect 0 27208 800 27328
rect 0 26664 800 26784
rect 0 26120 800 26240
rect 69200 26256 70000 26376
rect 0 25576 800 25696
rect 0 25032 800 25152
rect 69200 25168 70000 25288
rect 0 24352 800 24472
rect 69200 24080 70000 24200
rect 0 23808 800 23928
rect 0 23264 800 23384
rect 69200 22992 70000 23112
rect 0 22720 800 22840
rect 0 22176 800 22296
rect 0 21632 800 21752
rect 69200 21768 70000 21888
rect 0 21088 800 21208
rect 0 20544 800 20664
rect 69200 20680 70000 20800
rect 0 20000 800 20120
rect 0 19456 800 19576
rect 69200 19592 70000 19712
rect 0 18912 800 19032
rect 0 18368 800 18488
rect 69200 18504 70000 18624
rect 0 17824 800 17944
rect 0 17280 800 17400
rect 69200 17280 70000 17400
rect 0 16736 800 16856
rect 0 16192 800 16312
rect 69200 16192 70000 16312
rect 0 15648 800 15768
rect 0 15104 800 15224
rect 69200 15104 70000 15224
rect 0 14560 800 14680
rect 0 14016 800 14136
rect 69200 14016 70000 14136
rect 0 13472 800 13592
rect 0 12928 800 13048
rect 69200 12792 70000 12912
rect 0 12248 800 12368
rect 0 11704 800 11824
rect 69200 11704 70000 11824
rect 0 11160 800 11280
rect 0 10616 800 10736
rect 69200 10616 70000 10736
rect 0 10072 800 10192
rect 0 9528 800 9648
rect 69200 9528 70000 9648
rect 0 8984 800 9104
rect 0 8440 800 8560
rect 69200 8304 70000 8424
rect 0 7896 800 8016
rect 0 7352 800 7472
rect 69200 7216 70000 7336
rect 0 6808 800 6928
rect 0 6264 800 6384
rect 69200 6128 70000 6248
rect 0 5720 800 5840
rect 0 5176 800 5296
rect 69200 5040 70000 5160
rect 0 4632 800 4752
rect 0 4088 800 4208
rect 69200 3816 70000 3936
rect 0 3544 800 3664
rect 0 3000 800 3120
rect 69200 2728 70000 2848
rect 0 2456 800 2576
rect 0 1912 800 2032
rect 69200 1640 70000 1760
rect 0 1368 800 1488
rect 0 824 800 944
rect 69200 552 70000 672
rect 0 280 800 400
<< obsm3 >>
rect 880 219576 69200 219741
rect 880 219568 69120 219576
rect 289 219304 69120 219568
rect 880 219296 69120 219304
rect 880 219024 69200 219296
rect 289 218760 69200 219024
rect 880 218488 69200 218760
rect 880 218480 69120 218488
rect 289 218216 69120 218480
rect 880 218208 69120 218216
rect 880 217936 69200 218208
rect 289 217672 69200 217936
rect 880 217400 69200 217672
rect 880 217392 69120 217400
rect 289 217128 69120 217392
rect 880 217120 69120 217128
rect 880 216848 69200 217120
rect 289 216584 69200 216848
rect 880 216304 69200 216584
rect 289 216176 69200 216304
rect 289 216040 69120 216176
rect 880 215896 69120 216040
rect 880 215760 69200 215896
rect 289 215496 69200 215760
rect 880 215216 69200 215496
rect 289 215088 69200 215216
rect 289 214952 69120 215088
rect 880 214808 69120 214952
rect 880 214672 69200 214808
rect 289 214408 69200 214672
rect 880 214128 69200 214408
rect 289 214000 69200 214128
rect 289 213864 69120 214000
rect 880 213720 69120 213864
rect 880 213584 69200 213720
rect 289 213320 69200 213584
rect 880 213040 69200 213320
rect 289 212912 69200 213040
rect 289 212776 69120 212912
rect 880 212632 69120 212776
rect 880 212496 69200 212632
rect 289 212232 69200 212496
rect 880 211952 69200 212232
rect 289 211688 69200 211952
rect 880 211408 69120 211688
rect 289 211144 69200 211408
rect 880 210864 69200 211144
rect 289 210600 69200 210864
rect 880 210320 69120 210600
rect 289 210056 69200 210320
rect 880 209776 69200 210056
rect 289 209512 69200 209776
rect 880 209232 69120 209512
rect 289 208968 69200 209232
rect 880 208688 69200 208968
rect 289 208424 69200 208688
rect 880 208144 69120 208424
rect 289 207744 69200 208144
rect 880 207464 69200 207744
rect 289 207200 69200 207464
rect 880 206920 69120 207200
rect 289 206656 69200 206920
rect 880 206376 69200 206656
rect 289 206112 69200 206376
rect 880 205832 69120 206112
rect 289 205568 69200 205832
rect 880 205288 69200 205568
rect 289 205024 69200 205288
rect 880 204744 69120 205024
rect 289 204480 69200 204744
rect 880 204200 69200 204480
rect 289 203936 69200 204200
rect 880 203656 69120 203936
rect 289 203392 69200 203656
rect 880 203112 69200 203392
rect 289 202848 69200 203112
rect 880 202712 69200 202848
rect 880 202568 69120 202712
rect 289 202432 69120 202568
rect 289 202304 69200 202432
rect 880 202024 69200 202304
rect 289 201760 69200 202024
rect 880 201624 69200 201760
rect 880 201480 69120 201624
rect 289 201344 69120 201480
rect 289 201216 69200 201344
rect 880 200936 69200 201216
rect 289 200672 69200 200936
rect 880 200536 69200 200672
rect 880 200392 69120 200536
rect 289 200256 69120 200392
rect 289 200128 69200 200256
rect 880 199848 69200 200128
rect 289 199584 69200 199848
rect 880 199448 69200 199584
rect 880 199304 69120 199448
rect 289 199168 69120 199304
rect 289 199040 69200 199168
rect 880 198760 69200 199040
rect 289 198496 69200 198760
rect 880 198224 69200 198496
rect 880 198216 69120 198224
rect 289 197952 69120 198216
rect 880 197944 69120 197952
rect 880 197672 69200 197944
rect 289 197408 69200 197672
rect 880 197136 69200 197408
rect 880 197128 69120 197136
rect 289 196864 69120 197128
rect 880 196856 69120 196864
rect 880 196584 69200 196856
rect 289 196320 69200 196584
rect 880 196048 69200 196320
rect 880 196040 69120 196048
rect 289 195768 69120 196040
rect 289 195640 69200 195768
rect 880 195360 69200 195640
rect 289 195096 69200 195360
rect 880 194960 69200 195096
rect 880 194816 69120 194960
rect 289 194680 69120 194816
rect 289 194552 69200 194680
rect 880 194272 69200 194552
rect 289 194008 69200 194272
rect 880 193736 69200 194008
rect 880 193728 69120 193736
rect 289 193464 69120 193728
rect 880 193456 69120 193464
rect 880 193184 69200 193456
rect 289 192920 69200 193184
rect 880 192648 69200 192920
rect 880 192640 69120 192648
rect 289 192376 69120 192640
rect 880 192368 69120 192376
rect 880 192096 69200 192368
rect 289 191832 69200 192096
rect 880 191560 69200 191832
rect 880 191552 69120 191560
rect 289 191288 69120 191552
rect 880 191280 69120 191288
rect 880 191008 69200 191280
rect 289 190744 69200 191008
rect 880 190472 69200 190744
rect 880 190464 69120 190472
rect 289 190200 69120 190464
rect 880 190192 69120 190200
rect 880 189920 69200 190192
rect 289 189656 69200 189920
rect 880 189376 69200 189656
rect 289 189248 69200 189376
rect 289 189112 69120 189248
rect 880 188968 69120 189112
rect 880 188832 69200 188968
rect 289 188568 69200 188832
rect 880 188288 69200 188568
rect 289 188160 69200 188288
rect 289 188024 69120 188160
rect 880 187880 69120 188024
rect 880 187744 69200 187880
rect 289 187480 69200 187744
rect 880 187200 69200 187480
rect 289 187072 69200 187200
rect 289 186936 69120 187072
rect 880 186792 69120 186936
rect 880 186656 69200 186792
rect 289 186392 69200 186656
rect 880 186112 69200 186392
rect 289 185984 69200 186112
rect 289 185848 69120 185984
rect 880 185704 69120 185848
rect 880 185568 69200 185704
rect 289 185304 69200 185568
rect 880 185024 69200 185304
rect 289 184760 69200 185024
rect 880 184480 69120 184760
rect 289 184216 69200 184480
rect 880 183936 69200 184216
rect 289 183672 69200 183936
rect 289 183536 69120 183672
rect 880 183392 69120 183536
rect 880 183256 69200 183392
rect 289 182992 69200 183256
rect 880 182712 69200 182992
rect 289 182584 69200 182712
rect 289 182448 69120 182584
rect 880 182304 69120 182448
rect 880 182168 69200 182304
rect 289 181904 69200 182168
rect 880 181624 69200 181904
rect 289 181496 69200 181624
rect 289 181360 69120 181496
rect 880 181216 69120 181360
rect 880 181080 69200 181216
rect 289 180816 69200 181080
rect 880 180536 69200 180816
rect 289 180272 69200 180536
rect 880 179992 69120 180272
rect 289 179728 69200 179992
rect 880 179448 69200 179728
rect 289 179184 69200 179448
rect 880 178904 69120 179184
rect 289 178640 69200 178904
rect 880 178360 69200 178640
rect 289 178096 69200 178360
rect 880 177816 69120 178096
rect 289 177552 69200 177816
rect 880 177272 69200 177552
rect 289 177008 69200 177272
rect 880 176728 69120 177008
rect 289 176464 69200 176728
rect 880 176184 69200 176464
rect 289 175920 69200 176184
rect 880 175784 69200 175920
rect 880 175640 69120 175784
rect 289 175504 69120 175640
rect 289 175376 69200 175504
rect 880 175096 69200 175376
rect 289 174832 69200 175096
rect 880 174696 69200 174832
rect 880 174552 69120 174696
rect 289 174416 69120 174552
rect 289 174288 69200 174416
rect 880 174008 69200 174288
rect 289 173744 69200 174008
rect 880 173608 69200 173744
rect 880 173464 69120 173608
rect 289 173328 69120 173464
rect 289 173200 69200 173328
rect 880 172920 69200 173200
rect 289 172656 69200 172920
rect 880 172520 69200 172656
rect 880 172376 69120 172520
rect 289 172240 69120 172376
rect 289 172112 69200 172240
rect 880 171832 69200 172112
rect 289 171432 69200 171832
rect 880 171296 69200 171432
rect 880 171152 69120 171296
rect 289 171016 69120 171152
rect 289 170888 69200 171016
rect 880 170608 69200 170888
rect 289 170344 69200 170608
rect 880 170208 69200 170344
rect 880 170064 69120 170208
rect 289 169928 69120 170064
rect 289 169800 69200 169928
rect 880 169520 69200 169800
rect 289 169256 69200 169520
rect 880 169120 69200 169256
rect 880 168976 69120 169120
rect 289 168840 69120 168976
rect 289 168712 69200 168840
rect 880 168432 69200 168712
rect 289 168168 69200 168432
rect 880 168032 69200 168168
rect 880 167888 69120 168032
rect 289 167752 69120 167888
rect 289 167624 69200 167752
rect 880 167344 69200 167624
rect 289 167080 69200 167344
rect 880 166808 69200 167080
rect 880 166800 69120 166808
rect 289 166536 69120 166800
rect 880 166528 69120 166536
rect 880 166256 69200 166528
rect 289 165992 69200 166256
rect 880 165720 69200 165992
rect 880 165712 69120 165720
rect 289 165448 69120 165712
rect 880 165440 69120 165448
rect 880 165168 69200 165440
rect 289 164904 69200 165168
rect 880 164632 69200 164904
rect 880 164624 69120 164632
rect 289 164360 69120 164624
rect 880 164352 69120 164360
rect 880 164080 69200 164352
rect 289 163816 69200 164080
rect 880 163536 69200 163816
rect 289 163408 69200 163536
rect 289 163272 69120 163408
rect 880 163128 69120 163272
rect 880 162992 69200 163128
rect 289 162728 69200 162992
rect 880 162448 69200 162728
rect 289 162320 69200 162448
rect 289 162184 69120 162320
rect 880 162040 69120 162184
rect 880 161904 69200 162040
rect 289 161640 69200 161904
rect 880 161360 69200 161640
rect 289 161232 69200 161360
rect 289 161096 69120 161232
rect 880 160952 69120 161096
rect 880 160816 69200 160952
rect 289 160552 69200 160816
rect 880 160272 69200 160552
rect 289 160144 69200 160272
rect 289 160008 69120 160144
rect 880 159864 69120 160008
rect 880 159728 69200 159864
rect 289 159464 69200 159728
rect 880 159184 69200 159464
rect 289 158920 69200 159184
rect 289 158784 69120 158920
rect 880 158640 69120 158784
rect 880 158504 69200 158640
rect 289 158240 69200 158504
rect 880 157960 69200 158240
rect 289 157832 69200 157960
rect 289 157696 69120 157832
rect 880 157552 69120 157696
rect 880 157416 69200 157552
rect 289 157152 69200 157416
rect 880 156872 69200 157152
rect 289 156744 69200 156872
rect 289 156608 69120 156744
rect 880 156464 69120 156608
rect 880 156328 69200 156464
rect 289 156064 69200 156328
rect 880 155784 69200 156064
rect 289 155656 69200 155784
rect 289 155520 69120 155656
rect 880 155376 69120 155520
rect 880 155240 69200 155376
rect 289 154976 69200 155240
rect 880 154696 69200 154976
rect 289 154432 69200 154696
rect 880 154152 69120 154432
rect 289 153888 69200 154152
rect 880 153608 69200 153888
rect 289 153344 69200 153608
rect 880 153064 69120 153344
rect 289 152800 69200 153064
rect 880 152520 69200 152800
rect 289 152256 69200 152520
rect 880 151976 69120 152256
rect 289 151712 69200 151976
rect 880 151432 69200 151712
rect 289 151168 69200 151432
rect 880 150888 69120 151168
rect 289 150624 69200 150888
rect 880 150344 69200 150624
rect 289 150080 69200 150344
rect 880 149944 69200 150080
rect 880 149800 69120 149944
rect 289 149664 69120 149800
rect 289 149536 69200 149664
rect 880 149256 69200 149536
rect 289 148992 69200 149256
rect 880 148856 69200 148992
rect 880 148712 69120 148856
rect 289 148576 69120 148712
rect 289 148448 69200 148576
rect 880 148168 69200 148448
rect 289 147904 69200 148168
rect 880 147768 69200 147904
rect 880 147624 69120 147768
rect 289 147488 69120 147624
rect 289 147360 69200 147488
rect 880 147080 69200 147360
rect 289 146680 69200 147080
rect 880 146400 69120 146680
rect 289 146136 69200 146400
rect 880 145856 69200 146136
rect 289 145592 69200 145856
rect 880 145456 69200 145592
rect 880 145312 69120 145456
rect 289 145176 69120 145312
rect 289 145048 69200 145176
rect 880 144768 69200 145048
rect 289 144504 69200 144768
rect 880 144368 69200 144504
rect 880 144224 69120 144368
rect 289 144088 69120 144224
rect 289 143960 69200 144088
rect 880 143680 69200 143960
rect 289 143416 69200 143680
rect 880 143280 69200 143416
rect 880 143136 69120 143280
rect 289 143000 69120 143136
rect 289 142872 69200 143000
rect 880 142592 69200 142872
rect 289 142328 69200 142592
rect 880 142192 69200 142328
rect 880 142048 69120 142192
rect 289 141912 69120 142048
rect 289 141784 69200 141912
rect 880 141504 69200 141784
rect 289 141240 69200 141504
rect 880 140968 69200 141240
rect 880 140960 69120 140968
rect 289 140696 69120 140960
rect 880 140688 69120 140696
rect 880 140416 69200 140688
rect 289 140152 69200 140416
rect 880 139880 69200 140152
rect 880 139872 69120 139880
rect 289 139608 69120 139872
rect 880 139600 69120 139608
rect 880 139328 69200 139600
rect 289 139064 69200 139328
rect 880 138792 69200 139064
rect 880 138784 69120 138792
rect 289 138520 69120 138784
rect 880 138512 69120 138520
rect 880 138240 69200 138512
rect 289 137976 69200 138240
rect 880 137704 69200 137976
rect 880 137696 69120 137704
rect 289 137432 69120 137696
rect 880 137424 69120 137432
rect 880 137152 69200 137424
rect 289 136888 69200 137152
rect 880 136608 69200 136888
rect 289 136480 69200 136608
rect 289 136344 69120 136480
rect 880 136200 69120 136344
rect 880 136064 69200 136200
rect 289 135800 69200 136064
rect 880 135520 69200 135800
rect 289 135392 69200 135520
rect 289 135256 69120 135392
rect 880 135112 69120 135256
rect 880 134976 69200 135112
rect 289 134576 69200 134976
rect 880 134304 69200 134576
rect 880 134296 69120 134304
rect 289 134032 69120 134296
rect 880 134024 69120 134032
rect 880 133752 69200 134024
rect 289 133488 69200 133752
rect 880 133216 69200 133488
rect 880 133208 69120 133216
rect 289 132944 69120 133208
rect 880 132936 69120 132944
rect 880 132664 69200 132936
rect 289 132400 69200 132664
rect 880 132120 69200 132400
rect 289 131992 69200 132120
rect 289 131856 69120 131992
rect 880 131712 69120 131856
rect 880 131576 69200 131712
rect 289 131312 69200 131576
rect 880 131032 69200 131312
rect 289 130904 69200 131032
rect 289 130768 69120 130904
rect 880 130624 69120 130768
rect 880 130488 69200 130624
rect 289 130224 69200 130488
rect 880 129944 69200 130224
rect 289 129816 69200 129944
rect 289 129680 69120 129816
rect 880 129536 69120 129680
rect 880 129400 69200 129536
rect 289 129136 69200 129400
rect 880 128856 69200 129136
rect 289 128728 69200 128856
rect 289 128592 69120 128728
rect 880 128448 69120 128592
rect 880 128312 69200 128448
rect 289 128048 69200 128312
rect 880 127768 69200 128048
rect 289 127504 69200 127768
rect 880 127224 69120 127504
rect 289 126960 69200 127224
rect 880 126680 69200 126960
rect 289 126416 69200 126680
rect 880 126136 69120 126416
rect 289 125872 69200 126136
rect 880 125592 69200 125872
rect 289 125328 69200 125592
rect 880 125048 69120 125328
rect 289 124784 69200 125048
rect 880 124504 69200 124784
rect 289 124240 69200 124504
rect 880 123960 69120 124240
rect 289 123696 69200 123960
rect 880 123416 69200 123696
rect 289 123152 69200 123416
rect 880 123016 69200 123152
rect 880 122872 69120 123016
rect 289 122736 69120 122872
rect 289 122472 69200 122736
rect 880 122192 69200 122472
rect 289 121928 69200 122192
rect 880 121648 69120 121928
rect 289 121384 69200 121648
rect 880 121104 69200 121384
rect 289 120840 69200 121104
rect 880 120560 69120 120840
rect 289 120296 69200 120560
rect 880 120016 69200 120296
rect 289 119752 69200 120016
rect 880 119472 69120 119752
rect 289 119208 69200 119472
rect 880 118928 69200 119208
rect 289 118664 69200 118928
rect 880 118528 69200 118664
rect 880 118384 69120 118528
rect 289 118248 69120 118384
rect 289 118120 69200 118248
rect 880 117840 69200 118120
rect 289 117576 69200 117840
rect 880 117440 69200 117576
rect 880 117296 69120 117440
rect 289 117160 69120 117296
rect 289 117032 69200 117160
rect 880 116752 69200 117032
rect 289 116488 69200 116752
rect 880 116352 69200 116488
rect 880 116208 69120 116352
rect 289 116072 69120 116208
rect 289 115944 69200 116072
rect 880 115664 69200 115944
rect 289 115400 69200 115664
rect 880 115264 69200 115400
rect 880 115120 69120 115264
rect 289 114984 69120 115120
rect 289 114856 69200 114984
rect 880 114576 69200 114856
rect 289 114312 69200 114576
rect 880 114040 69200 114312
rect 880 114032 69120 114040
rect 289 113768 69120 114032
rect 880 113760 69120 113768
rect 880 113488 69200 113760
rect 289 113224 69200 113488
rect 880 112952 69200 113224
rect 880 112944 69120 112952
rect 289 112680 69120 112944
rect 880 112672 69120 112680
rect 880 112400 69200 112672
rect 289 112136 69200 112400
rect 880 111864 69200 112136
rect 880 111856 69120 111864
rect 289 111592 69120 111856
rect 880 111584 69120 111592
rect 880 111312 69200 111584
rect 289 111048 69200 111312
rect 880 110776 69200 111048
rect 880 110768 69120 110776
rect 289 110504 69120 110768
rect 880 110496 69120 110504
rect 880 110224 69200 110496
rect 289 109824 69200 110224
rect 880 109552 69200 109824
rect 880 109544 69120 109552
rect 289 109280 69120 109544
rect 880 109272 69120 109280
rect 880 109000 69200 109272
rect 289 108736 69200 109000
rect 880 108464 69200 108736
rect 880 108456 69120 108464
rect 289 108192 69120 108456
rect 880 108184 69120 108192
rect 880 107912 69200 108184
rect 289 107648 69200 107912
rect 880 107376 69200 107648
rect 880 107368 69120 107376
rect 289 107104 69120 107368
rect 880 107096 69120 107104
rect 880 106824 69200 107096
rect 289 106560 69200 106824
rect 880 106280 69200 106560
rect 289 106152 69200 106280
rect 289 106016 69120 106152
rect 880 105872 69120 106016
rect 880 105736 69200 105872
rect 289 105472 69200 105736
rect 880 105192 69200 105472
rect 289 105064 69200 105192
rect 289 104928 69120 105064
rect 880 104784 69120 104928
rect 880 104648 69200 104784
rect 289 104384 69200 104648
rect 880 104104 69200 104384
rect 289 103976 69200 104104
rect 289 103840 69120 103976
rect 880 103696 69120 103840
rect 880 103560 69200 103696
rect 289 103296 69200 103560
rect 880 103016 69200 103296
rect 289 102888 69200 103016
rect 289 102752 69120 102888
rect 880 102608 69120 102752
rect 880 102472 69200 102608
rect 289 102208 69200 102472
rect 880 101928 69200 102208
rect 289 101664 69200 101928
rect 880 101384 69120 101664
rect 289 101120 69200 101384
rect 880 100840 69200 101120
rect 289 100576 69200 100840
rect 880 100296 69120 100576
rect 289 100032 69200 100296
rect 880 99752 69200 100032
rect 289 99488 69200 99752
rect 880 99208 69120 99488
rect 289 98944 69200 99208
rect 880 98664 69200 98944
rect 289 98400 69200 98664
rect 880 98120 69120 98400
rect 289 97720 69200 98120
rect 880 97440 69200 97720
rect 289 97176 69200 97440
rect 880 96896 69120 97176
rect 289 96632 69200 96896
rect 880 96352 69200 96632
rect 289 96088 69200 96352
rect 880 95808 69120 96088
rect 289 95544 69200 95808
rect 880 95264 69200 95544
rect 289 95000 69200 95264
rect 880 94720 69120 95000
rect 289 94456 69200 94720
rect 880 94176 69200 94456
rect 289 93912 69200 94176
rect 880 93632 69120 93912
rect 289 93368 69200 93632
rect 880 93088 69200 93368
rect 289 92824 69200 93088
rect 880 92688 69200 92824
rect 880 92544 69120 92688
rect 289 92408 69120 92544
rect 289 92280 69200 92408
rect 880 92000 69200 92280
rect 289 91736 69200 92000
rect 880 91600 69200 91736
rect 880 91456 69120 91600
rect 289 91320 69120 91456
rect 289 91192 69200 91320
rect 880 90912 69200 91192
rect 289 90648 69200 90912
rect 880 90512 69200 90648
rect 880 90368 69120 90512
rect 289 90232 69120 90368
rect 289 90104 69200 90232
rect 880 89824 69200 90104
rect 289 89560 69200 89824
rect 880 89424 69200 89560
rect 880 89280 69120 89424
rect 289 89144 69120 89280
rect 289 89016 69200 89144
rect 880 88736 69200 89016
rect 289 88472 69200 88736
rect 880 88200 69200 88472
rect 880 88192 69120 88200
rect 289 87928 69120 88192
rect 880 87920 69120 87928
rect 880 87648 69200 87920
rect 289 87384 69200 87648
rect 880 87112 69200 87384
rect 880 87104 69120 87112
rect 289 86840 69120 87104
rect 880 86832 69120 86840
rect 880 86560 69200 86832
rect 289 86296 69200 86560
rect 880 86024 69200 86296
rect 880 86016 69120 86024
rect 289 85744 69120 86016
rect 289 85616 69200 85744
rect 880 85336 69200 85616
rect 289 85072 69200 85336
rect 880 84936 69200 85072
rect 880 84792 69120 84936
rect 289 84656 69120 84792
rect 289 84528 69200 84656
rect 880 84248 69200 84528
rect 289 83984 69200 84248
rect 880 83712 69200 83984
rect 880 83704 69120 83712
rect 289 83440 69120 83704
rect 880 83432 69120 83440
rect 880 83160 69200 83432
rect 289 82896 69200 83160
rect 880 82624 69200 82896
rect 880 82616 69120 82624
rect 289 82352 69120 82616
rect 880 82344 69120 82352
rect 880 82072 69200 82344
rect 289 81808 69200 82072
rect 880 81536 69200 81808
rect 880 81528 69120 81536
rect 289 81264 69120 81528
rect 880 81256 69120 81264
rect 880 80984 69200 81256
rect 289 80720 69200 80984
rect 880 80448 69200 80720
rect 880 80440 69120 80448
rect 289 80176 69120 80440
rect 880 80168 69120 80176
rect 880 79896 69200 80168
rect 289 79632 69200 79896
rect 880 79352 69200 79632
rect 289 79224 69200 79352
rect 289 79088 69120 79224
rect 880 78944 69120 79088
rect 880 78808 69200 78944
rect 289 78544 69200 78808
rect 880 78264 69200 78544
rect 289 78136 69200 78264
rect 289 78000 69120 78136
rect 880 77856 69120 78000
rect 880 77720 69200 77856
rect 289 77456 69200 77720
rect 880 77176 69200 77456
rect 289 77048 69200 77176
rect 289 76912 69120 77048
rect 880 76768 69120 76912
rect 880 76632 69200 76768
rect 289 76368 69200 76632
rect 880 76088 69200 76368
rect 289 75960 69200 76088
rect 289 75824 69120 75960
rect 880 75680 69120 75824
rect 880 75544 69200 75680
rect 289 75280 69200 75544
rect 880 75000 69200 75280
rect 289 74736 69200 75000
rect 880 74456 69120 74736
rect 289 74192 69200 74456
rect 880 73912 69200 74192
rect 289 73648 69200 73912
rect 289 73512 69120 73648
rect 880 73368 69120 73512
rect 880 73232 69200 73368
rect 289 72968 69200 73232
rect 880 72688 69200 72968
rect 289 72560 69200 72688
rect 289 72424 69120 72560
rect 880 72280 69120 72424
rect 880 72144 69200 72280
rect 289 71880 69200 72144
rect 880 71600 69200 71880
rect 289 71472 69200 71600
rect 289 71336 69120 71472
rect 880 71192 69120 71336
rect 880 71056 69200 71192
rect 289 70792 69200 71056
rect 880 70512 69200 70792
rect 289 70248 69200 70512
rect 880 69968 69120 70248
rect 289 69704 69200 69968
rect 880 69424 69200 69704
rect 289 69160 69200 69424
rect 880 68880 69120 69160
rect 289 68616 69200 68880
rect 880 68336 69200 68616
rect 289 68072 69200 68336
rect 880 67792 69120 68072
rect 289 67528 69200 67792
rect 880 67248 69200 67528
rect 289 66984 69200 67248
rect 880 66704 69120 66984
rect 289 66440 69200 66704
rect 880 66160 69200 66440
rect 289 65896 69200 66160
rect 880 65760 69200 65896
rect 880 65616 69120 65760
rect 289 65480 69120 65616
rect 289 65352 69200 65480
rect 880 65072 69200 65352
rect 289 64808 69200 65072
rect 880 64672 69200 64808
rect 880 64528 69120 64672
rect 289 64392 69120 64528
rect 289 64264 69200 64392
rect 880 63984 69200 64264
rect 289 63720 69200 63984
rect 880 63584 69200 63720
rect 880 63440 69120 63584
rect 289 63304 69120 63440
rect 289 63176 69200 63304
rect 880 62896 69200 63176
rect 289 62632 69200 62896
rect 880 62496 69200 62632
rect 880 62352 69120 62496
rect 289 62216 69120 62352
rect 289 62088 69200 62216
rect 880 61808 69200 62088
rect 289 61408 69200 61808
rect 880 61272 69200 61408
rect 880 61128 69120 61272
rect 289 60992 69120 61128
rect 289 60864 69200 60992
rect 880 60584 69200 60864
rect 289 60320 69200 60584
rect 880 60184 69200 60320
rect 880 60040 69120 60184
rect 289 59904 69120 60040
rect 289 59776 69200 59904
rect 880 59496 69200 59776
rect 289 59232 69200 59496
rect 880 59096 69200 59232
rect 880 58952 69120 59096
rect 289 58816 69120 58952
rect 289 58688 69200 58816
rect 880 58408 69200 58688
rect 289 58144 69200 58408
rect 880 58008 69200 58144
rect 880 57864 69120 58008
rect 289 57728 69120 57864
rect 289 57600 69200 57728
rect 880 57320 69200 57600
rect 289 57056 69200 57320
rect 880 56784 69200 57056
rect 880 56776 69120 56784
rect 289 56512 69120 56776
rect 880 56504 69120 56512
rect 880 56232 69200 56504
rect 289 55968 69200 56232
rect 880 55696 69200 55968
rect 880 55688 69120 55696
rect 289 55424 69120 55688
rect 880 55416 69120 55424
rect 880 55144 69200 55416
rect 289 54880 69200 55144
rect 880 54608 69200 54880
rect 880 54600 69120 54608
rect 289 54336 69120 54600
rect 880 54328 69120 54336
rect 880 54056 69200 54328
rect 289 53792 69200 54056
rect 880 53512 69200 53792
rect 289 53384 69200 53512
rect 289 53248 69120 53384
rect 880 53104 69120 53248
rect 880 52968 69200 53104
rect 289 52704 69200 52968
rect 880 52424 69200 52704
rect 289 52296 69200 52424
rect 289 52160 69120 52296
rect 880 52016 69120 52160
rect 880 51880 69200 52016
rect 289 51616 69200 51880
rect 880 51336 69200 51616
rect 289 51208 69200 51336
rect 289 51072 69120 51208
rect 880 50928 69120 51072
rect 880 50792 69200 50928
rect 289 50528 69200 50792
rect 880 50248 69200 50528
rect 289 50120 69200 50248
rect 289 49984 69120 50120
rect 880 49840 69120 49984
rect 880 49704 69200 49840
rect 289 49440 69200 49704
rect 880 49160 69200 49440
rect 289 48896 69200 49160
rect 289 48760 69120 48896
rect 880 48616 69120 48760
rect 880 48480 69200 48616
rect 289 48216 69200 48480
rect 880 47936 69200 48216
rect 289 47808 69200 47936
rect 289 47672 69120 47808
rect 880 47528 69120 47672
rect 880 47392 69200 47528
rect 289 47128 69200 47392
rect 880 46848 69200 47128
rect 289 46720 69200 46848
rect 289 46584 69120 46720
rect 880 46440 69120 46584
rect 880 46304 69200 46440
rect 289 46040 69200 46304
rect 880 45760 69200 46040
rect 289 45632 69200 45760
rect 289 45496 69120 45632
rect 880 45352 69120 45496
rect 880 45216 69200 45352
rect 289 44952 69200 45216
rect 880 44672 69200 44952
rect 289 44408 69200 44672
rect 880 44128 69120 44408
rect 289 43864 69200 44128
rect 880 43584 69200 43864
rect 289 43320 69200 43584
rect 880 43040 69120 43320
rect 289 42776 69200 43040
rect 880 42496 69200 42776
rect 289 42232 69200 42496
rect 880 41952 69120 42232
rect 289 41688 69200 41952
rect 880 41408 69200 41688
rect 289 41144 69200 41408
rect 880 40864 69120 41144
rect 289 40600 69200 40864
rect 880 40320 69200 40600
rect 289 40056 69200 40320
rect 880 39920 69200 40056
rect 880 39776 69120 39920
rect 289 39640 69120 39776
rect 289 39512 69200 39640
rect 880 39232 69200 39512
rect 289 38968 69200 39232
rect 880 38832 69200 38968
rect 880 38688 69120 38832
rect 289 38552 69120 38688
rect 289 38424 69200 38552
rect 880 38144 69200 38424
rect 289 37880 69200 38144
rect 880 37744 69200 37880
rect 880 37600 69120 37744
rect 289 37464 69120 37600
rect 289 37336 69200 37464
rect 880 37056 69200 37336
rect 289 36656 69200 37056
rect 880 36376 69120 36656
rect 289 36112 69200 36376
rect 880 35832 69200 36112
rect 289 35568 69200 35832
rect 880 35432 69200 35568
rect 880 35288 69120 35432
rect 289 35152 69120 35288
rect 289 35024 69200 35152
rect 880 34744 69200 35024
rect 289 34480 69200 34744
rect 880 34344 69200 34480
rect 880 34200 69120 34344
rect 289 34064 69120 34200
rect 289 33936 69200 34064
rect 880 33656 69200 33936
rect 289 33392 69200 33656
rect 880 33256 69200 33392
rect 880 33112 69120 33256
rect 289 32976 69120 33112
rect 289 32848 69200 32976
rect 880 32568 69200 32848
rect 289 32304 69200 32568
rect 880 32168 69200 32304
rect 880 32024 69120 32168
rect 289 31888 69120 32024
rect 289 31760 69200 31888
rect 880 31480 69200 31760
rect 289 31216 69200 31480
rect 880 30944 69200 31216
rect 880 30936 69120 30944
rect 289 30672 69120 30936
rect 880 30664 69120 30672
rect 880 30392 69200 30664
rect 289 30128 69200 30392
rect 880 29856 69200 30128
rect 880 29848 69120 29856
rect 289 29584 69120 29848
rect 880 29576 69120 29584
rect 880 29304 69200 29576
rect 289 29040 69200 29304
rect 880 28768 69200 29040
rect 880 28760 69120 28768
rect 289 28496 69120 28760
rect 880 28488 69120 28496
rect 880 28216 69200 28488
rect 289 27952 69200 28216
rect 880 27680 69200 27952
rect 880 27672 69120 27680
rect 289 27408 69120 27672
rect 880 27400 69120 27408
rect 880 27128 69200 27400
rect 289 26864 69200 27128
rect 880 26584 69200 26864
rect 289 26456 69200 26584
rect 289 26320 69120 26456
rect 880 26176 69120 26320
rect 880 26040 69200 26176
rect 289 25776 69200 26040
rect 880 25496 69200 25776
rect 289 25368 69200 25496
rect 289 25232 69120 25368
rect 880 25088 69120 25232
rect 880 24952 69200 25088
rect 289 24552 69200 24952
rect 880 24280 69200 24552
rect 880 24272 69120 24280
rect 289 24008 69120 24272
rect 880 24000 69120 24008
rect 880 23728 69200 24000
rect 289 23464 69200 23728
rect 880 23192 69200 23464
rect 880 23184 69120 23192
rect 289 22920 69120 23184
rect 880 22912 69120 22920
rect 880 22640 69200 22912
rect 289 22376 69200 22640
rect 880 22096 69200 22376
rect 289 21968 69200 22096
rect 289 21832 69120 21968
rect 880 21688 69120 21832
rect 880 21552 69200 21688
rect 289 21288 69200 21552
rect 880 21008 69200 21288
rect 289 20880 69200 21008
rect 289 20744 69120 20880
rect 880 20600 69120 20744
rect 880 20464 69200 20600
rect 289 20200 69200 20464
rect 880 19920 69200 20200
rect 289 19792 69200 19920
rect 289 19656 69120 19792
rect 880 19512 69120 19656
rect 880 19376 69200 19512
rect 289 19112 69200 19376
rect 880 18832 69200 19112
rect 289 18704 69200 18832
rect 289 18568 69120 18704
rect 880 18424 69120 18568
rect 880 18288 69200 18424
rect 289 18024 69200 18288
rect 880 17744 69200 18024
rect 289 17480 69200 17744
rect 880 17200 69120 17480
rect 289 16936 69200 17200
rect 880 16656 69200 16936
rect 289 16392 69200 16656
rect 880 16112 69120 16392
rect 289 15848 69200 16112
rect 880 15568 69200 15848
rect 289 15304 69200 15568
rect 880 15024 69120 15304
rect 289 14760 69200 15024
rect 880 14480 69200 14760
rect 289 14216 69200 14480
rect 880 13936 69120 14216
rect 289 13672 69200 13936
rect 880 13392 69200 13672
rect 289 13128 69200 13392
rect 880 12992 69200 13128
rect 880 12848 69120 12992
rect 289 12712 69120 12848
rect 289 12448 69200 12712
rect 880 12168 69200 12448
rect 289 11904 69200 12168
rect 880 11624 69120 11904
rect 289 11360 69200 11624
rect 880 11080 69200 11360
rect 289 10816 69200 11080
rect 880 10536 69120 10816
rect 289 10272 69200 10536
rect 880 9992 69200 10272
rect 289 9728 69200 9992
rect 880 9448 69120 9728
rect 289 9184 69200 9448
rect 880 8904 69200 9184
rect 289 8640 69200 8904
rect 880 8504 69200 8640
rect 880 8360 69120 8504
rect 289 8224 69120 8360
rect 289 8096 69200 8224
rect 880 7816 69200 8096
rect 289 7552 69200 7816
rect 880 7416 69200 7552
rect 880 7272 69120 7416
rect 289 7136 69120 7272
rect 289 7008 69200 7136
rect 880 6728 69200 7008
rect 289 6464 69200 6728
rect 880 6328 69200 6464
rect 880 6184 69120 6328
rect 289 6048 69120 6184
rect 289 5920 69200 6048
rect 880 5640 69200 5920
rect 289 5376 69200 5640
rect 880 5240 69200 5376
rect 880 5096 69120 5240
rect 289 4960 69120 5096
rect 289 4832 69200 4960
rect 880 4552 69200 4832
rect 289 4288 69200 4552
rect 880 4016 69200 4288
rect 880 4008 69120 4016
rect 289 3744 69120 4008
rect 880 3736 69120 3744
rect 880 3464 69200 3736
rect 289 3200 69200 3464
rect 880 2928 69200 3200
rect 880 2920 69120 2928
rect 289 2656 69120 2920
rect 880 2648 69120 2656
rect 880 2376 69200 2648
rect 289 2112 69200 2376
rect 880 1840 69200 2112
rect 880 1832 69120 1840
rect 289 1568 69120 1832
rect 880 1560 69120 1568
rect 880 1288 69200 1560
rect 289 1024 69200 1288
rect 880 752 69200 1024
rect 880 744 69120 752
rect 289 480 69120 744
rect 880 472 69120 480
rect 880 307 69200 472
<< metal4 >>
rect 4208 2128 4528 217648
rect 19568 2128 19888 217648
rect 34928 2128 35248 217648
rect 50288 2128 50608 217648
rect 65648 2128 65968 217648
<< obsm4 >>
rect 430 3299 4128 217429
rect 4608 3299 19488 217429
rect 19968 3299 34848 217429
rect 35328 3299 50208 217429
rect 50688 3299 61765 217429
<< labels >>
rlabel metal2 s 10782 0 10838 800 6 master0_wb_ack_i
port 1 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 master0_wb_adr_o[0]
port 2 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 master0_wb_adr_o[10]
port 3 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 master0_wb_adr_o[11]
port 4 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 master0_wb_adr_o[12]
port 5 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 master0_wb_adr_o[13]
port 6 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 master0_wb_adr_o[14]
port 7 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 master0_wb_adr_o[15]
port 8 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 master0_wb_adr_o[16]
port 9 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 master0_wb_adr_o[17]
port 10 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 master0_wb_adr_o[18]
port 11 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 master0_wb_adr_o[19]
port 12 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 master0_wb_adr_o[1]
port 13 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 master0_wb_adr_o[20]
port 14 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 master0_wb_adr_o[21]
port 15 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 master0_wb_adr_o[22]
port 16 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 master0_wb_adr_o[23]
port 17 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 master0_wb_adr_o[24]
port 18 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 master0_wb_adr_o[25]
port 19 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 master0_wb_adr_o[26]
port 20 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 master0_wb_adr_o[27]
port 21 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 master0_wb_adr_o[2]
port 22 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 master0_wb_adr_o[3]
port 23 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 master0_wb_adr_o[4]
port 24 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 master0_wb_adr_o[5]
port 25 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 master0_wb_adr_o[6]
port 26 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 master0_wb_adr_o[7]
port 27 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 master0_wb_adr_o[8]
port 28 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 master0_wb_adr_o[9]
port 29 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 master0_wb_cyc_o
port 30 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 master0_wb_data_i[0]
port 31 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 master0_wb_data_i[10]
port 32 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 master0_wb_data_i[11]
port 33 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 master0_wb_data_i[12]
port 34 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 master0_wb_data_i[13]
port 35 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 master0_wb_data_i[14]
port 36 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 master0_wb_data_i[15]
port 37 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 master0_wb_data_i[16]
port 38 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 master0_wb_data_i[17]
port 39 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 master0_wb_data_i[18]
port 40 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 master0_wb_data_i[19]
port 41 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 master0_wb_data_i[1]
port 42 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 master0_wb_data_i[20]
port 43 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 master0_wb_data_i[21]
port 44 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 master0_wb_data_i[22]
port 45 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 master0_wb_data_i[23]
port 46 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 master0_wb_data_i[24]
port 47 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 master0_wb_data_i[25]
port 48 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 master0_wb_data_i[26]
port 49 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 master0_wb_data_i[27]
port 50 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 master0_wb_data_i[28]
port 51 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 master0_wb_data_i[29]
port 52 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 master0_wb_data_i[2]
port 53 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 master0_wb_data_i[30]
port 54 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 master0_wb_data_i[31]
port 55 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 master0_wb_data_i[3]
port 56 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 master0_wb_data_i[4]
port 57 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 master0_wb_data_i[5]
port 58 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 master0_wb_data_i[6]
port 59 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 master0_wb_data_i[7]
port 60 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 master0_wb_data_i[8]
port 61 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 master0_wb_data_i[9]
port 62 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 master0_wb_data_o[0]
port 63 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 master0_wb_data_o[10]
port 64 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 master0_wb_data_o[11]
port 65 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 master0_wb_data_o[12]
port 66 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 master0_wb_data_o[13]
port 67 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 master0_wb_data_o[14]
port 68 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 master0_wb_data_o[15]
port 69 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 master0_wb_data_o[16]
port 70 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 master0_wb_data_o[17]
port 71 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 master0_wb_data_o[18]
port 72 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 master0_wb_data_o[19]
port 73 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 master0_wb_data_o[1]
port 74 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 master0_wb_data_o[20]
port 75 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 master0_wb_data_o[21]
port 76 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 master0_wb_data_o[22]
port 77 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 master0_wb_data_o[23]
port 78 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 master0_wb_data_o[24]
port 79 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 master0_wb_data_o[25]
port 80 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 master0_wb_data_o[26]
port 81 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 master0_wb_data_o[27]
port 82 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 master0_wb_data_o[28]
port 83 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 master0_wb_data_o[29]
port 84 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 master0_wb_data_o[2]
port 85 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 master0_wb_data_o[30]
port 86 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 master0_wb_data_o[31]
port 87 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 master0_wb_data_o[3]
port 88 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 master0_wb_data_o[4]
port 89 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 master0_wb_data_o[5]
port 90 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 master0_wb_data_o[6]
port 91 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 master0_wb_data_o[7]
port 92 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 master0_wb_data_o[8]
port 93 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 master0_wb_data_o[9]
port 94 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 master0_wb_error_i
port 95 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 master0_wb_sel_o[0]
port 96 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 master0_wb_sel_o[1]
port 97 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 master0_wb_sel_o[2]
port 98 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 master0_wb_sel_o[3]
port 99 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 master0_wb_stall_i
port 100 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 master0_wb_stb_o
port 101 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 master0_wb_we_o
port 102 nsew signal input
rlabel metal3 s 0 110304 800 110424 6 master1_wb_ack_i
port 103 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 master1_wb_adr_o[0]
port 104 nsew signal input
rlabel metal3 s 0 132200 800 132320 6 master1_wb_adr_o[10]
port 105 nsew signal input
rlabel metal3 s 0 133832 800 133952 6 master1_wb_adr_o[11]
port 106 nsew signal input
rlabel metal3 s 0 135600 800 135720 6 master1_wb_adr_o[12]
port 107 nsew signal input
rlabel metal3 s 0 137232 800 137352 6 master1_wb_adr_o[13]
port 108 nsew signal input
rlabel metal3 s 0 138864 800 138984 6 master1_wb_adr_o[14]
port 109 nsew signal input
rlabel metal3 s 0 140496 800 140616 6 master1_wb_adr_o[15]
port 110 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 master1_wb_adr_o[16]
port 111 nsew signal input
rlabel metal3 s 0 143760 800 143880 6 master1_wb_adr_o[17]
port 112 nsew signal input
rlabel metal3 s 0 145392 800 145512 6 master1_wb_adr_o[18]
port 113 nsew signal input
rlabel metal3 s 0 147160 800 147280 6 master1_wb_adr_o[19]
port 114 nsew signal input
rlabel metal3 s 0 115744 800 115864 6 master1_wb_adr_o[1]
port 115 nsew signal input
rlabel metal3 s 0 148792 800 148912 6 master1_wb_adr_o[20]
port 116 nsew signal input
rlabel metal3 s 0 150424 800 150544 6 master1_wb_adr_o[21]
port 117 nsew signal input
rlabel metal3 s 0 152056 800 152176 6 master1_wb_adr_o[22]
port 118 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 master1_wb_adr_o[23]
port 119 nsew signal input
rlabel metal3 s 0 155320 800 155440 6 master1_wb_adr_o[24]
port 120 nsew signal input
rlabel metal3 s 0 156952 800 157072 6 master1_wb_adr_o[25]
port 121 nsew signal input
rlabel metal3 s 0 158584 800 158704 6 master1_wb_adr_o[26]
port 122 nsew signal input
rlabel metal3 s 0 160352 800 160472 6 master1_wb_adr_o[27]
port 123 nsew signal input
rlabel metal3 s 0 117920 800 118040 6 master1_wb_adr_o[2]
port 124 nsew signal input
rlabel metal3 s 0 120096 800 120216 6 master1_wb_adr_o[3]
port 125 nsew signal input
rlabel metal3 s 0 122272 800 122392 6 master1_wb_adr_o[4]
port 126 nsew signal input
rlabel metal3 s 0 124040 800 124160 6 master1_wb_adr_o[5]
port 127 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 master1_wb_adr_o[6]
port 128 nsew signal input
rlabel metal3 s 0 127304 800 127424 6 master1_wb_adr_o[7]
port 129 nsew signal input
rlabel metal3 s 0 128936 800 129056 6 master1_wb_adr_o[8]
port 130 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 master1_wb_adr_o[9]
port 131 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 master1_wb_cyc_o
port 132 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 master1_wb_data_i[0]
port 133 nsew signal output
rlabel metal3 s 0 132744 800 132864 6 master1_wb_data_i[10]
port 134 nsew signal output
rlabel metal3 s 0 134376 800 134496 6 master1_wb_data_i[11]
port 135 nsew signal output
rlabel metal3 s 0 136144 800 136264 6 master1_wb_data_i[12]
port 136 nsew signal output
rlabel metal3 s 0 137776 800 137896 6 master1_wb_data_i[13]
port 137 nsew signal output
rlabel metal3 s 0 139408 800 139528 6 master1_wb_data_i[14]
port 138 nsew signal output
rlabel metal3 s 0 141040 800 141160 6 master1_wb_data_i[15]
port 139 nsew signal output
rlabel metal3 s 0 142672 800 142792 6 master1_wb_data_i[16]
port 140 nsew signal output
rlabel metal3 s 0 144304 800 144424 6 master1_wb_data_i[17]
port 141 nsew signal output
rlabel metal3 s 0 145936 800 146056 6 master1_wb_data_i[18]
port 142 nsew signal output
rlabel metal3 s 0 147704 800 147824 6 master1_wb_data_i[19]
port 143 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 master1_wb_data_i[1]
port 144 nsew signal output
rlabel metal3 s 0 149336 800 149456 6 master1_wb_data_i[20]
port 145 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 master1_wb_data_i[21]
port 146 nsew signal output
rlabel metal3 s 0 152600 800 152720 6 master1_wb_data_i[22]
port 147 nsew signal output
rlabel metal3 s 0 154232 800 154352 6 master1_wb_data_i[23]
port 148 nsew signal output
rlabel metal3 s 0 155864 800 155984 6 master1_wb_data_i[24]
port 149 nsew signal output
rlabel metal3 s 0 157496 800 157616 6 master1_wb_data_i[25]
port 150 nsew signal output
rlabel metal3 s 0 159264 800 159384 6 master1_wb_data_i[26]
port 151 nsew signal output
rlabel metal3 s 0 160896 800 161016 6 master1_wb_data_i[27]
port 152 nsew signal output
rlabel metal3 s 0 161984 800 162104 6 master1_wb_data_i[28]
port 153 nsew signal output
rlabel metal3 s 0 163072 800 163192 6 master1_wb_data_i[29]
port 154 nsew signal output
rlabel metal3 s 0 118464 800 118584 6 master1_wb_data_i[2]
port 155 nsew signal output
rlabel metal3 s 0 164160 800 164280 6 master1_wb_data_i[30]
port 156 nsew signal output
rlabel metal3 s 0 165248 800 165368 6 master1_wb_data_i[31]
port 157 nsew signal output
rlabel metal3 s 0 120640 800 120760 6 master1_wb_data_i[3]
port 158 nsew signal output
rlabel metal3 s 0 122952 800 123072 6 master1_wb_data_i[4]
port 159 nsew signal output
rlabel metal3 s 0 124584 800 124704 6 master1_wb_data_i[5]
port 160 nsew signal output
rlabel metal3 s 0 126216 800 126336 6 master1_wb_data_i[6]
port 161 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 master1_wb_data_i[7]
port 162 nsew signal output
rlabel metal3 s 0 129480 800 129600 6 master1_wb_data_i[8]
port 163 nsew signal output
rlabel metal3 s 0 131112 800 131232 6 master1_wb_data_i[9]
port 164 nsew signal output
rlabel metal3 s 0 114656 800 114776 6 master1_wb_data_o[0]
port 165 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 master1_wb_data_o[10]
port 166 nsew signal input
rlabel metal3 s 0 135056 800 135176 6 master1_wb_data_o[11]
port 167 nsew signal input
rlabel metal3 s 0 136688 800 136808 6 master1_wb_data_o[12]
port 168 nsew signal input
rlabel metal3 s 0 138320 800 138440 6 master1_wb_data_o[13]
port 169 nsew signal input
rlabel metal3 s 0 139952 800 140072 6 master1_wb_data_o[14]
port 170 nsew signal input
rlabel metal3 s 0 141584 800 141704 6 master1_wb_data_o[15]
port 171 nsew signal input
rlabel metal3 s 0 143216 800 143336 6 master1_wb_data_o[16]
port 172 nsew signal input
rlabel metal3 s 0 144848 800 144968 6 master1_wb_data_o[17]
port 173 nsew signal input
rlabel metal3 s 0 146480 800 146600 6 master1_wb_data_o[18]
port 174 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 master1_wb_data_o[19]
port 175 nsew signal input
rlabel metal3 s 0 116832 800 116952 6 master1_wb_data_o[1]
port 176 nsew signal input
rlabel metal3 s 0 149880 800 150000 6 master1_wb_data_o[20]
port 177 nsew signal input
rlabel metal3 s 0 151512 800 151632 6 master1_wb_data_o[21]
port 178 nsew signal input
rlabel metal3 s 0 153144 800 153264 6 master1_wb_data_o[22]
port 179 nsew signal input
rlabel metal3 s 0 154776 800 154896 6 master1_wb_data_o[23]
port 180 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 master1_wb_data_o[24]
port 181 nsew signal input
rlabel metal3 s 0 158040 800 158160 6 master1_wb_data_o[25]
port 182 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 master1_wb_data_o[26]
port 183 nsew signal input
rlabel metal3 s 0 161440 800 161560 6 master1_wb_data_o[27]
port 184 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 master1_wb_data_o[28]
port 185 nsew signal input
rlabel metal3 s 0 163616 800 163736 6 master1_wb_data_o[29]
port 186 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 master1_wb_data_o[2]
port 187 nsew signal input
rlabel metal3 s 0 164704 800 164824 6 master1_wb_data_o[30]
port 188 nsew signal input
rlabel metal3 s 0 165792 800 165912 6 master1_wb_data_o[31]
port 189 nsew signal input
rlabel metal3 s 0 121184 800 121304 6 master1_wb_data_o[3]
port 190 nsew signal input
rlabel metal3 s 0 123496 800 123616 6 master1_wb_data_o[4]
port 191 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 master1_wb_data_o[5]
port 192 nsew signal input
rlabel metal3 s 0 126760 800 126880 6 master1_wb_data_o[6]
port 193 nsew signal input
rlabel metal3 s 0 128392 800 128512 6 master1_wb_data_o[7]
port 194 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 master1_wb_data_o[8]
port 195 nsew signal input
rlabel metal3 s 0 131656 800 131776 6 master1_wb_data_o[9]
port 196 nsew signal input
rlabel metal3 s 0 111392 800 111512 6 master1_wb_error_i
port 197 nsew signal output
rlabel metal3 s 0 115200 800 115320 6 master1_wb_sel_o[0]
port 198 nsew signal input
rlabel metal3 s 0 117376 800 117496 6 master1_wb_sel_o[1]
port 199 nsew signal input
rlabel metal3 s 0 119552 800 119672 6 master1_wb_sel_o[2]
port 200 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 master1_wb_sel_o[3]
port 201 nsew signal input
rlabel metal3 s 0 111936 800 112056 6 master1_wb_stall_i
port 202 nsew signal output
rlabel metal3 s 0 112480 800 112600 6 master1_wb_stb_o
port 203 nsew signal input
rlabel metal3 s 0 113024 800 113144 6 master1_wb_we_o
port 204 nsew signal input
rlabel metal3 s 0 280 800 400 6 master2_wb_ack_i
port 205 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 master2_wb_adr_o[0]
port 206 nsew signal input
rlabel metal3 s 0 22176 800 22296 6 master2_wb_adr_o[10]
port 207 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 master2_wb_adr_o[11]
port 208 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 master2_wb_adr_o[12]
port 209 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 master2_wb_adr_o[13]
port 210 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 master2_wb_adr_o[14]
port 211 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 master2_wb_adr_o[15]
port 212 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 master2_wb_adr_o[16]
port 213 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 master2_wb_adr_o[17]
port 214 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 master2_wb_adr_o[18]
port 215 nsew signal input
rlabel metal3 s 0 37136 800 37256 6 master2_wb_adr_o[19]
port 216 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 master2_wb_adr_o[1]
port 217 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 master2_wb_adr_o[20]
port 218 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 master2_wb_adr_o[21]
port 219 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 master2_wb_adr_o[22]
port 220 nsew signal input
rlabel metal3 s 0 43664 800 43784 6 master2_wb_adr_o[23]
port 221 nsew signal input
rlabel metal3 s 0 45296 800 45416 6 master2_wb_adr_o[24]
port 222 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 master2_wb_adr_o[25]
port 223 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 master2_wb_adr_o[26]
port 224 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 master2_wb_adr_o[27]
port 225 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 master2_wb_adr_o[2]
port 226 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 master2_wb_adr_o[3]
port 227 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 master2_wb_adr_o[4]
port 228 nsew signal input
rlabel metal3 s 0 14016 800 14136 6 master2_wb_adr_o[5]
port 229 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 master2_wb_adr_o[6]
port 230 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 master2_wb_adr_o[7]
port 231 nsew signal input
rlabel metal3 s 0 18912 800 19032 6 master2_wb_adr_o[8]
port 232 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 master2_wb_adr_o[9]
port 233 nsew signal input
rlabel metal3 s 0 824 800 944 6 master2_wb_cyc_o
port 234 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 master2_wb_data_i[0]
port 235 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 master2_wb_data_i[10]
port 236 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 master2_wb_data_i[11]
port 237 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 master2_wb_data_i[12]
port 238 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 master2_wb_data_i[13]
port 239 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 master2_wb_data_i[14]
port 240 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 master2_wb_data_i[15]
port 241 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 master2_wb_data_i[16]
port 242 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 master2_wb_data_i[17]
port 243 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 master2_wb_data_i[18]
port 244 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 master2_wb_data_i[19]
port 245 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 master2_wb_data_i[1]
port 246 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 master2_wb_data_i[20]
port 247 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 master2_wb_data_i[21]
port 248 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 master2_wb_data_i[22]
port 249 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 master2_wb_data_i[23]
port 250 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 master2_wb_data_i[24]
port 251 nsew signal output
rlabel metal3 s 0 47472 800 47592 6 master2_wb_data_i[25]
port 252 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 master2_wb_data_i[26]
port 253 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 master2_wb_data_i[27]
port 254 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 master2_wb_data_i[28]
port 255 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 master2_wb_data_i[29]
port 256 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 master2_wb_data_i[2]
port 257 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 master2_wb_data_i[30]
port 258 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 master2_wb_data_i[31]
port 259 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 master2_wb_data_i[3]
port 260 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 master2_wb_data_i[4]
port 261 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 master2_wb_data_i[5]
port 262 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 master2_wb_data_i[6]
port 263 nsew signal output
rlabel metal3 s 0 17824 800 17944 6 master2_wb_data_i[7]
port 264 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 master2_wb_data_i[8]
port 265 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 master2_wb_data_i[9]
port 266 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 master2_wb_data_o[0]
port 267 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 master2_wb_data_o[10]
port 268 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 master2_wb_data_o[11]
port 269 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 master2_wb_data_o[12]
port 270 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 master2_wb_data_o[13]
port 271 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 master2_wb_data_o[14]
port 272 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 master2_wb_data_o[15]
port 273 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 master2_wb_data_o[16]
port 274 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 master2_wb_data_o[17]
port 275 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 master2_wb_data_o[18]
port 276 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 master2_wb_data_o[19]
port 277 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 master2_wb_data_o[1]
port 278 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 master2_wb_data_o[20]
port 279 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 master2_wb_data_o[21]
port 280 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 master2_wb_data_o[22]
port 281 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 master2_wb_data_o[23]
port 282 nsew signal input
rlabel metal3 s 0 46384 800 46504 6 master2_wb_data_o[24]
port 283 nsew signal input
rlabel metal3 s 0 48016 800 48136 6 master2_wb_data_o[25]
port 284 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 master2_wb_data_o[26]
port 285 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 master2_wb_data_o[27]
port 286 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 master2_wb_data_o[28]
port 287 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 master2_wb_data_o[29]
port 288 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 master2_wb_data_o[2]
port 289 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 master2_wb_data_o[30]
port 290 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 master2_wb_data_o[31]
port 291 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 master2_wb_data_o[3]
port 292 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 master2_wb_data_o[4]
port 293 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 master2_wb_data_o[5]
port 294 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 master2_wb_data_o[6]
port 295 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 master2_wb_data_o[7]
port 296 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 master2_wb_data_o[8]
port 297 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 master2_wb_data_o[9]
port 298 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 master2_wb_error_i
port 299 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 master2_wb_sel_o[0]
port 300 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 master2_wb_sel_o[1]
port 301 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 master2_wb_sel_o[2]
port 302 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 master2_wb_sel_o[3]
port 303 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 master2_wb_stall_i
port 304 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 master2_wb_stb_o
port 305 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 master2_wb_we_o
port 306 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 probe_master0_currentSlave[0]
port 307 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 probe_master0_currentSlave[1]
port 308 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 probe_master1_currentSlave[0]
port 309 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 probe_master1_currentSlave[1]
port 310 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 probe_master2_currentSlave[0]
port 311 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 probe_master2_currentSlave[1]
port 312 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 probe_master3_currentSlave[0]
port 313 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 probe_master3_currentSlave[1]
port 314 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 probe_slave0_currentMaster[0]
port 315 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 probe_slave0_currentMaster[1]
port 316 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 probe_slave1_currentMaster[0]
port 317 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 probe_slave1_currentMaster[1]
port 318 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 probe_slave2_currentMaster[0]
port 319 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 probe_slave2_currentMaster[1]
port 320 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 probe_slave3_currentMaster[0]
port 321 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 probe_slave3_currentMaster[1]
port 322 nsew signal output
rlabel metal3 s 0 166336 800 166456 6 slave0_wb_ack_o
port 323 nsew signal input
rlabel metal3 s 0 169600 800 169720 6 slave0_wb_adr_i[0]
port 324 nsew signal output
rlabel metal3 s 0 188368 800 188488 6 slave0_wb_adr_i[10]
port 325 nsew signal output
rlabel metal3 s 0 190000 800 190120 6 slave0_wb_adr_i[11]
port 326 nsew signal output
rlabel metal3 s 0 191632 800 191752 6 slave0_wb_adr_i[12]
port 327 nsew signal output
rlabel metal3 s 0 193264 800 193384 6 slave0_wb_adr_i[13]
port 328 nsew signal output
rlabel metal3 s 0 194896 800 195016 6 slave0_wb_adr_i[14]
port 329 nsew signal output
rlabel metal3 s 0 196664 800 196784 6 slave0_wb_adr_i[15]
port 330 nsew signal output
rlabel metal3 s 0 198296 800 198416 6 slave0_wb_adr_i[16]
port 331 nsew signal output
rlabel metal3 s 0 199928 800 200048 6 slave0_wb_adr_i[17]
port 332 nsew signal output
rlabel metal3 s 0 201560 800 201680 6 slave0_wb_adr_i[18]
port 333 nsew signal output
rlabel metal3 s 0 203192 800 203312 6 slave0_wb_adr_i[19]
port 334 nsew signal output
rlabel metal3 s 0 171912 800 172032 6 slave0_wb_adr_i[1]
port 335 nsew signal output
rlabel metal3 s 0 204824 800 204944 6 slave0_wb_adr_i[20]
port 336 nsew signal output
rlabel metal3 s 0 206456 800 206576 6 slave0_wb_adr_i[21]
port 337 nsew signal output
rlabel metal3 s 0 208224 800 208344 6 slave0_wb_adr_i[22]
port 338 nsew signal output
rlabel metal3 s 0 209856 800 209976 6 slave0_wb_adr_i[23]
port 339 nsew signal output
rlabel metal3 s 0 174088 800 174208 6 slave0_wb_adr_i[2]
port 340 nsew signal output
rlabel metal3 s 0 176264 800 176384 6 slave0_wb_adr_i[3]
port 341 nsew signal output
rlabel metal3 s 0 178440 800 178560 6 slave0_wb_adr_i[4]
port 342 nsew signal output
rlabel metal3 s 0 180072 800 180192 6 slave0_wb_adr_i[5]
port 343 nsew signal output
rlabel metal3 s 0 181704 800 181824 6 slave0_wb_adr_i[6]
port 344 nsew signal output
rlabel metal3 s 0 183336 800 183456 6 slave0_wb_adr_i[7]
port 345 nsew signal output
rlabel metal3 s 0 185104 800 185224 6 slave0_wb_adr_i[8]
port 346 nsew signal output
rlabel metal3 s 0 186736 800 186856 6 slave0_wb_adr_i[9]
port 347 nsew signal output
rlabel metal3 s 0 166880 800 167000 6 slave0_wb_cyc_i
port 348 nsew signal output
rlabel metal3 s 0 170144 800 170264 6 slave0_wb_data_i[0]
port 349 nsew signal output
rlabel metal3 s 0 188912 800 189032 6 slave0_wb_data_i[10]
port 350 nsew signal output
rlabel metal3 s 0 190544 800 190664 6 slave0_wb_data_i[11]
port 351 nsew signal output
rlabel metal3 s 0 192176 800 192296 6 slave0_wb_data_i[12]
port 352 nsew signal output
rlabel metal3 s 0 193808 800 193928 6 slave0_wb_data_i[13]
port 353 nsew signal output
rlabel metal3 s 0 195440 800 195560 6 slave0_wb_data_i[14]
port 354 nsew signal output
rlabel metal3 s 0 197208 800 197328 6 slave0_wb_data_i[15]
port 355 nsew signal output
rlabel metal3 s 0 198840 800 198960 6 slave0_wb_data_i[16]
port 356 nsew signal output
rlabel metal3 s 0 200472 800 200592 6 slave0_wb_data_i[17]
port 357 nsew signal output
rlabel metal3 s 0 202104 800 202224 6 slave0_wb_data_i[18]
port 358 nsew signal output
rlabel metal3 s 0 203736 800 203856 6 slave0_wb_data_i[19]
port 359 nsew signal output
rlabel metal3 s 0 172456 800 172576 6 slave0_wb_data_i[1]
port 360 nsew signal output
rlabel metal3 s 0 205368 800 205488 6 slave0_wb_data_i[20]
port 361 nsew signal output
rlabel metal3 s 0 207000 800 207120 6 slave0_wb_data_i[21]
port 362 nsew signal output
rlabel metal3 s 0 208768 800 208888 6 slave0_wb_data_i[22]
port 363 nsew signal output
rlabel metal3 s 0 210400 800 210520 6 slave0_wb_data_i[23]
port 364 nsew signal output
rlabel metal3 s 0 211488 800 211608 6 slave0_wb_data_i[24]
port 365 nsew signal output
rlabel metal3 s 0 212576 800 212696 6 slave0_wb_data_i[25]
port 366 nsew signal output
rlabel metal3 s 0 213664 800 213784 6 slave0_wb_data_i[26]
port 367 nsew signal output
rlabel metal3 s 0 214752 800 214872 6 slave0_wb_data_i[27]
port 368 nsew signal output
rlabel metal3 s 0 215840 800 215960 6 slave0_wb_data_i[28]
port 369 nsew signal output
rlabel metal3 s 0 216928 800 217048 6 slave0_wb_data_i[29]
port 370 nsew signal output
rlabel metal3 s 0 174632 800 174752 6 slave0_wb_data_i[2]
port 371 nsew signal output
rlabel metal3 s 0 218016 800 218136 6 slave0_wb_data_i[30]
port 372 nsew signal output
rlabel metal3 s 0 219104 800 219224 6 slave0_wb_data_i[31]
port 373 nsew signal output
rlabel metal3 s 0 176808 800 176928 6 slave0_wb_data_i[3]
port 374 nsew signal output
rlabel metal3 s 0 178984 800 179104 6 slave0_wb_data_i[4]
port 375 nsew signal output
rlabel metal3 s 0 180616 800 180736 6 slave0_wb_data_i[5]
port 376 nsew signal output
rlabel metal3 s 0 182248 800 182368 6 slave0_wb_data_i[6]
port 377 nsew signal output
rlabel metal3 s 0 184016 800 184136 6 slave0_wb_data_i[7]
port 378 nsew signal output
rlabel metal3 s 0 185648 800 185768 6 slave0_wb_data_i[8]
port 379 nsew signal output
rlabel metal3 s 0 187280 800 187400 6 slave0_wb_data_i[9]
port 380 nsew signal output
rlabel metal3 s 0 170688 800 170808 6 slave0_wb_data_o[0]
port 381 nsew signal input
rlabel metal3 s 0 189456 800 189576 6 slave0_wb_data_o[10]
port 382 nsew signal input
rlabel metal3 s 0 191088 800 191208 6 slave0_wb_data_o[11]
port 383 nsew signal input
rlabel metal3 s 0 192720 800 192840 6 slave0_wb_data_o[12]
port 384 nsew signal input
rlabel metal3 s 0 194352 800 194472 6 slave0_wb_data_o[13]
port 385 nsew signal input
rlabel metal3 s 0 196120 800 196240 6 slave0_wb_data_o[14]
port 386 nsew signal input
rlabel metal3 s 0 197752 800 197872 6 slave0_wb_data_o[15]
port 387 nsew signal input
rlabel metal3 s 0 199384 800 199504 6 slave0_wb_data_o[16]
port 388 nsew signal input
rlabel metal3 s 0 201016 800 201136 6 slave0_wb_data_o[17]
port 389 nsew signal input
rlabel metal3 s 0 202648 800 202768 6 slave0_wb_data_o[18]
port 390 nsew signal input
rlabel metal3 s 0 204280 800 204400 6 slave0_wb_data_o[19]
port 391 nsew signal input
rlabel metal3 s 0 173000 800 173120 6 slave0_wb_data_o[1]
port 392 nsew signal input
rlabel metal3 s 0 205912 800 206032 6 slave0_wb_data_o[20]
port 393 nsew signal input
rlabel metal3 s 0 207544 800 207664 6 slave0_wb_data_o[21]
port 394 nsew signal input
rlabel metal3 s 0 209312 800 209432 6 slave0_wb_data_o[22]
port 395 nsew signal input
rlabel metal3 s 0 210944 800 211064 6 slave0_wb_data_o[23]
port 396 nsew signal input
rlabel metal3 s 0 212032 800 212152 6 slave0_wb_data_o[24]
port 397 nsew signal input
rlabel metal3 s 0 213120 800 213240 6 slave0_wb_data_o[25]
port 398 nsew signal input
rlabel metal3 s 0 214208 800 214328 6 slave0_wb_data_o[26]
port 399 nsew signal input
rlabel metal3 s 0 215296 800 215416 6 slave0_wb_data_o[27]
port 400 nsew signal input
rlabel metal3 s 0 216384 800 216504 6 slave0_wb_data_o[28]
port 401 nsew signal input
rlabel metal3 s 0 217472 800 217592 6 slave0_wb_data_o[29]
port 402 nsew signal input
rlabel metal3 s 0 175176 800 175296 6 slave0_wb_data_o[2]
port 403 nsew signal input
rlabel metal3 s 0 218560 800 218680 6 slave0_wb_data_o[30]
port 404 nsew signal input
rlabel metal3 s 0 219648 800 219768 6 slave0_wb_data_o[31]
port 405 nsew signal input
rlabel metal3 s 0 177352 800 177472 6 slave0_wb_data_o[3]
port 406 nsew signal input
rlabel metal3 s 0 179528 800 179648 6 slave0_wb_data_o[4]
port 407 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 slave0_wb_data_o[5]
port 408 nsew signal input
rlabel metal3 s 0 182792 800 182912 6 slave0_wb_data_o[6]
port 409 nsew signal input
rlabel metal3 s 0 184560 800 184680 6 slave0_wb_data_o[7]
port 410 nsew signal input
rlabel metal3 s 0 186192 800 186312 6 slave0_wb_data_o[8]
port 411 nsew signal input
rlabel metal3 s 0 187824 800 187944 6 slave0_wb_data_o[9]
port 412 nsew signal input
rlabel metal3 s 0 167424 800 167544 6 slave0_wb_error_o
port 413 nsew signal input
rlabel metal3 s 0 171232 800 171352 6 slave0_wb_sel_i[0]
port 414 nsew signal output
rlabel metal3 s 0 173544 800 173664 6 slave0_wb_sel_i[1]
port 415 nsew signal output
rlabel metal3 s 0 175720 800 175840 6 slave0_wb_sel_i[2]
port 416 nsew signal output
rlabel metal3 s 0 177896 800 178016 6 slave0_wb_sel_i[3]
port 417 nsew signal output
rlabel metal3 s 0 167968 800 168088 6 slave0_wb_stall_o
port 418 nsew signal input
rlabel metal3 s 0 168512 800 168632 6 slave0_wb_stb_i
port 419 nsew signal output
rlabel metal3 s 0 169056 800 169176 6 slave0_wb_we_i
port 420 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 slave1_wb_ack_o
port 421 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 slave1_wb_adr_i[0]
port 422 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 slave1_wb_adr_i[10]
port 423 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 slave1_wb_adr_i[11]
port 424 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 slave1_wb_adr_i[12]
port 425 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 slave1_wb_adr_i[13]
port 426 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 slave1_wb_adr_i[14]
port 427 nsew signal output
rlabel metal3 s 0 86640 800 86760 6 slave1_wb_adr_i[15]
port 428 nsew signal output
rlabel metal3 s 0 88272 800 88392 6 slave1_wb_adr_i[16]
port 429 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 slave1_wb_adr_i[17]
port 430 nsew signal output
rlabel metal3 s 0 91536 800 91656 6 slave1_wb_adr_i[18]
port 431 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 slave1_wb_adr_i[19]
port 432 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 slave1_wb_adr_i[1]
port 433 nsew signal output
rlabel metal3 s 0 94800 800 94920 6 slave1_wb_adr_i[20]
port 434 nsew signal output
rlabel metal3 s 0 96432 800 96552 6 slave1_wb_adr_i[21]
port 435 nsew signal output
rlabel metal3 s 0 98200 800 98320 6 slave1_wb_adr_i[22]
port 436 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 slave1_wb_adr_i[23]
port 437 nsew signal output
rlabel metal3 s 0 64064 800 64184 6 slave1_wb_adr_i[2]
port 438 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 slave1_wb_adr_i[3]
port 439 nsew signal output
rlabel metal3 s 0 68416 800 68536 6 slave1_wb_adr_i[4]
port 440 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 slave1_wb_adr_i[5]
port 441 nsew signal output
rlabel metal3 s 0 71680 800 71800 6 slave1_wb_adr_i[6]
port 442 nsew signal output
rlabel metal3 s 0 73312 800 73432 6 slave1_wb_adr_i[7]
port 443 nsew signal output
rlabel metal3 s 0 75080 800 75200 6 slave1_wb_adr_i[8]
port 444 nsew signal output
rlabel metal3 s 0 76712 800 76832 6 slave1_wb_adr_i[9]
port 445 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 slave1_wb_cyc_i
port 446 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 slave1_wb_data_i[0]
port 447 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 slave1_wb_data_i[10]
port 448 nsew signal output
rlabel metal3 s 0 80520 800 80640 6 slave1_wb_data_i[11]
port 449 nsew signal output
rlabel metal3 s 0 82152 800 82272 6 slave1_wb_data_i[12]
port 450 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 slave1_wb_data_i[13]
port 451 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 slave1_wb_data_i[14]
port 452 nsew signal output
rlabel metal3 s 0 87184 800 87304 6 slave1_wb_data_i[15]
port 453 nsew signal output
rlabel metal3 s 0 88816 800 88936 6 slave1_wb_data_i[16]
port 454 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 slave1_wb_data_i[17]
port 455 nsew signal output
rlabel metal3 s 0 92080 800 92200 6 slave1_wb_data_i[18]
port 456 nsew signal output
rlabel metal3 s 0 93712 800 93832 6 slave1_wb_data_i[19]
port 457 nsew signal output
rlabel metal3 s 0 62432 800 62552 6 slave1_wb_data_i[1]
port 458 nsew signal output
rlabel metal3 s 0 95344 800 95464 6 slave1_wb_data_i[20]
port 459 nsew signal output
rlabel metal3 s 0 96976 800 97096 6 slave1_wb_data_i[21]
port 460 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 slave1_wb_data_i[22]
port 461 nsew signal output
rlabel metal3 s 0 100376 800 100496 6 slave1_wb_data_i[23]
port 462 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 slave1_wb_data_i[24]
port 463 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 slave1_wb_data_i[25]
port 464 nsew signal output
rlabel metal3 s 0 103640 800 103760 6 slave1_wb_data_i[26]
port 465 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 slave1_wb_data_i[27]
port 466 nsew signal output
rlabel metal3 s 0 105816 800 105936 6 slave1_wb_data_i[28]
port 467 nsew signal output
rlabel metal3 s 0 106904 800 107024 6 slave1_wb_data_i[29]
port 468 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 slave1_wb_data_i[2]
port 469 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 slave1_wb_data_i[30]
port 470 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 slave1_wb_data_i[31]
port 471 nsew signal output
rlabel metal3 s 0 66784 800 66904 6 slave1_wb_data_i[3]
port 472 nsew signal output
rlabel metal3 s 0 68960 800 69080 6 slave1_wb_data_i[4]
port 473 nsew signal output
rlabel metal3 s 0 70592 800 70712 6 slave1_wb_data_i[5]
port 474 nsew signal output
rlabel metal3 s 0 72224 800 72344 6 slave1_wb_data_i[6]
port 475 nsew signal output
rlabel metal3 s 0 73992 800 74112 6 slave1_wb_data_i[7]
port 476 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 slave1_wb_data_i[8]
port 477 nsew signal output
rlabel metal3 s 0 77256 800 77376 6 slave1_wb_data_i[9]
port 478 nsew signal output
rlabel metal3 s 0 60664 800 60784 6 slave1_wb_data_o[0]
port 479 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 slave1_wb_data_o[10]
port 480 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 slave1_wb_data_o[11]
port 481 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 slave1_wb_data_o[12]
port 482 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 slave1_wb_data_o[13]
port 483 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 slave1_wb_data_o[14]
port 484 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 slave1_wb_data_o[15]
port 485 nsew signal input
rlabel metal3 s 0 89360 800 89480 6 slave1_wb_data_o[16]
port 486 nsew signal input
rlabel metal3 s 0 90992 800 91112 6 slave1_wb_data_o[17]
port 487 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 slave1_wb_data_o[18]
port 488 nsew signal input
rlabel metal3 s 0 94256 800 94376 6 slave1_wb_data_o[19]
port 489 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 slave1_wb_data_o[1]
port 490 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 slave1_wb_data_o[20]
port 491 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 slave1_wb_data_o[21]
port 492 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 slave1_wb_data_o[22]
port 493 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 slave1_wb_data_o[23]
port 494 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 slave1_wb_data_o[24]
port 495 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 slave1_wb_data_o[25]
port 496 nsew signal input
rlabel metal3 s 0 104184 800 104304 6 slave1_wb_data_o[26]
port 497 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 slave1_wb_data_o[27]
port 498 nsew signal input
rlabel metal3 s 0 106360 800 106480 6 slave1_wb_data_o[28]
port 499 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 slave1_wb_data_o[29]
port 500 nsew signal input
rlabel metal3 s 0 65152 800 65272 6 slave1_wb_data_o[2]
port 501 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 slave1_wb_data_o[30]
port 502 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 slave1_wb_data_o[31]
port 503 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 slave1_wb_data_o[3]
port 504 nsew signal input
rlabel metal3 s 0 69504 800 69624 6 slave1_wb_data_o[4]
port 505 nsew signal input
rlabel metal3 s 0 71136 800 71256 6 slave1_wb_data_o[5]
port 506 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 slave1_wb_data_o[6]
port 507 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 slave1_wb_data_o[7]
port 508 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 slave1_wb_data_o[8]
port 509 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 slave1_wb_data_o[9]
port 510 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 slave1_wb_error_o
port 511 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 slave1_wb_sel_i[0]
port 512 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 slave1_wb_sel_i[1]
port 513 nsew signal output
rlabel metal3 s 0 65696 800 65816 6 slave1_wb_sel_i[2]
port 514 nsew signal output
rlabel metal3 s 0 67872 800 67992 6 slave1_wb_sel_i[3]
port 515 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 slave1_wb_stall_o
port 516 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 slave1_wb_stb_i
port 517 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 slave1_wb_we_i
port 518 nsew signal output
rlabel metal2 s 294 219200 350 220000 6 slave2_wb_ack_o
port 519 nsew signal input
rlabel metal2 s 4526 219200 4582 220000 6 slave2_wb_adr_i[0]
port 520 nsew signal output
rlabel metal2 s 28814 219200 28870 220000 6 slave2_wb_adr_i[10]
port 521 nsew signal output
rlabel metal2 s 30930 219200 30986 220000 6 slave2_wb_adr_i[11]
port 522 nsew signal output
rlabel metal2 s 33138 219200 33194 220000 6 slave2_wb_adr_i[12]
port 523 nsew signal output
rlabel metal2 s 35254 219200 35310 220000 6 slave2_wb_adr_i[13]
port 524 nsew signal output
rlabel metal2 s 37370 219200 37426 220000 6 slave2_wb_adr_i[14]
port 525 nsew signal output
rlabel metal2 s 39578 219200 39634 220000 6 slave2_wb_adr_i[15]
port 526 nsew signal output
rlabel metal2 s 41694 219200 41750 220000 6 slave2_wb_adr_i[16]
port 527 nsew signal output
rlabel metal2 s 43810 219200 43866 220000 6 slave2_wb_adr_i[17]
port 528 nsew signal output
rlabel metal2 s 45926 219200 45982 220000 6 slave2_wb_adr_i[18]
port 529 nsew signal output
rlabel metal2 s 48134 219200 48190 220000 6 slave2_wb_adr_i[19]
port 530 nsew signal output
rlabel metal2 s 7378 219200 7434 220000 6 slave2_wb_adr_i[1]
port 531 nsew signal output
rlabel metal2 s 50250 219200 50306 220000 6 slave2_wb_adr_i[20]
port 532 nsew signal output
rlabel metal2 s 52366 219200 52422 220000 6 slave2_wb_adr_i[21]
port 533 nsew signal output
rlabel metal2 s 54574 219200 54630 220000 6 slave2_wb_adr_i[22]
port 534 nsew signal output
rlabel metal2 s 56690 219200 56746 220000 6 slave2_wb_adr_i[23]
port 535 nsew signal output
rlabel metal2 s 10230 219200 10286 220000 6 slave2_wb_adr_i[2]
port 536 nsew signal output
rlabel metal2 s 13082 219200 13138 220000 6 slave2_wb_adr_i[3]
port 537 nsew signal output
rlabel metal2 s 15934 219200 15990 220000 6 slave2_wb_adr_i[4]
port 538 nsew signal output
rlabel metal2 s 18142 219200 18198 220000 6 slave2_wb_adr_i[5]
port 539 nsew signal output
rlabel metal2 s 20258 219200 20314 220000 6 slave2_wb_adr_i[6]
port 540 nsew signal output
rlabel metal2 s 22374 219200 22430 220000 6 slave2_wb_adr_i[7]
port 541 nsew signal output
rlabel metal2 s 24582 219200 24638 220000 6 slave2_wb_adr_i[8]
port 542 nsew signal output
rlabel metal2 s 26698 219200 26754 220000 6 slave2_wb_adr_i[9]
port 543 nsew signal output
rlabel metal2 s 938 219200 994 220000 6 slave2_wb_cyc_i
port 544 nsew signal output
rlabel metal2 s 5262 219200 5318 220000 6 slave2_wb_data_i[0]
port 545 nsew signal output
rlabel metal2 s 29550 219200 29606 220000 6 slave2_wb_data_i[10]
port 546 nsew signal output
rlabel metal2 s 31666 219200 31722 220000 6 slave2_wb_data_i[11]
port 547 nsew signal output
rlabel metal2 s 33782 219200 33838 220000 6 slave2_wb_data_i[12]
port 548 nsew signal output
rlabel metal2 s 35990 219200 36046 220000 6 slave2_wb_data_i[13]
port 549 nsew signal output
rlabel metal2 s 38106 219200 38162 220000 6 slave2_wb_data_i[14]
port 550 nsew signal output
rlabel metal2 s 40222 219200 40278 220000 6 slave2_wb_data_i[15]
port 551 nsew signal output
rlabel metal2 s 42430 219200 42486 220000 6 slave2_wb_data_i[16]
port 552 nsew signal output
rlabel metal2 s 44546 219200 44602 220000 6 slave2_wb_data_i[17]
port 553 nsew signal output
rlabel metal2 s 46662 219200 46718 220000 6 slave2_wb_data_i[18]
port 554 nsew signal output
rlabel metal2 s 48870 219200 48926 220000 6 slave2_wb_data_i[19]
port 555 nsew signal output
rlabel metal2 s 8114 219200 8170 220000 6 slave2_wb_data_i[1]
port 556 nsew signal output
rlabel metal2 s 50986 219200 51042 220000 6 slave2_wb_data_i[20]
port 557 nsew signal output
rlabel metal2 s 53102 219200 53158 220000 6 slave2_wb_data_i[21]
port 558 nsew signal output
rlabel metal2 s 55218 219200 55274 220000 6 slave2_wb_data_i[22]
port 559 nsew signal output
rlabel metal2 s 57426 219200 57482 220000 6 slave2_wb_data_i[23]
port 560 nsew signal output
rlabel metal2 s 58806 219200 58862 220000 6 slave2_wb_data_i[24]
port 561 nsew signal output
rlabel metal2 s 60278 219200 60334 220000 6 slave2_wb_data_i[25]
port 562 nsew signal output
rlabel metal2 s 61658 219200 61714 220000 6 slave2_wb_data_i[26]
port 563 nsew signal output
rlabel metal2 s 63130 219200 63186 220000 6 slave2_wb_data_i[27]
port 564 nsew signal output
rlabel metal2 s 64510 219200 64566 220000 6 slave2_wb_data_i[28]
port 565 nsew signal output
rlabel metal2 s 65982 219200 66038 220000 6 slave2_wb_data_i[29]
port 566 nsew signal output
rlabel metal2 s 10966 219200 11022 220000 6 slave2_wb_data_i[2]
port 567 nsew signal output
rlabel metal2 s 67362 219200 67418 220000 6 slave2_wb_data_i[30]
port 568 nsew signal output
rlabel metal2 s 68834 219200 68890 220000 6 slave2_wb_data_i[31]
port 569 nsew signal output
rlabel metal2 s 13818 219200 13874 220000 6 slave2_wb_data_i[3]
port 570 nsew signal output
rlabel metal2 s 16670 219200 16726 220000 6 slave2_wb_data_i[4]
port 571 nsew signal output
rlabel metal2 s 18786 219200 18842 220000 6 slave2_wb_data_i[5]
port 572 nsew signal output
rlabel metal2 s 20994 219200 21050 220000 6 slave2_wb_data_i[6]
port 573 nsew signal output
rlabel metal2 s 23110 219200 23166 220000 6 slave2_wb_data_i[7]
port 574 nsew signal output
rlabel metal2 s 25226 219200 25282 220000 6 slave2_wb_data_i[8]
port 575 nsew signal output
rlabel metal2 s 27434 219200 27490 220000 6 slave2_wb_data_i[9]
port 576 nsew signal output
rlabel metal2 s 5998 219200 6054 220000 6 slave2_wb_data_o[0]
port 577 nsew signal input
rlabel metal2 s 30286 219200 30342 220000 6 slave2_wb_data_o[10]
port 578 nsew signal input
rlabel metal2 s 32402 219200 32458 220000 6 slave2_wb_data_o[11]
port 579 nsew signal input
rlabel metal2 s 34518 219200 34574 220000 6 slave2_wb_data_o[12]
port 580 nsew signal input
rlabel metal2 s 36726 219200 36782 220000 6 slave2_wb_data_o[13]
port 581 nsew signal input
rlabel metal2 s 38842 219200 38898 220000 6 slave2_wb_data_o[14]
port 582 nsew signal input
rlabel metal2 s 40958 219200 41014 220000 6 slave2_wb_data_o[15]
port 583 nsew signal input
rlabel metal2 s 43074 219200 43130 220000 6 slave2_wb_data_o[16]
port 584 nsew signal input
rlabel metal2 s 45282 219200 45338 220000 6 slave2_wb_data_o[17]
port 585 nsew signal input
rlabel metal2 s 47398 219200 47454 220000 6 slave2_wb_data_o[18]
port 586 nsew signal input
rlabel metal2 s 49514 219200 49570 220000 6 slave2_wb_data_o[19]
port 587 nsew signal input
rlabel metal2 s 8850 219200 8906 220000 6 slave2_wb_data_o[1]
port 588 nsew signal input
rlabel metal2 s 51722 219200 51778 220000 6 slave2_wb_data_o[20]
port 589 nsew signal input
rlabel metal2 s 53838 219200 53894 220000 6 slave2_wb_data_o[21]
port 590 nsew signal input
rlabel metal2 s 55954 219200 56010 220000 6 slave2_wb_data_o[22]
port 591 nsew signal input
rlabel metal2 s 58070 219200 58126 220000 6 slave2_wb_data_o[23]
port 592 nsew signal input
rlabel metal2 s 59542 219200 59598 220000 6 slave2_wb_data_o[24]
port 593 nsew signal input
rlabel metal2 s 61014 219200 61070 220000 6 slave2_wb_data_o[25]
port 594 nsew signal input
rlabel metal2 s 62394 219200 62450 220000 6 slave2_wb_data_o[26]
port 595 nsew signal input
rlabel metal2 s 63866 219200 63922 220000 6 slave2_wb_data_o[27]
port 596 nsew signal input
rlabel metal2 s 65246 219200 65302 220000 6 slave2_wb_data_o[28]
port 597 nsew signal input
rlabel metal2 s 66718 219200 66774 220000 6 slave2_wb_data_o[29]
port 598 nsew signal input
rlabel metal2 s 11702 219200 11758 220000 6 slave2_wb_data_o[2]
port 599 nsew signal input
rlabel metal2 s 68098 219200 68154 220000 6 slave2_wb_data_o[30]
port 600 nsew signal input
rlabel metal2 s 69570 219200 69626 220000 6 slave2_wb_data_o[31]
port 601 nsew signal input
rlabel metal2 s 14554 219200 14610 220000 6 slave2_wb_data_o[3]
port 602 nsew signal input
rlabel metal2 s 17406 219200 17462 220000 6 slave2_wb_data_o[4]
port 603 nsew signal input
rlabel metal2 s 19522 219200 19578 220000 6 slave2_wb_data_o[5]
port 604 nsew signal input
rlabel metal2 s 21638 219200 21694 220000 6 slave2_wb_data_o[6]
port 605 nsew signal input
rlabel metal2 s 23846 219200 23902 220000 6 slave2_wb_data_o[7]
port 606 nsew signal input
rlabel metal2 s 25962 219200 26018 220000 6 slave2_wb_data_o[8]
port 607 nsew signal input
rlabel metal2 s 28078 219200 28134 220000 6 slave2_wb_data_o[9]
port 608 nsew signal input
rlabel metal2 s 1674 219200 1730 220000 6 slave2_wb_error_o
port 609 nsew signal input
rlabel metal2 s 6642 219200 6698 220000 6 slave2_wb_sel_i[0]
port 610 nsew signal output
rlabel metal2 s 9494 219200 9550 220000 6 slave2_wb_sel_i[1]
port 611 nsew signal output
rlabel metal2 s 12438 219200 12494 220000 6 slave2_wb_sel_i[2]
port 612 nsew signal output
rlabel metal2 s 15290 219200 15346 220000 6 slave2_wb_sel_i[3]
port 613 nsew signal output
rlabel metal2 s 2410 219200 2466 220000 6 slave2_wb_stall_o
port 614 nsew signal input
rlabel metal2 s 3146 219200 3202 220000 6 slave2_wb_stb_i
port 615 nsew signal output
rlabel metal2 s 3790 219200 3846 220000 6 slave2_wb_we_i
port 616 nsew signal output
rlabel metal3 s 69200 110576 70000 110696 6 slave3_wb_ack_o
port 617 nsew signal input
rlabel metal3 s 69200 117240 70000 117360 6 slave3_wb_adr_i[0]
port 618 nsew signal output
rlabel metal3 s 69200 155456 70000 155576 6 slave3_wb_adr_i[10]
port 619 nsew signal output
rlabel metal3 s 69200 158720 70000 158840 6 slave3_wb_adr_i[11]
port 620 nsew signal output
rlabel metal3 s 69200 162120 70000 162240 6 slave3_wb_adr_i[12]
port 621 nsew signal output
rlabel metal3 s 69200 165520 70000 165640 6 slave3_wb_adr_i[13]
port 622 nsew signal output
rlabel metal3 s 69200 168920 70000 169040 6 slave3_wb_adr_i[14]
port 623 nsew signal output
rlabel metal3 s 69200 172320 70000 172440 6 slave3_wb_adr_i[15]
port 624 nsew signal output
rlabel metal3 s 69200 175584 70000 175704 6 slave3_wb_adr_i[16]
port 625 nsew signal output
rlabel metal3 s 69200 178984 70000 179104 6 slave3_wb_adr_i[17]
port 626 nsew signal output
rlabel metal3 s 69200 182384 70000 182504 6 slave3_wb_adr_i[18]
port 627 nsew signal output
rlabel metal3 s 69200 185784 70000 185904 6 slave3_wb_adr_i[19]
port 628 nsew signal output
rlabel metal3 s 69200 121728 70000 121848 6 slave3_wb_adr_i[1]
port 629 nsew signal output
rlabel metal3 s 69200 189048 70000 189168 6 slave3_wb_adr_i[20]
port 630 nsew signal output
rlabel metal3 s 69200 192448 70000 192568 6 slave3_wb_adr_i[21]
port 631 nsew signal output
rlabel metal3 s 69200 195848 70000 195968 6 slave3_wb_adr_i[22]
port 632 nsew signal output
rlabel metal3 s 69200 199248 70000 199368 6 slave3_wb_adr_i[23]
port 633 nsew signal output
rlabel metal3 s 69200 126216 70000 126336 6 slave3_wb_adr_i[2]
port 634 nsew signal output
rlabel metal3 s 69200 130704 70000 130824 6 slave3_wb_adr_i[3]
port 635 nsew signal output
rlabel metal3 s 69200 135192 70000 135312 6 slave3_wb_adr_i[4]
port 636 nsew signal output
rlabel metal3 s 69200 138592 70000 138712 6 slave3_wb_adr_i[5]
port 637 nsew signal output
rlabel metal3 s 69200 141992 70000 142112 6 slave3_wb_adr_i[6]
port 638 nsew signal output
rlabel metal3 s 69200 145256 70000 145376 6 slave3_wb_adr_i[7]
port 639 nsew signal output
rlabel metal3 s 69200 148656 70000 148776 6 slave3_wb_adr_i[8]
port 640 nsew signal output
rlabel metal3 s 69200 152056 70000 152176 6 slave3_wb_adr_i[9]
port 641 nsew signal output
rlabel metal3 s 69200 111664 70000 111784 6 slave3_wb_cyc_i
port 642 nsew signal output
rlabel metal3 s 69200 118328 70000 118448 6 slave3_wb_data_i[0]
port 643 nsew signal output
rlabel metal3 s 69200 156544 70000 156664 6 slave3_wb_data_i[10]
port 644 nsew signal output
rlabel metal3 s 69200 159944 70000 160064 6 slave3_wb_data_i[11]
port 645 nsew signal output
rlabel metal3 s 69200 163208 70000 163328 6 slave3_wb_data_i[12]
port 646 nsew signal output
rlabel metal3 s 69200 166608 70000 166728 6 slave3_wb_data_i[13]
port 647 nsew signal output
rlabel metal3 s 69200 170008 70000 170128 6 slave3_wb_data_i[14]
port 648 nsew signal output
rlabel metal3 s 69200 173408 70000 173528 6 slave3_wb_data_i[15]
port 649 nsew signal output
rlabel metal3 s 69200 176808 70000 176928 6 slave3_wb_data_i[16]
port 650 nsew signal output
rlabel metal3 s 69200 180072 70000 180192 6 slave3_wb_data_i[17]
port 651 nsew signal output
rlabel metal3 s 69200 183472 70000 183592 6 slave3_wb_data_i[18]
port 652 nsew signal output
rlabel metal3 s 69200 186872 70000 186992 6 slave3_wb_data_i[19]
port 653 nsew signal output
rlabel metal3 s 69200 122816 70000 122936 6 slave3_wb_data_i[1]
port 654 nsew signal output
rlabel metal3 s 69200 190272 70000 190392 6 slave3_wb_data_i[20]
port 655 nsew signal output
rlabel metal3 s 69200 193536 70000 193656 6 slave3_wb_data_i[21]
port 656 nsew signal output
rlabel metal3 s 69200 196936 70000 197056 6 slave3_wb_data_i[22]
port 657 nsew signal output
rlabel metal3 s 69200 200336 70000 200456 6 slave3_wb_data_i[23]
port 658 nsew signal output
rlabel metal3 s 69200 202512 70000 202632 6 slave3_wb_data_i[24]
port 659 nsew signal output
rlabel metal3 s 69200 204824 70000 204944 6 slave3_wb_data_i[25]
port 660 nsew signal output
rlabel metal3 s 69200 207000 70000 207120 6 slave3_wb_data_i[26]
port 661 nsew signal output
rlabel metal3 s 69200 209312 70000 209432 6 slave3_wb_data_i[27]
port 662 nsew signal output
rlabel metal3 s 69200 211488 70000 211608 6 slave3_wb_data_i[28]
port 663 nsew signal output
rlabel metal3 s 69200 213800 70000 213920 6 slave3_wb_data_i[29]
port 664 nsew signal output
rlabel metal3 s 69200 127304 70000 127424 6 slave3_wb_data_i[2]
port 665 nsew signal output
rlabel metal3 s 69200 215976 70000 216096 6 slave3_wb_data_i[30]
port 666 nsew signal output
rlabel metal3 s 69200 218288 70000 218408 6 slave3_wb_data_i[31]
port 667 nsew signal output
rlabel metal3 s 69200 131792 70000 131912 6 slave3_wb_data_i[3]
port 668 nsew signal output
rlabel metal3 s 69200 136280 70000 136400 6 slave3_wb_data_i[4]
port 669 nsew signal output
rlabel metal3 s 69200 139680 70000 139800 6 slave3_wb_data_i[5]
port 670 nsew signal output
rlabel metal3 s 69200 143080 70000 143200 6 slave3_wb_data_i[6]
port 671 nsew signal output
rlabel metal3 s 69200 146480 70000 146600 6 slave3_wb_data_i[7]
port 672 nsew signal output
rlabel metal3 s 69200 149744 70000 149864 6 slave3_wb_data_i[8]
port 673 nsew signal output
rlabel metal3 s 69200 153144 70000 153264 6 slave3_wb_data_i[9]
port 674 nsew signal output
rlabel metal3 s 69200 119552 70000 119672 6 slave3_wb_data_o[0]
port 675 nsew signal input
rlabel metal3 s 69200 157632 70000 157752 6 slave3_wb_data_o[10]
port 676 nsew signal input
rlabel metal3 s 69200 161032 70000 161152 6 slave3_wb_data_o[11]
port 677 nsew signal input
rlabel metal3 s 69200 164432 70000 164552 6 slave3_wb_data_o[12]
port 678 nsew signal input
rlabel metal3 s 69200 167832 70000 167952 6 slave3_wb_data_o[13]
port 679 nsew signal input
rlabel metal3 s 69200 171096 70000 171216 6 slave3_wb_data_o[14]
port 680 nsew signal input
rlabel metal3 s 69200 174496 70000 174616 6 slave3_wb_data_o[15]
port 681 nsew signal input
rlabel metal3 s 69200 177896 70000 178016 6 slave3_wb_data_o[16]
port 682 nsew signal input
rlabel metal3 s 69200 181296 70000 181416 6 slave3_wb_data_o[17]
port 683 nsew signal input
rlabel metal3 s 69200 184560 70000 184680 6 slave3_wb_data_o[18]
port 684 nsew signal input
rlabel metal3 s 69200 187960 70000 188080 6 slave3_wb_data_o[19]
port 685 nsew signal input
rlabel metal3 s 69200 124040 70000 124160 6 slave3_wb_data_o[1]
port 686 nsew signal input
rlabel metal3 s 69200 191360 70000 191480 6 slave3_wb_data_o[20]
port 687 nsew signal input
rlabel metal3 s 69200 194760 70000 194880 6 slave3_wb_data_o[21]
port 688 nsew signal input
rlabel metal3 s 69200 198024 70000 198144 6 slave3_wb_data_o[22]
port 689 nsew signal input
rlabel metal3 s 69200 201424 70000 201544 6 slave3_wb_data_o[23]
port 690 nsew signal input
rlabel metal3 s 69200 203736 70000 203856 6 slave3_wb_data_o[24]
port 691 nsew signal input
rlabel metal3 s 69200 205912 70000 206032 6 slave3_wb_data_o[25]
port 692 nsew signal input
rlabel metal3 s 69200 208224 70000 208344 6 slave3_wb_data_o[26]
port 693 nsew signal input
rlabel metal3 s 69200 210400 70000 210520 6 slave3_wb_data_o[27]
port 694 nsew signal input
rlabel metal3 s 69200 212712 70000 212832 6 slave3_wb_data_o[28]
port 695 nsew signal input
rlabel metal3 s 69200 214888 70000 215008 6 slave3_wb_data_o[29]
port 696 nsew signal input
rlabel metal3 s 69200 128528 70000 128648 6 slave3_wb_data_o[2]
port 697 nsew signal input
rlabel metal3 s 69200 217200 70000 217320 6 slave3_wb_data_o[30]
port 698 nsew signal input
rlabel metal3 s 69200 219376 70000 219496 6 slave3_wb_data_o[31]
port 699 nsew signal input
rlabel metal3 s 69200 133016 70000 133136 6 slave3_wb_data_o[3]
port 700 nsew signal input
rlabel metal3 s 69200 137504 70000 137624 6 slave3_wb_data_o[4]
port 701 nsew signal input
rlabel metal3 s 69200 140768 70000 140888 6 slave3_wb_data_o[5]
port 702 nsew signal input
rlabel metal3 s 69200 144168 70000 144288 6 slave3_wb_data_o[6]
port 703 nsew signal input
rlabel metal3 s 69200 147568 70000 147688 6 slave3_wb_data_o[7]
port 704 nsew signal input
rlabel metal3 s 69200 150968 70000 151088 6 slave3_wb_data_o[8]
port 705 nsew signal input
rlabel metal3 s 69200 154232 70000 154352 6 slave3_wb_data_o[9]
port 706 nsew signal input
rlabel metal3 s 69200 112752 70000 112872 6 slave3_wb_error_o
port 707 nsew signal input
rlabel metal3 s 69200 120640 70000 120760 6 slave3_wb_sel_i[0]
port 708 nsew signal output
rlabel metal3 s 69200 125128 70000 125248 6 slave3_wb_sel_i[1]
port 709 nsew signal output
rlabel metal3 s 69200 129616 70000 129736 6 slave3_wb_sel_i[2]
port 710 nsew signal output
rlabel metal3 s 69200 134104 70000 134224 6 slave3_wb_sel_i[3]
port 711 nsew signal output
rlabel metal3 s 69200 113840 70000 113960 6 slave3_wb_stall_o
port 712 nsew signal input
rlabel metal3 s 69200 115064 70000 115184 6 slave3_wb_stb_i
port 713 nsew signal output
rlabel metal3 s 69200 116152 70000 116272 6 slave3_wb_we_i
port 714 nsew signal output
rlabel metal3 s 69200 552 70000 672 6 slave4_wb_ack_o
port 715 nsew signal input
rlabel metal3 s 69200 7216 70000 7336 6 slave4_wb_adr_i[0]
port 716 nsew signal output
rlabel metal3 s 69200 45432 70000 45552 6 slave4_wb_adr_i[10]
port 717 nsew signal output
rlabel metal3 s 69200 48696 70000 48816 6 slave4_wb_adr_i[11]
port 718 nsew signal output
rlabel metal3 s 69200 52096 70000 52216 6 slave4_wb_adr_i[12]
port 719 nsew signal output
rlabel metal3 s 69200 55496 70000 55616 6 slave4_wb_adr_i[13]
port 720 nsew signal output
rlabel metal3 s 69200 58896 70000 59016 6 slave4_wb_adr_i[14]
port 721 nsew signal output
rlabel metal3 s 69200 62296 70000 62416 6 slave4_wb_adr_i[15]
port 722 nsew signal output
rlabel metal3 s 69200 65560 70000 65680 6 slave4_wb_adr_i[16]
port 723 nsew signal output
rlabel metal3 s 69200 68960 70000 69080 6 slave4_wb_adr_i[17]
port 724 nsew signal output
rlabel metal3 s 69200 72360 70000 72480 6 slave4_wb_adr_i[18]
port 725 nsew signal output
rlabel metal3 s 69200 75760 70000 75880 6 slave4_wb_adr_i[19]
port 726 nsew signal output
rlabel metal3 s 69200 11704 70000 11824 6 slave4_wb_adr_i[1]
port 727 nsew signal output
rlabel metal3 s 69200 79024 70000 79144 6 slave4_wb_adr_i[20]
port 728 nsew signal output
rlabel metal3 s 69200 82424 70000 82544 6 slave4_wb_adr_i[21]
port 729 nsew signal output
rlabel metal3 s 69200 85824 70000 85944 6 slave4_wb_adr_i[22]
port 730 nsew signal output
rlabel metal3 s 69200 89224 70000 89344 6 slave4_wb_adr_i[23]
port 731 nsew signal output
rlabel metal3 s 69200 16192 70000 16312 6 slave4_wb_adr_i[2]
port 732 nsew signal output
rlabel metal3 s 69200 20680 70000 20800 6 slave4_wb_adr_i[3]
port 733 nsew signal output
rlabel metal3 s 69200 25168 70000 25288 6 slave4_wb_adr_i[4]
port 734 nsew signal output
rlabel metal3 s 69200 28568 70000 28688 6 slave4_wb_adr_i[5]
port 735 nsew signal output
rlabel metal3 s 69200 31968 70000 32088 6 slave4_wb_adr_i[6]
port 736 nsew signal output
rlabel metal3 s 69200 35232 70000 35352 6 slave4_wb_adr_i[7]
port 737 nsew signal output
rlabel metal3 s 69200 38632 70000 38752 6 slave4_wb_adr_i[8]
port 738 nsew signal output
rlabel metal3 s 69200 42032 70000 42152 6 slave4_wb_adr_i[9]
port 739 nsew signal output
rlabel metal3 s 69200 1640 70000 1760 6 slave4_wb_cyc_i
port 740 nsew signal output
rlabel metal3 s 69200 8304 70000 8424 6 slave4_wb_data_i[0]
port 741 nsew signal output
rlabel metal3 s 69200 46520 70000 46640 6 slave4_wb_data_i[10]
port 742 nsew signal output
rlabel metal3 s 69200 49920 70000 50040 6 slave4_wb_data_i[11]
port 743 nsew signal output
rlabel metal3 s 69200 53184 70000 53304 6 slave4_wb_data_i[12]
port 744 nsew signal output
rlabel metal3 s 69200 56584 70000 56704 6 slave4_wb_data_i[13]
port 745 nsew signal output
rlabel metal3 s 69200 59984 70000 60104 6 slave4_wb_data_i[14]
port 746 nsew signal output
rlabel metal3 s 69200 63384 70000 63504 6 slave4_wb_data_i[15]
port 747 nsew signal output
rlabel metal3 s 69200 66784 70000 66904 6 slave4_wb_data_i[16]
port 748 nsew signal output
rlabel metal3 s 69200 70048 70000 70168 6 slave4_wb_data_i[17]
port 749 nsew signal output
rlabel metal3 s 69200 73448 70000 73568 6 slave4_wb_data_i[18]
port 750 nsew signal output
rlabel metal3 s 69200 76848 70000 76968 6 slave4_wb_data_i[19]
port 751 nsew signal output
rlabel metal3 s 69200 12792 70000 12912 6 slave4_wb_data_i[1]
port 752 nsew signal output
rlabel metal3 s 69200 80248 70000 80368 6 slave4_wb_data_i[20]
port 753 nsew signal output
rlabel metal3 s 69200 83512 70000 83632 6 slave4_wb_data_i[21]
port 754 nsew signal output
rlabel metal3 s 69200 86912 70000 87032 6 slave4_wb_data_i[22]
port 755 nsew signal output
rlabel metal3 s 69200 90312 70000 90432 6 slave4_wb_data_i[23]
port 756 nsew signal output
rlabel metal3 s 69200 92488 70000 92608 6 slave4_wb_data_i[24]
port 757 nsew signal output
rlabel metal3 s 69200 94800 70000 94920 6 slave4_wb_data_i[25]
port 758 nsew signal output
rlabel metal3 s 69200 96976 70000 97096 6 slave4_wb_data_i[26]
port 759 nsew signal output
rlabel metal3 s 69200 99288 70000 99408 6 slave4_wb_data_i[27]
port 760 nsew signal output
rlabel metal3 s 69200 101464 70000 101584 6 slave4_wb_data_i[28]
port 761 nsew signal output
rlabel metal3 s 69200 103776 70000 103896 6 slave4_wb_data_i[29]
port 762 nsew signal output
rlabel metal3 s 69200 17280 70000 17400 6 slave4_wb_data_i[2]
port 763 nsew signal output
rlabel metal3 s 69200 105952 70000 106072 6 slave4_wb_data_i[30]
port 764 nsew signal output
rlabel metal3 s 69200 108264 70000 108384 6 slave4_wb_data_i[31]
port 765 nsew signal output
rlabel metal3 s 69200 21768 70000 21888 6 slave4_wb_data_i[3]
port 766 nsew signal output
rlabel metal3 s 69200 26256 70000 26376 6 slave4_wb_data_i[4]
port 767 nsew signal output
rlabel metal3 s 69200 29656 70000 29776 6 slave4_wb_data_i[5]
port 768 nsew signal output
rlabel metal3 s 69200 33056 70000 33176 6 slave4_wb_data_i[6]
port 769 nsew signal output
rlabel metal3 s 69200 36456 70000 36576 6 slave4_wb_data_i[7]
port 770 nsew signal output
rlabel metal3 s 69200 39720 70000 39840 6 slave4_wb_data_i[8]
port 771 nsew signal output
rlabel metal3 s 69200 43120 70000 43240 6 slave4_wb_data_i[9]
port 772 nsew signal output
rlabel metal3 s 69200 9528 70000 9648 6 slave4_wb_data_o[0]
port 773 nsew signal input
rlabel metal3 s 69200 47608 70000 47728 6 slave4_wb_data_o[10]
port 774 nsew signal input
rlabel metal3 s 69200 51008 70000 51128 6 slave4_wb_data_o[11]
port 775 nsew signal input
rlabel metal3 s 69200 54408 70000 54528 6 slave4_wb_data_o[12]
port 776 nsew signal input
rlabel metal3 s 69200 57808 70000 57928 6 slave4_wb_data_o[13]
port 777 nsew signal input
rlabel metal3 s 69200 61072 70000 61192 6 slave4_wb_data_o[14]
port 778 nsew signal input
rlabel metal3 s 69200 64472 70000 64592 6 slave4_wb_data_o[15]
port 779 nsew signal input
rlabel metal3 s 69200 67872 70000 67992 6 slave4_wb_data_o[16]
port 780 nsew signal input
rlabel metal3 s 69200 71272 70000 71392 6 slave4_wb_data_o[17]
port 781 nsew signal input
rlabel metal3 s 69200 74536 70000 74656 6 slave4_wb_data_o[18]
port 782 nsew signal input
rlabel metal3 s 69200 77936 70000 78056 6 slave4_wb_data_o[19]
port 783 nsew signal input
rlabel metal3 s 69200 14016 70000 14136 6 slave4_wb_data_o[1]
port 784 nsew signal input
rlabel metal3 s 69200 81336 70000 81456 6 slave4_wb_data_o[20]
port 785 nsew signal input
rlabel metal3 s 69200 84736 70000 84856 6 slave4_wb_data_o[21]
port 786 nsew signal input
rlabel metal3 s 69200 88000 70000 88120 6 slave4_wb_data_o[22]
port 787 nsew signal input
rlabel metal3 s 69200 91400 70000 91520 6 slave4_wb_data_o[23]
port 788 nsew signal input
rlabel metal3 s 69200 93712 70000 93832 6 slave4_wb_data_o[24]
port 789 nsew signal input
rlabel metal3 s 69200 95888 70000 96008 6 slave4_wb_data_o[25]
port 790 nsew signal input
rlabel metal3 s 69200 98200 70000 98320 6 slave4_wb_data_o[26]
port 791 nsew signal input
rlabel metal3 s 69200 100376 70000 100496 6 slave4_wb_data_o[27]
port 792 nsew signal input
rlabel metal3 s 69200 102688 70000 102808 6 slave4_wb_data_o[28]
port 793 nsew signal input
rlabel metal3 s 69200 104864 70000 104984 6 slave4_wb_data_o[29]
port 794 nsew signal input
rlabel metal3 s 69200 18504 70000 18624 6 slave4_wb_data_o[2]
port 795 nsew signal input
rlabel metal3 s 69200 107176 70000 107296 6 slave4_wb_data_o[30]
port 796 nsew signal input
rlabel metal3 s 69200 109352 70000 109472 6 slave4_wb_data_o[31]
port 797 nsew signal input
rlabel metal3 s 69200 22992 70000 23112 6 slave4_wb_data_o[3]
port 798 nsew signal input
rlabel metal3 s 69200 27480 70000 27600 6 slave4_wb_data_o[4]
port 799 nsew signal input
rlabel metal3 s 69200 30744 70000 30864 6 slave4_wb_data_o[5]
port 800 nsew signal input
rlabel metal3 s 69200 34144 70000 34264 6 slave4_wb_data_o[6]
port 801 nsew signal input
rlabel metal3 s 69200 37544 70000 37664 6 slave4_wb_data_o[7]
port 802 nsew signal input
rlabel metal3 s 69200 40944 70000 41064 6 slave4_wb_data_o[8]
port 803 nsew signal input
rlabel metal3 s 69200 44208 70000 44328 6 slave4_wb_data_o[9]
port 804 nsew signal input
rlabel metal3 s 69200 2728 70000 2848 6 slave4_wb_error_o
port 805 nsew signal input
rlabel metal3 s 69200 10616 70000 10736 6 slave4_wb_sel_i[0]
port 806 nsew signal output
rlabel metal3 s 69200 15104 70000 15224 6 slave4_wb_sel_i[1]
port 807 nsew signal output
rlabel metal3 s 69200 19592 70000 19712 6 slave4_wb_sel_i[2]
port 808 nsew signal output
rlabel metal3 s 69200 24080 70000 24200 6 slave4_wb_sel_i[3]
port 809 nsew signal output
rlabel metal3 s 69200 3816 70000 3936 6 slave4_wb_stall_o
port 810 nsew signal input
rlabel metal3 s 69200 5040 70000 5160 6 slave4_wb_stb_i
port 811 nsew signal output
rlabel metal3 s 69200 6128 70000 6248 6 slave4_wb_we_i
port 812 nsew signal output
rlabel metal4 s 4208 2128 4528 217648 6 vccd1
port 813 nsew power input
rlabel metal4 s 34928 2128 35248 217648 6 vccd1
port 813 nsew power input
rlabel metal4 s 65648 2128 65968 217648 6 vccd1
port 813 nsew power input
rlabel metal4 s 19568 2128 19888 217648 6 vssd1
port 814 nsew ground input
rlabel metal4 s 50288 2128 50608 217648 6 vssd1
port 814 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 815 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 816 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 220000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13096680
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/WishboneInterconnect/runs/WishboneInterconnect/results/finishing/WishboneInterconnect.magic.gds
string GDS_START 714876
<< end >>

